magic
tech sky130A
magscale 1 2
timestamp 1608764397
<< checkpaint >>
rect -1260 -1260 18260 21260
<< locali >>
rect 12265 14943 12299 15113
rect 12265 9435 12299 9673
rect 12265 8279 12299 8381
rect 12265 2907 12299 3077
rect 12357 1479 12391 1853
<< viali >>
rect 5641 17289 5675 17323
rect 6929 17289 6963 17323
rect 10701 17289 10735 17323
rect 11437 17221 11471 17255
rect 2329 17153 2363 17187
rect 3157 17153 3191 17187
rect 4261 17153 4295 17187
rect 6285 17153 6319 17187
rect 7481 17153 7515 17187
rect 2063 17085 2097 17119
rect 2973 17085 3007 17119
rect 4077 17085 4111 17119
rect 4997 17085 5031 17119
rect 7297 17085 7331 17119
rect 8125 17085 8159 17119
rect 8861 17085 8895 17119
rect 9781 17085 9815 17119
rect 10517 17085 10551 17119
rect 11253 17085 11287 17119
rect 12633 17085 12667 17119
rect 6009 17017 6043 17051
rect 7389 17017 7423 17051
rect 6101 16949 6135 16983
rect 8309 16949 8343 16983
rect 9045 16949 9079 16983
rect 9965 16949 9999 16983
rect 12817 16949 12851 16983
rect 5273 16745 5307 16779
rect 7665 16745 7699 16779
rect 8033 16745 8067 16779
rect 12081 16745 12115 16779
rect 12817 16745 12851 16779
rect 13553 16745 13587 16779
rect 5641 16677 5675 16711
rect 8125 16677 8159 16711
rect 1777 16609 1811 16643
rect 2053 16609 2087 16643
rect 2697 16609 2731 16643
rect 4077 16609 4111 16643
rect 5181 16609 5215 16643
rect 5733 16609 5767 16643
rect 6837 16609 6871 16643
rect 8867 16609 8901 16643
rect 9689 16609 9723 16643
rect 10425 16609 10459 16643
rect 11161 16609 11195 16643
rect 11897 16609 11931 16643
rect 12633 16609 12667 16643
rect 13369 16609 13403 16643
rect 2973 16541 3007 16575
rect 4261 16541 4295 16575
rect 5825 16541 5859 16575
rect 6929 16541 6963 16575
rect 7021 16541 7055 16575
rect 8217 16541 8251 16575
rect 9045 16473 9079 16507
rect 11345 16473 11379 16507
rect 4997 16405 5031 16439
rect 6469 16405 6503 16439
rect 9873 16405 9907 16439
rect 10609 16405 10643 16439
rect 3985 16201 4019 16235
rect 8033 16201 8067 16235
rect 14105 16201 14139 16235
rect 9229 16133 9263 16167
rect 10609 16133 10643 16167
rect 11345 16133 11379 16167
rect 12633 16133 12667 16167
rect 4629 16065 4663 16099
rect 5733 16065 5767 16099
rect 7389 16065 7423 16099
rect 8677 16065 8711 16099
rect 9781 16065 9815 16099
rect 1777 15997 1811 16031
rect 2697 15997 2731 16031
rect 4353 15997 4387 16031
rect 5549 15997 5583 16031
rect 6653 15997 6687 16031
rect 8493 15997 8527 16031
rect 9597 15997 9631 16031
rect 9689 15997 9723 16031
rect 10425 15997 10459 16031
rect 11161 15997 11195 16031
rect 12449 15997 12483 16031
rect 13185 15997 13219 16031
rect 13921 15997 13955 16031
rect 2053 15929 2087 15963
rect 2973 15929 3007 15963
rect 4445 15929 4479 15963
rect 5641 15929 5675 15963
rect 8401 15929 8435 15963
rect 5181 15861 5215 15895
rect 6469 15861 6503 15895
rect 6837 15861 6871 15895
rect 7205 15861 7239 15895
rect 7297 15861 7331 15895
rect 13369 15861 13403 15895
rect 4721 15657 4755 15691
rect 6929 15657 6963 15691
rect 9321 15657 9355 15691
rect 13277 15657 13311 15691
rect 1961 15589 1995 15623
rect 7849 15589 7883 15623
rect 10057 15589 10091 15623
rect 1685 15521 1719 15555
rect 2615 15521 2649 15555
rect 3893 15521 3927 15555
rect 5549 15521 5583 15555
rect 5816 15521 5850 15555
rect 7757 15521 7791 15555
rect 8585 15521 8619 15555
rect 9505 15521 9539 15555
rect 10149 15521 10183 15555
rect 10885 15521 10919 15555
rect 11621 15521 11655 15555
rect 12357 15521 12391 15555
rect 13093 15521 13127 15555
rect 2881 15453 2915 15487
rect 4813 15453 4847 15487
rect 4997 15453 5031 15487
rect 7941 15453 7975 15487
rect 10241 15453 10275 15487
rect 8769 15385 8803 15419
rect 9689 15385 9723 15419
rect 11069 15385 11103 15419
rect 11805 15385 11839 15419
rect 3709 15317 3743 15351
rect 4353 15317 4387 15351
rect 7389 15317 7423 15351
rect 12541 15317 12575 15351
rect 2513 15113 2547 15147
rect 3709 15113 3743 15147
rect 8677 15113 8711 15147
rect 9873 15113 9907 15147
rect 11069 15113 11103 15147
rect 12265 15113 12299 15147
rect 12633 15113 12667 15147
rect 3065 14977 3099 15011
rect 4169 14977 4203 15011
rect 4353 14977 4387 15011
rect 9321 14977 9355 15011
rect 10425 14977 10459 15011
rect 11529 14977 11563 15011
rect 11621 14977 11655 15011
rect 1593 14909 1627 14943
rect 2973 14909 3007 14943
rect 4905 14909 4939 14943
rect 6837 14909 6871 14943
rect 7104 14909 7138 14943
rect 9045 14909 9079 14943
rect 10333 14909 10367 14943
rect 12265 14909 12299 14943
rect 12449 14909 12483 14943
rect 1869 14841 1903 14875
rect 2881 14841 2915 14875
rect 5172 14841 5206 14875
rect 4077 14773 4111 14807
rect 6285 14773 6319 14807
rect 8217 14773 8251 14807
rect 9137 14773 9171 14807
rect 10241 14773 10275 14807
rect 11437 14773 11471 14807
rect 13185 14773 13219 14807
rect 3249 14569 3283 14603
rect 9137 14569 9171 14603
rect 10885 14569 10919 14603
rect 11253 14569 11287 14603
rect 3157 14501 3191 14535
rect 10149 14501 10183 14535
rect 1869 14433 1903 14467
rect 4629 14433 4663 14467
rect 5457 14433 5491 14467
rect 5724 14433 5758 14467
rect 7553 14433 7587 14467
rect 9321 14433 9355 14467
rect 10057 14433 10091 14467
rect 12081 14433 12115 14467
rect 12817 14433 12851 14467
rect 2145 14365 2179 14399
rect 3433 14365 3467 14399
rect 4721 14365 4755 14399
rect 4905 14365 4939 14399
rect 7297 14365 7331 14399
rect 10241 14365 10275 14399
rect 11345 14365 11379 14399
rect 11437 14365 11471 14399
rect 13553 14365 13587 14399
rect 14197 14365 14231 14399
rect 8677 14297 8711 14331
rect 9689 14297 9723 14331
rect 13001 14297 13035 14331
rect 2789 14229 2823 14263
rect 4261 14229 4295 14263
rect 6837 14229 6871 14263
rect 12265 14229 12299 14263
rect 1869 14025 1903 14059
rect 4445 14025 4479 14059
rect 6285 14025 6319 14059
rect 10057 14025 10091 14059
rect 10517 14025 10551 14059
rect 12449 14025 12483 14059
rect 8217 13957 8251 13991
rect 2513 13889 2547 13923
rect 4905 13889 4939 13923
rect 8677 13889 8711 13923
rect 11161 13889 11195 13923
rect 13093 13889 13127 13923
rect 3065 13821 3099 13855
rect 5172 13821 5206 13855
rect 6837 13821 6871 13855
rect 14657 13821 14691 13855
rect 14933 13821 14967 13855
rect 2237 13753 2271 13787
rect 3332 13753 3366 13787
rect 7104 13753 7138 13787
rect 8922 13753 8956 13787
rect 10977 13753 11011 13787
rect 11713 13753 11747 13787
rect 12909 13753 12943 13787
rect 13645 13753 13679 13787
rect 2329 13685 2363 13719
rect 10885 13685 10919 13719
rect 12817 13685 12851 13719
rect 2053 13481 2087 13515
rect 2789 13481 2823 13515
rect 3157 13481 3191 13515
rect 9321 13481 9355 13515
rect 10057 13481 10091 13515
rect 10885 13481 10919 13515
rect 12081 13481 12115 13515
rect 13277 13481 13311 13515
rect 13737 13481 13771 13515
rect 14473 13481 14507 13515
rect 4813 13413 4847 13447
rect 7748 13413 7782 13447
rect 11345 13413 11379 13447
rect 13645 13413 13679 13447
rect 1961 13345 1995 13379
rect 5908 13345 5942 13379
rect 7481 13345 7515 13379
rect 9505 13345 9539 13379
rect 11253 13345 11287 13379
rect 12449 13345 12483 13379
rect 2237 13277 2271 13311
rect 3249 13277 3283 13311
rect 3341 13277 3375 13311
rect 4905 13277 4939 13311
rect 5089 13277 5123 13311
rect 5641 13277 5675 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 11529 13277 11563 13311
rect 12541 13277 12575 13311
rect 12725 13277 12759 13311
rect 13829 13277 13863 13311
rect 8861 13209 8895 13243
rect 1593 13141 1627 13175
rect 4445 13141 4479 13175
rect 7021 13141 7055 13175
rect 9689 13141 9723 13175
rect 2513 12937 2547 12971
rect 12449 12937 12483 12971
rect 3709 12869 3743 12903
rect 6285 12869 6319 12903
rect 8217 12869 8251 12903
rect 10057 12869 10091 12903
rect 10517 12869 10551 12903
rect 3157 12801 3191 12835
rect 4353 12801 4387 12835
rect 8677 12801 8711 12835
rect 11069 12801 11103 12835
rect 11713 12801 11747 12835
rect 13001 12801 13035 12835
rect 13829 12801 13863 12835
rect 1593 12733 1627 12767
rect 4077 12733 4111 12767
rect 4905 12733 4939 12767
rect 5172 12733 5206 12767
rect 6837 12733 6871 12767
rect 12817 12733 12851 12767
rect 12909 12733 12943 12767
rect 13645 12733 13679 12767
rect 14565 12733 14599 12767
rect 1869 12665 1903 12699
rect 2881 12665 2915 12699
rect 4169 12665 4203 12699
rect 7104 12665 7138 12699
rect 8944 12665 8978 12699
rect 10977 12665 11011 12699
rect 14841 12665 14875 12699
rect 2973 12597 3007 12631
rect 10885 12597 10919 12631
rect 1593 12393 1627 12427
rect 1961 12393 1995 12427
rect 2789 12393 2823 12427
rect 3157 12393 3191 12427
rect 4353 12393 4387 12427
rect 6929 12393 6963 12427
rect 8769 12393 8803 12427
rect 9229 12393 9263 12427
rect 9689 12393 9723 12427
rect 12081 12393 12115 12427
rect 12541 12393 12575 12427
rect 13277 12393 13311 12427
rect 14657 12393 14691 12427
rect 4721 12325 4755 12359
rect 7634 12325 7668 12359
rect 2053 12257 2087 12291
rect 5816 12257 5850 12291
rect 7389 12257 7423 12291
rect 9413 12257 9447 12291
rect 10057 12257 10091 12291
rect 11253 12257 11287 12291
rect 12449 12257 12483 12291
rect 13645 12257 13679 12291
rect 14473 12257 14507 12291
rect 2237 12189 2271 12223
rect 3249 12189 3283 12223
rect 3433 12189 3467 12223
rect 4813 12189 4847 12223
rect 4997 12189 5031 12223
rect 5549 12189 5583 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 11345 12189 11379 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 13737 12189 13771 12223
rect 13829 12189 13863 12223
rect 10885 12053 10919 12087
rect 1869 11849 1903 11883
rect 8217 11849 8251 11883
rect 10517 11849 10551 11883
rect 15025 11849 15059 11883
rect 12449 11781 12483 11815
rect 13645 11781 13679 11815
rect 2513 11713 2547 11747
rect 6837 11713 6871 11747
rect 11069 11713 11103 11747
rect 11713 11713 11747 11747
rect 13001 11713 13035 11747
rect 14197 11713 14231 11747
rect 2329 11645 2363 11679
rect 3065 11645 3099 11679
rect 4905 11645 4939 11679
rect 8677 11645 8711 11679
rect 12817 11645 12851 11679
rect 14841 11645 14875 11679
rect 2237 11577 2271 11611
rect 3332 11577 3366 11611
rect 5172 11577 5206 11611
rect 7082 11577 7116 11611
rect 8944 11577 8978 11611
rect 14013 11577 14047 11611
rect 4445 11509 4479 11543
rect 6285 11509 6319 11543
rect 10057 11509 10091 11543
rect 10885 11509 10919 11543
rect 10977 11509 11011 11543
rect 12909 11509 12943 11543
rect 14105 11509 14139 11543
rect 1593 11305 1627 11339
rect 2053 11305 2087 11339
rect 2789 11305 2823 11339
rect 3157 11305 3191 11339
rect 4077 11305 4111 11339
rect 4537 11305 4571 11339
rect 6653 11305 6687 11339
rect 8493 11305 8527 11339
rect 10057 11305 10091 11339
rect 12449 11305 12483 11339
rect 13277 11305 13311 11339
rect 2697 11237 2731 11271
rect 3249 11237 3283 11271
rect 5518 11237 5552 11271
rect 7358 11237 7392 11271
rect 8953 11237 8987 11271
rect 10149 11237 10183 11271
rect 1961 11169 1995 11203
rect 4445 11169 4479 11203
rect 7113 11169 7147 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 12541 11169 12575 11203
rect 13645 11169 13679 11203
rect 14473 11169 14507 11203
rect 2237 11101 2271 11135
rect 3433 11101 3467 11135
rect 4721 11101 4755 11135
rect 5273 11101 5307 11135
rect 10241 11101 10275 11135
rect 11437 11101 11471 11135
rect 12633 11101 12667 11135
rect 13737 11101 13771 11135
rect 13921 11101 13955 11135
rect 9689 11033 9723 11067
rect 14657 11033 14691 11067
rect 10885 10965 10919 10999
rect 12081 10965 12115 10999
rect 1869 10761 1903 10795
rect 4997 10761 5031 10795
rect 10057 10761 10091 10795
rect 13645 10761 13679 10795
rect 4445 10693 4479 10727
rect 2513 10625 2547 10659
rect 5273 10625 5307 10659
rect 6837 10625 6871 10659
rect 10977 10625 11011 10659
rect 11161 10625 11195 10659
rect 11713 10625 11747 10659
rect 12909 10625 12943 10659
rect 13093 10625 13127 10659
rect 14105 10625 14139 10659
rect 14197 10625 14231 10659
rect 3065 10557 3099 10591
rect 5181 10557 5215 10591
rect 8677 10557 8711 10591
rect 12817 10557 12851 10591
rect 14841 10557 14875 10591
rect 2329 10489 2363 10523
rect 3332 10489 3366 10523
rect 5518 10489 5552 10523
rect 7082 10489 7116 10523
rect 8944 10489 8978 10523
rect 2237 10421 2271 10455
rect 6653 10421 6687 10455
rect 8217 10421 8251 10455
rect 10517 10421 10551 10455
rect 10885 10421 10919 10455
rect 12449 10421 12483 10455
rect 14013 10421 14047 10455
rect 15025 10421 15059 10455
rect 1593 10217 1627 10251
rect 2053 10217 2087 10251
rect 5825 10217 5859 10251
rect 7297 10217 7331 10251
rect 9045 10217 9079 10251
rect 10149 10217 10183 10251
rect 10885 10217 10919 10251
rect 11253 10217 11287 10251
rect 12449 10217 12483 10251
rect 13737 10217 13771 10251
rect 1961 10149 1995 10183
rect 4712 10149 4746 10183
rect 3157 10081 3191 10115
rect 3249 10081 3283 10115
rect 6184 10081 6218 10115
rect 7932 10081 7966 10115
rect 10057 10081 10091 10115
rect 13645 10081 13679 10115
rect 14473 10081 14507 10115
rect 2237 10013 2271 10047
rect 3341 10013 3375 10047
rect 4445 10013 4479 10047
rect 5917 10013 5951 10047
rect 7665 10013 7699 10047
rect 10333 10013 10367 10047
rect 11345 10013 11379 10047
rect 11437 10013 11471 10047
rect 12541 10013 12575 10047
rect 12725 10013 12759 10047
rect 13829 10013 13863 10047
rect 9689 9945 9723 9979
rect 2789 9877 2823 9911
rect 12081 9877 12115 9911
rect 13277 9877 13311 9911
rect 14657 9877 14691 9911
rect 6285 9673 6319 9707
rect 8677 9673 8711 9707
rect 11069 9673 11103 9707
rect 12265 9673 12299 9707
rect 4077 9605 4111 9639
rect 9873 9605 9907 9639
rect 2973 9537 3007 9571
rect 3801 9537 3835 9571
rect 4537 9537 4571 9571
rect 4721 9537 4755 9571
rect 6837 9537 6871 9571
rect 9321 9537 9355 9571
rect 10425 9537 10459 9571
rect 11713 9537 11747 9571
rect 1593 9469 1627 9503
rect 2789 9469 2823 9503
rect 4905 9469 4939 9503
rect 9045 9469 9079 9503
rect 10241 9469 10275 9503
rect 12909 9537 12943 9571
rect 13001 9537 13035 9571
rect 14197 9537 14231 9571
rect 14105 9469 14139 9503
rect 14841 9469 14875 9503
rect 1869 9401 1903 9435
rect 2881 9401 2915 9435
rect 3617 9401 3651 9435
rect 4445 9401 4479 9435
rect 5172 9401 5206 9435
rect 7104 9401 7138 9435
rect 11529 9401 11563 9435
rect 12265 9401 12299 9435
rect 12817 9401 12851 9435
rect 2421 9333 2455 9367
rect 3249 9333 3283 9367
rect 3709 9333 3743 9367
rect 8217 9333 8251 9367
rect 9137 9333 9171 9367
rect 10333 9333 10367 9367
rect 11437 9333 11471 9367
rect 12449 9333 12483 9367
rect 13645 9333 13679 9367
rect 14013 9333 14047 9367
rect 15025 9333 15059 9367
rect 1593 9129 1627 9163
rect 2053 9129 2087 9163
rect 3157 9129 3191 9163
rect 5457 9129 5491 9163
rect 10057 9129 10091 9163
rect 12081 9129 12115 9163
rect 13737 9129 13771 9163
rect 1961 9061 1995 9095
rect 7665 9061 7699 9095
rect 8024 9061 8058 9095
rect 4077 8993 4111 9027
rect 4333 8993 4367 9027
rect 5917 8993 5951 9027
rect 11253 8993 11287 9027
rect 12449 8993 12483 9027
rect 13645 8993 13679 9027
rect 14473 8993 14507 9027
rect 2237 8925 2271 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 7757 8925 7791 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 12541 8925 12575 8959
rect 12725 8925 12759 8959
rect 13829 8925 13863 8959
rect 2789 8857 2823 8891
rect 10885 8857 10919 8891
rect 9137 8789 9171 8823
rect 9689 8789 9723 8823
rect 13277 8789 13311 8823
rect 14657 8789 14691 8823
rect 6285 8585 6319 8619
rect 8677 8585 8711 8619
rect 11069 8585 11103 8619
rect 12449 8585 12483 8619
rect 13645 8585 13679 8619
rect 8217 8517 8251 8551
rect 15025 8517 15059 8551
rect 3157 8449 3191 8483
rect 4353 8449 4387 8483
rect 9229 8449 9263 8483
rect 10425 8449 10459 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 14197 8449 14231 8483
rect 1593 8381 1627 8415
rect 1869 8381 1903 8415
rect 4077 8381 4111 8415
rect 4905 8381 4939 8415
rect 6837 8381 6871 8415
rect 9137 8381 9171 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 14105 8381 14139 8415
rect 14841 8381 14875 8415
rect 2881 8313 2915 8347
rect 4169 8313 4203 8347
rect 5172 8313 5206 8347
rect 7104 8313 7138 8347
rect 10333 8313 10367 8347
rect 11437 8313 11471 8347
rect 2513 8245 2547 8279
rect 2973 8245 3007 8279
rect 3709 8245 3743 8279
rect 9045 8245 9079 8279
rect 9873 8245 9907 8279
rect 10241 8245 10275 8279
rect 12265 8245 12299 8279
rect 14013 8245 14047 8279
rect 1593 8041 1627 8075
rect 2789 8041 2823 8075
rect 10057 8041 10091 8075
rect 11253 8041 11287 8075
rect 11345 8041 11379 8075
rect 13277 8041 13311 8075
rect 13737 8041 13771 8075
rect 3157 7973 3191 8007
rect 10149 7973 10183 8007
rect 1961 7905 1995 7939
rect 4813 7905 4847 7939
rect 5641 7905 5675 7939
rect 5908 7905 5942 7939
rect 7481 7905 7515 7939
rect 7748 7905 7782 7939
rect 9505 7905 9539 7939
rect 12449 7905 12483 7939
rect 12541 7905 12575 7939
rect 13645 7905 13679 7939
rect 14473 7905 14507 7939
rect 2053 7837 2087 7871
rect 2237 7837 2271 7871
rect 3249 7837 3283 7871
rect 3433 7837 3467 7871
rect 4905 7837 4939 7871
rect 5089 7837 5123 7871
rect 10241 7837 10275 7871
rect 11437 7837 11471 7871
rect 12725 7837 12759 7871
rect 13921 7837 13955 7871
rect 10885 7769 10919 7803
rect 4445 7701 4479 7735
rect 7021 7701 7055 7735
rect 8861 7701 8895 7735
rect 9321 7701 9355 7735
rect 9689 7701 9723 7735
rect 12081 7701 12115 7735
rect 14657 7701 14691 7735
rect 1869 7497 1903 7531
rect 12449 7497 12483 7531
rect 4445 7429 4479 7463
rect 8217 7429 8251 7463
rect 10517 7429 10551 7463
rect 2513 7361 2547 7395
rect 6837 7361 6871 7395
rect 8677 7361 8711 7395
rect 10977 7361 11011 7395
rect 11161 7361 11195 7395
rect 11713 7361 11747 7395
rect 13001 7361 13035 7395
rect 14105 7361 14139 7395
rect 14197 7361 14231 7395
rect 2237 7293 2271 7327
rect 3065 7293 3099 7327
rect 4905 7293 4939 7327
rect 8933 7293 8967 7327
rect 10885 7293 10919 7327
rect 14841 7293 14875 7327
rect 3332 7225 3366 7259
rect 5172 7225 5206 7259
rect 7082 7225 7116 7259
rect 12817 7225 12851 7259
rect 2329 7157 2363 7191
rect 6285 7157 6319 7191
rect 10057 7157 10091 7191
rect 12909 7157 12943 7191
rect 13645 7157 13679 7191
rect 14013 7157 14047 7191
rect 15025 7157 15059 7191
rect 1961 6953 1995 6987
rect 13185 6953 13219 6987
rect 13921 6953 13955 6987
rect 3157 6885 3191 6919
rect 4997 6885 5031 6919
rect 6092 6885 6126 6919
rect 7932 6885 7966 6919
rect 9956 6885 9990 6919
rect 11897 6885 11931 6919
rect 13093 6885 13127 6919
rect 2053 6817 2087 6851
rect 7665 6817 7699 6851
rect 9689 6817 9723 6851
rect 14289 6817 14323 6851
rect 2237 6749 2271 6783
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 5089 6749 5123 6783
rect 5273 6749 5307 6783
rect 5825 6749 5859 6783
rect 11989 6749 12023 6783
rect 12081 6749 12115 6783
rect 13369 6749 13403 6783
rect 14381 6749 14415 6783
rect 14473 6749 14507 6783
rect 1593 6681 1627 6715
rect 12725 6681 12759 6715
rect 2789 6613 2823 6647
rect 4629 6613 4663 6647
rect 7205 6613 7239 6647
rect 9045 6613 9079 6647
rect 11069 6613 11103 6647
rect 11529 6613 11563 6647
rect 1869 6409 1903 6443
rect 10057 6409 10091 6443
rect 10517 6409 10551 6443
rect 12449 6409 12483 6443
rect 4445 6341 4479 6375
rect 2421 6273 2455 6307
rect 8684 6273 8718 6307
rect 11069 6273 11103 6307
rect 13093 6273 13127 6307
rect 14197 6273 14231 6307
rect 2329 6205 2363 6239
rect 3065 6205 3099 6239
rect 4905 6205 4939 6239
rect 6837 6205 6871 6239
rect 10885 6205 10919 6239
rect 14841 6205 14875 6239
rect 3332 6137 3366 6171
rect 5172 6137 5206 6171
rect 7104 6137 7138 6171
rect 8922 6137 8956 6171
rect 12909 6137 12943 6171
rect 14013 6137 14047 6171
rect 2237 6069 2271 6103
rect 6285 6069 6319 6103
rect 8217 6069 8251 6103
rect 10977 6069 11011 6103
rect 11713 6069 11747 6103
rect 12817 6069 12851 6103
rect 13645 6069 13679 6103
rect 14105 6069 14139 6103
rect 15025 6069 15059 6103
rect 1593 5865 1627 5899
rect 2053 5865 2087 5899
rect 3157 5865 3191 5899
rect 8493 5865 8527 5899
rect 8953 5865 8987 5899
rect 12357 5865 12391 5899
rect 13553 5865 13587 5899
rect 14013 5865 14047 5899
rect 1961 5797 1995 5831
rect 4445 5729 4479 5763
rect 5540 5729 5574 5763
rect 7113 5729 7147 5763
rect 7369 5729 7403 5763
rect 9689 5729 9723 5763
rect 11529 5729 11563 5763
rect 12725 5729 12759 5763
rect 12817 5729 12851 5763
rect 13921 5729 13955 5763
rect 14933 5729 14967 5763
rect 2237 5661 2271 5695
rect 3249 5661 3283 5695
rect 3433 5661 3467 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 5273 5661 5307 5695
rect 10057 5661 10091 5695
rect 11621 5661 11655 5695
rect 11805 5661 11839 5695
rect 12909 5661 12943 5695
rect 14105 5661 14139 5695
rect 2789 5525 2823 5559
rect 4077 5525 4111 5559
rect 6653 5525 6687 5559
rect 11161 5525 11195 5559
rect 14749 5525 14783 5559
rect 4445 5321 4479 5355
rect 13645 5321 13679 5355
rect 8217 5253 8251 5287
rect 10057 5253 10091 5287
rect 12449 5253 12483 5287
rect 2513 5185 2547 5219
rect 3065 5185 3099 5219
rect 8677 5185 8711 5219
rect 11161 5185 11195 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 14197 5185 14231 5219
rect 3321 5117 3355 5151
rect 4905 5117 4939 5151
rect 6837 5117 6871 5151
rect 8933 5117 8967 5151
rect 10977 5117 11011 5151
rect 14013 5117 14047 5151
rect 14841 5117 14875 5151
rect 2237 5049 2271 5083
rect 5172 5049 5206 5083
rect 7104 5049 7138 5083
rect 10885 5049 10919 5083
rect 12817 5049 12851 5083
rect 1869 4981 1903 5015
rect 2329 4981 2363 5015
rect 6285 4981 6319 5015
rect 10517 4981 10551 5015
rect 11713 4981 11747 5015
rect 14105 4981 14139 5015
rect 15025 4981 15059 5015
rect 2053 4777 2087 4811
rect 8677 4777 8711 4811
rect 10057 4777 10091 4811
rect 12081 4777 12115 4811
rect 13277 4777 13311 4811
rect 13645 4777 13679 4811
rect 12449 4709 12483 4743
rect 12541 4709 12575 4743
rect 13737 4709 13771 4743
rect 1961 4641 1995 4675
rect 3157 4641 3191 4675
rect 3249 4641 3283 4675
rect 4629 4641 4663 4675
rect 4721 4641 4755 4675
rect 5457 4641 5491 4675
rect 5713 4641 5747 4675
rect 7564 4641 7598 4675
rect 9321 4641 9355 4675
rect 11253 4641 11287 4675
rect 11345 4641 11379 4675
rect 14473 4641 14507 4675
rect 2237 4573 2271 4607
rect 3433 4573 3467 4607
rect 4905 4573 4939 4607
rect 7297 4573 7331 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11437 4573 11471 4607
rect 12633 4573 12667 4607
rect 13829 4573 13863 4607
rect 1593 4505 1627 4539
rect 9689 4505 9723 4539
rect 10885 4505 10919 4539
rect 14657 4505 14691 4539
rect 2789 4437 2823 4471
rect 4261 4437 4295 4471
rect 6837 4437 6871 4471
rect 9137 4437 9171 4471
rect 8217 4233 8251 4267
rect 10057 4233 10091 4267
rect 10517 4233 10551 4267
rect 6285 4165 6319 4199
rect 2973 4097 3007 4131
rect 3157 4097 3191 4131
rect 4353 4097 4387 4131
rect 11069 4097 11103 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 14749 4097 14783 4131
rect 1593 4029 1627 4063
rect 4905 4029 4939 4063
rect 5172 4029 5206 4063
rect 6837 4029 6871 4063
rect 8677 4029 8711 4063
rect 13645 4029 13679 4063
rect 14565 4029 14599 4063
rect 1869 3961 1903 3995
rect 7082 3961 7116 3995
rect 8944 3961 8978 3995
rect 10885 3961 10919 3995
rect 13921 3961 13955 3995
rect 2513 3893 2547 3927
rect 2881 3893 2915 3927
rect 3709 3893 3743 3927
rect 4077 3893 4111 3927
rect 4169 3893 4203 3927
rect 10977 3893 11011 3927
rect 11713 3893 11747 3927
rect 12449 3893 12483 3927
rect 12817 3893 12851 3927
rect 2053 3689 2087 3723
rect 3157 3689 3191 3723
rect 3249 3689 3283 3723
rect 4537 3689 4571 3723
rect 8585 3689 8619 3723
rect 9045 3689 9079 3723
rect 11253 3689 11287 3723
rect 11345 3689 11379 3723
rect 13553 3621 13587 3655
rect 1961 3553 1995 3587
rect 4629 3553 4663 3587
rect 5365 3553 5399 3587
rect 5632 3553 5666 3587
rect 7461 3553 7495 3587
rect 9229 3553 9263 3587
rect 10057 3553 10091 3587
rect 12449 3553 12483 3587
rect 13277 3553 13311 3587
rect 14289 3553 14323 3587
rect 2237 3485 2271 3519
rect 3341 3485 3375 3519
rect 4813 3485 4847 3519
rect 7205 3485 7239 3519
rect 10149 3485 10183 3519
rect 10241 3485 10275 3519
rect 11437 3485 11471 3519
rect 12541 3485 12575 3519
rect 12633 3485 12667 3519
rect 14473 3485 14507 3519
rect 2789 3417 2823 3451
rect 9689 3417 9723 3451
rect 1593 3349 1627 3383
rect 4169 3349 4203 3383
rect 6745 3349 6779 3383
rect 10885 3349 10919 3383
rect 12081 3349 12115 3383
rect 2513 3145 2547 3179
rect 8217 3145 8251 3179
rect 8677 3145 8711 3179
rect 11069 3145 11103 3179
rect 3709 3077 3743 3111
rect 9873 3077 9907 3111
rect 12265 3077 12299 3111
rect 2973 3009 3007 3043
rect 3157 3009 3191 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 9229 3009 9263 3043
rect 10425 3009 10459 3043
rect 11621 3009 11655 3043
rect 1593 2941 1627 2975
rect 4905 2941 4939 2975
rect 5172 2941 5206 2975
rect 6837 2941 6871 2975
rect 9137 2941 9171 2975
rect 10333 2941 10367 2975
rect 13645 3009 13679 3043
rect 12449 2941 12483 2975
rect 13369 2941 13403 2975
rect 14289 2941 14323 2975
rect 1869 2873 1903 2907
rect 2881 2873 2915 2907
rect 7104 2873 7138 2907
rect 9045 2873 9079 2907
rect 12265 2873 12299 2907
rect 12725 2873 12759 2907
rect 14565 2873 14599 2907
rect 4077 2805 4111 2839
rect 6285 2805 6319 2839
rect 10241 2805 10275 2839
rect 11437 2805 11471 2839
rect 11529 2805 11563 2839
rect 4445 2601 4479 2635
rect 4905 2601 4939 2635
rect 5641 2601 5675 2635
rect 6101 2601 6135 2635
rect 6929 2601 6963 2635
rect 8125 2601 8159 2635
rect 10149 2601 10183 2635
rect 10241 2601 10275 2635
rect 10977 2601 11011 2635
rect 11437 2601 11471 2635
rect 4813 2533 4847 2567
rect 1409 2465 1443 2499
rect 2412 2465 2446 2499
rect 6009 2465 6043 2499
rect 7297 2465 7331 2499
rect 7389 2465 7423 2499
rect 8493 2465 8527 2499
rect 9505 2465 9539 2499
rect 11345 2465 11379 2499
rect 12357 2465 12391 2499
rect 12633 2465 12667 2499
rect 13921 2465 13955 2499
rect 2145 2397 2179 2431
rect 5089 2397 5123 2431
rect 6285 2397 6319 2431
rect 7481 2397 7515 2431
rect 8585 2397 8619 2431
rect 8769 2397 8803 2431
rect 10333 2397 10367 2431
rect 11529 2397 11563 2431
rect 12817 2397 12851 2431
rect 14197 2397 14231 2431
rect 3525 2329 3559 2363
rect 1593 2261 1627 2295
rect 9321 2261 9355 2295
rect 9781 2261 9815 2295
rect 12173 2261 12207 2295
rect 12357 1853 12391 1887
rect 12357 1445 12391 1479
<< metal1 >>
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 9398 18068 9404 18080
rect 4856 18040 9404 18068
rect 4856 18028 4862 18040
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 5166 17960 5172 18012
rect 5224 18000 5230 18012
rect 9490 18000 9496 18012
rect 5224 17972 9496 18000
rect 5224 17960 5230 17972
rect 9490 17960 9496 17972
rect 9548 17960 9554 18012
rect 7190 17892 7196 17944
rect 7248 17932 7254 17944
rect 12066 17932 12072 17944
rect 7248 17904 12072 17932
rect 7248 17892 7254 17904
rect 12066 17892 12072 17904
rect 12124 17892 12130 17944
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 9030 17864 9036 17876
rect 3568 17836 9036 17864
rect 3568 17824 3574 17836
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 5994 17756 6000 17808
rect 6052 17796 6058 17808
rect 11146 17796 11152 17808
rect 6052 17768 11152 17796
rect 6052 17756 6058 17768
rect 11146 17756 11152 17768
rect 11204 17756 11210 17808
rect 4522 17688 4528 17740
rect 4580 17728 4586 17740
rect 10226 17728 10232 17740
rect 4580 17700 10232 17728
rect 4580 17688 4586 17700
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 11330 17660 11336 17672
rect 6972 17632 11336 17660
rect 6972 17620 6978 17632
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 4154 17552 4160 17604
rect 4212 17592 4218 17604
rect 9858 17592 9864 17604
rect 4212 17564 9864 17592
rect 4212 17552 4218 17564
rect 9858 17552 9864 17564
rect 9916 17552 9922 17604
rect 10502 17552 10508 17604
rect 10560 17592 10566 17604
rect 12434 17592 12440 17604
rect 10560 17564 12440 17592
rect 10560 17552 10566 17564
rect 12434 17552 12440 17564
rect 12492 17552 12498 17604
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 10686 17524 10692 17536
rect 5592 17496 10692 17524
rect 5592 17484 5598 17496
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 11422 17484 11428 17536
rect 11480 17524 11486 17536
rect 16022 17524 16028 17536
rect 11480 17496 16028 17524
rect 11480 17484 11486 17496
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 3108 17292 5641 17320
rect 3108 17280 3114 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 5629 17283 5687 17289
rect 6178 17280 6184 17332
rect 6236 17280 6242 17332
rect 6914 17320 6920 17332
rect 6875 17292 6920 17320
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 10502 17320 10508 17332
rect 8076 17292 10508 17320
rect 8076 17280 8082 17292
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 10686 17320 10692 17332
rect 10647 17292 10692 17320
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 2130 17212 2136 17264
rect 2188 17252 2194 17264
rect 6196 17252 6224 17280
rect 11425 17255 11483 17261
rect 11425 17252 11437 17255
rect 2188 17224 3188 17252
rect 6196 17224 11437 17252
rect 2188 17212 2194 17224
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 2774 17184 2780 17196
rect 2363 17156 2780 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 3160 17193 3188 17224
rect 11425 17221 11437 17224
rect 11471 17221 11483 17255
rect 11425 17215 11483 17221
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 3234 17144 3240 17196
rect 3292 17184 3298 17196
rect 4249 17187 4307 17193
rect 4249 17184 4261 17187
rect 3292 17156 4261 17184
rect 3292 17144 3298 17156
rect 4249 17153 4261 17156
rect 4295 17153 4307 17187
rect 6270 17184 6276 17196
rect 6231 17156 6276 17184
rect 4249 17147 4307 17153
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 7466 17184 7472 17196
rect 7427 17156 7472 17184
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 8036 17156 8340 17184
rect 2051 17119 2109 17125
rect 2051 17085 2063 17119
rect 2097 17085 2109 17119
rect 2958 17116 2964 17128
rect 2871 17088 2964 17116
rect 2051 17079 2109 17085
rect 2056 17048 2084 17079
rect 2958 17076 2964 17088
rect 3016 17116 3022 17128
rect 3970 17116 3976 17128
rect 3016 17088 3976 17116
rect 3016 17076 3022 17088
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17085 4123 17119
rect 4065 17079 4123 17085
rect 4985 17119 5043 17125
rect 4985 17085 4997 17119
rect 5031 17116 5043 17119
rect 7098 17116 7104 17128
rect 5031 17088 7104 17116
rect 5031 17085 5043 17088
rect 4985 17079 5043 17085
rect 3878 17048 3884 17060
rect 2056 17020 3884 17048
rect 3878 17008 3884 17020
rect 3936 17048 3942 17060
rect 4080 17048 4108 17079
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 7248 17088 7297 17116
rect 7248 17076 7254 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 5994 17048 6000 17060
rect 3936 17020 4108 17048
rect 5955 17020 6000 17048
rect 3936 17008 3942 17020
rect 5994 17008 6000 17020
rect 6052 17008 6058 17060
rect 7374 17048 7380 17060
rect 7335 17020 7380 17048
rect 7374 17008 7380 17020
rect 7432 17048 7438 17060
rect 8036 17048 8064 17156
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8312 17116 8340 17156
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 12802 17184 12808 17196
rect 8444 17156 12808 17184
rect 8444 17144 8450 17156
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 8849 17119 8907 17125
rect 8849 17116 8861 17119
rect 8312 17088 8861 17116
rect 8113 17079 8171 17085
rect 8849 17085 8861 17088
rect 8895 17085 8907 17119
rect 9766 17116 9772 17128
rect 9727 17088 9772 17116
rect 8849 17079 8907 17085
rect 7432 17020 8064 17048
rect 8128 17048 8156 17079
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 10134 17076 10140 17128
rect 10192 17116 10198 17128
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 10192 17088 10517 17116
rect 10192 17076 10198 17088
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 11882 17116 11888 17128
rect 11287 17088 11888 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 11882 17076 11888 17088
rect 11940 17076 11946 17128
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12584 17088 12633 17116
rect 12584 17076 12590 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 8754 17048 8760 17060
rect 8128 17020 8760 17048
rect 7432 17008 7438 17020
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 9214 17008 9220 17060
rect 9272 17048 9278 17060
rect 13538 17048 13544 17060
rect 9272 17020 13544 17048
rect 9272 17008 9278 17020
rect 13538 17008 13544 17020
rect 13596 17008 13602 17060
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 7926 16980 7932 16992
rect 6135 16952 7932 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 7926 16940 7932 16952
rect 7984 16940 7990 16992
rect 8297 16983 8355 16989
rect 8297 16949 8309 16983
rect 8343 16980 8355 16983
rect 8662 16980 8668 16992
rect 8343 16952 8668 16980
rect 8343 16949 8355 16952
rect 8297 16943 8355 16949
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9732 16952 9965 16980
rect 9732 16940 9738 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 10560 16952 12817 16980
rect 10560 16940 10566 16952
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 12805 16943 12863 16949
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 4430 16736 4436 16788
rect 4488 16776 4494 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 4488 16748 5273 16776
rect 4488 16736 4494 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 5261 16739 5319 16745
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 5592 16748 7665 16776
rect 5592 16736 5598 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 7653 16739 7711 16745
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 11422 16776 11428 16788
rect 9364 16748 11428 16776
rect 9364 16736 9370 16748
rect 11422 16736 11428 16748
rect 11480 16736 11486 16788
rect 12066 16776 12072 16788
rect 12027 16748 12072 16776
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 13538 16776 13544 16788
rect 13499 16748 13544 16776
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 3326 16708 3332 16720
rect 1780 16680 3332 16708
rect 1780 16649 1808 16680
rect 3326 16668 3332 16680
rect 3384 16668 3390 16720
rect 5629 16711 5687 16717
rect 5629 16677 5641 16711
rect 5675 16708 5687 16711
rect 7834 16708 7840 16720
rect 5675 16680 7840 16708
rect 5675 16677 5687 16680
rect 5629 16671 5687 16677
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 8113 16711 8171 16717
rect 8113 16677 8125 16711
rect 8159 16708 8171 16711
rect 10042 16708 10048 16720
rect 8159 16680 10048 16708
rect 8159 16677 8171 16680
rect 8113 16671 8171 16677
rect 10042 16668 10048 16680
rect 10100 16708 10106 16720
rect 11238 16708 11244 16720
rect 10100 16680 11244 16708
rect 10100 16668 10106 16680
rect 11238 16668 11244 16680
rect 11296 16668 11302 16720
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16609 1823 16643
rect 1765 16603 1823 16609
rect 1946 16600 1952 16652
rect 2004 16640 2010 16652
rect 2041 16643 2099 16649
rect 2041 16640 2053 16643
rect 2004 16612 2053 16640
rect 2004 16600 2010 16612
rect 2041 16609 2053 16612
rect 2087 16609 2099 16643
rect 2041 16603 2099 16609
rect 2130 16600 2136 16652
rect 2188 16640 2194 16652
rect 2685 16643 2743 16649
rect 2685 16640 2697 16643
rect 2188 16612 2697 16640
rect 2188 16600 2194 16612
rect 2685 16609 2697 16612
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 4028 16612 4077 16640
rect 4028 16600 4034 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16640 5227 16643
rect 5350 16640 5356 16652
rect 5215 16612 5356 16640
rect 5215 16609 5227 16612
rect 5169 16603 5227 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5721 16643 5779 16649
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 6638 16640 6644 16652
rect 5767 16612 6644 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 6822 16640 6828 16652
rect 6783 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7742 16640 7748 16652
rect 7024 16612 7748 16640
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3142 16572 3148 16584
rect 3007 16544 3148 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 3292 16544 4261 16572
rect 3292 16532 3298 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 5828 16504 5856 16535
rect 5902 16532 5908 16584
rect 5960 16572 5966 16584
rect 6730 16572 6736 16584
rect 5960 16544 6736 16572
rect 5960 16532 5966 16544
rect 6730 16532 6736 16544
rect 6788 16532 6794 16584
rect 7024 16581 7052 16612
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 8386 16640 8392 16652
rect 8352 16612 8392 16640
rect 8352 16600 8358 16612
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 8855 16643 8913 16649
rect 8855 16609 8867 16643
rect 8901 16609 8913 16643
rect 8855 16603 8913 16609
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10318 16640 10324 16652
rect 9723 16612 10324 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 6917 16575 6975 16581
rect 6917 16541 6929 16575
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 6270 16504 6276 16516
rect 5828 16476 6276 16504
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 6932 16504 6960 16535
rect 8018 16532 8024 16584
rect 8076 16572 8082 16584
rect 8205 16575 8263 16581
rect 8205 16572 8217 16575
rect 8076 16544 8217 16572
rect 8076 16532 8082 16544
rect 8205 16541 8217 16544
rect 8251 16541 8263 16575
rect 8205 16535 8263 16541
rect 8570 16532 8576 16584
rect 8628 16572 8634 16584
rect 8864 16572 8892 16603
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 11149 16643 11207 16649
rect 10468 16612 10513 16640
rect 10468 16600 10474 16612
rect 11149 16609 11161 16643
rect 11195 16640 11207 16643
rect 11790 16640 11796 16652
rect 11195 16612 11796 16640
rect 11195 16609 11207 16612
rect 11149 16603 11207 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12066 16640 12072 16652
rect 11931 16612 12072 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 12066 16600 12072 16612
rect 12124 16600 12130 16652
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12400 16612 12633 16640
rect 12400 16600 12406 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 12710 16600 12716 16652
rect 12768 16640 12774 16652
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 12768 16612 13369 16640
rect 12768 16600 12774 16612
rect 13357 16609 13369 16612
rect 13403 16609 13415 16643
rect 13357 16603 13415 16609
rect 8628 16544 8892 16572
rect 8628 16532 8634 16544
rect 9122 16532 9128 16584
rect 9180 16572 9186 16584
rect 10502 16572 10508 16584
rect 9180 16544 10508 16572
rect 9180 16532 9186 16544
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 7650 16504 7656 16516
rect 6932 16476 7656 16504
rect 7650 16464 7656 16476
rect 7708 16464 7714 16516
rect 9030 16504 9036 16516
rect 8991 16476 9036 16504
rect 9030 16464 9036 16476
rect 9088 16464 9094 16516
rect 9398 16464 9404 16516
rect 9456 16504 9462 16516
rect 9674 16504 9680 16516
rect 9456 16476 9680 16504
rect 9456 16464 9462 16476
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 11333 16507 11391 16513
rect 11333 16504 11345 16507
rect 9784 16476 11345 16504
rect 4985 16439 5043 16445
rect 4985 16405 4997 16439
rect 5031 16436 5043 16439
rect 5442 16436 5448 16448
rect 5031 16408 5448 16436
rect 5031 16405 5043 16408
rect 4985 16399 5043 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6454 16436 6460 16448
rect 6415 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 6730 16396 6736 16448
rect 6788 16436 6794 16448
rect 9784 16436 9812 16476
rect 11333 16473 11345 16476
rect 11379 16473 11391 16507
rect 11333 16467 11391 16473
rect 6788 16408 9812 16436
rect 6788 16396 6794 16408
rect 9858 16396 9864 16448
rect 9916 16436 9922 16448
rect 9916 16408 9961 16436
rect 9916 16396 9922 16408
rect 10226 16396 10232 16448
rect 10284 16436 10290 16448
rect 10597 16439 10655 16445
rect 10597 16436 10609 16439
rect 10284 16408 10609 16436
rect 10284 16396 10290 16408
rect 10597 16405 10609 16408
rect 10643 16405 10655 16439
rect 10597 16399 10655 16405
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 3326 16192 3332 16244
rect 3384 16232 3390 16244
rect 3973 16235 4031 16241
rect 3973 16232 3985 16235
rect 3384 16204 3985 16232
rect 3384 16192 3390 16204
rect 3973 16201 3985 16204
rect 4019 16201 4031 16235
rect 3973 16195 4031 16201
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 6880 16204 8033 16232
rect 6880 16192 6886 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 8128 16204 9444 16232
rect 4246 16124 4252 16176
rect 4304 16164 4310 16176
rect 8128 16164 8156 16204
rect 9217 16167 9275 16173
rect 9217 16164 9229 16167
rect 4304 16136 8156 16164
rect 8220 16136 9229 16164
rect 4304 16124 4310 16136
rect 4614 16096 4620 16108
rect 4575 16068 4620 16096
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 5718 16096 5724 16108
rect 5679 16068 5724 16096
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 6972 16068 7389 16096
rect 6972 16056 6978 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 8220 16096 8248 16136
rect 9217 16133 9229 16136
rect 9263 16133 9275 16167
rect 9416 16164 9444 16204
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 10008 16204 14105 16232
rect 10008 16192 10014 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 10597 16167 10655 16173
rect 10597 16164 10609 16167
rect 9416 16136 10609 16164
rect 9217 16127 9275 16133
rect 10597 16133 10609 16136
rect 10643 16133 10655 16167
rect 10597 16127 10655 16133
rect 10778 16124 10784 16176
rect 10836 16164 10842 16176
rect 11333 16167 11391 16173
rect 11333 16164 11345 16167
rect 10836 16136 11345 16164
rect 10836 16124 10842 16136
rect 11333 16133 11345 16136
rect 11379 16133 11391 16167
rect 12618 16164 12624 16176
rect 12579 16136 12624 16164
rect 11333 16127 11391 16133
rect 12618 16124 12624 16136
rect 12676 16124 12682 16176
rect 7892 16068 8248 16096
rect 8665 16099 8723 16105
rect 7892 16056 7898 16068
rect 8665 16065 8677 16099
rect 8711 16096 8723 16099
rect 8846 16096 8852 16108
rect 8711 16068 8852 16096
rect 8711 16065 8723 16068
rect 8665 16059 8723 16065
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 9769 16099 9827 16105
rect 9769 16096 9781 16099
rect 9232 16068 9781 16096
rect 9232 16040 9260 16068
rect 9769 16065 9781 16068
rect 9815 16065 9827 16099
rect 10870 16096 10876 16108
rect 9769 16059 9827 16065
rect 9876 16068 10876 16096
rect 9876 16040 9904 16068
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2682 16028 2688 16040
rect 2643 16000 2688 16028
rect 2682 15988 2688 16000
rect 2740 15988 2746 16040
rect 4338 16028 4344 16040
rect 4299 16000 4344 16028
rect 4338 15988 4344 16000
rect 4396 15988 4402 16040
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 16028 5595 16031
rect 6454 16028 6460 16040
rect 5583 16000 6460 16028
rect 5583 15997 5595 16000
rect 5537 15991 5595 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 8294 16028 8300 16040
rect 6687 16000 8300 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8478 16028 8484 16040
rect 8439 16000 8484 16028
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 9214 15988 9220 16040
rect 9272 15988 9278 16040
rect 9306 15988 9312 16040
rect 9364 16028 9370 16040
rect 9585 16031 9643 16037
rect 9585 16028 9597 16031
rect 9364 16000 9597 16028
rect 9364 15988 9370 16000
rect 9585 15997 9597 16000
rect 9631 15997 9643 16031
rect 9585 15991 9643 15997
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 9858 16028 9864 16040
rect 9723 16000 9864 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 9858 15988 9864 16000
rect 9916 15988 9922 16040
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 10502 16028 10508 16040
rect 10459 16000 10508 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11238 16028 11244 16040
rect 11195 16000 11244 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 12434 16028 12440 16040
rect 12395 16000 12440 16028
rect 12434 15988 12440 16000
rect 12492 15988 12498 16040
rect 12894 15988 12900 16040
rect 12952 16028 12958 16040
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 12952 16000 13185 16028
rect 12952 15988 12958 16000
rect 13173 15997 13185 16000
rect 13219 15997 13231 16031
rect 13906 16028 13912 16040
rect 13867 16000 13912 16028
rect 13173 15991 13231 15997
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 2038 15960 2044 15972
rect 1999 15932 2044 15960
rect 2038 15920 2044 15932
rect 2096 15920 2102 15972
rect 2958 15960 2964 15972
rect 2919 15932 2964 15960
rect 2958 15920 2964 15932
rect 3016 15920 3022 15972
rect 3878 15920 3884 15972
rect 3936 15960 3942 15972
rect 4433 15963 4491 15969
rect 4433 15960 4445 15963
rect 3936 15932 4445 15960
rect 3936 15920 3942 15932
rect 4433 15929 4445 15932
rect 4479 15929 4491 15963
rect 5629 15963 5687 15969
rect 5629 15960 5641 15963
rect 4433 15923 4491 15929
rect 4540 15932 5641 15960
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 2314 15892 2320 15904
rect 1452 15864 2320 15892
rect 1452 15852 1458 15864
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 4540 15892 4568 15932
rect 5629 15929 5641 15932
rect 5675 15929 5687 15963
rect 8389 15963 8447 15969
rect 5629 15923 5687 15929
rect 6840 15932 8248 15960
rect 5166 15892 5172 15904
rect 4212 15864 4568 15892
rect 5127 15864 5172 15892
rect 4212 15852 4218 15864
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6840 15901 6868 15932
rect 6457 15895 6515 15901
rect 6457 15892 6469 15895
rect 6420 15864 6469 15892
rect 6420 15852 6426 15864
rect 6457 15861 6469 15864
rect 6503 15861 6515 15895
rect 6457 15855 6515 15861
rect 6825 15895 6883 15901
rect 6825 15861 6837 15895
rect 6871 15861 6883 15895
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 6825 15855 6883 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7374 15892 7380 15904
rect 7331 15864 7380 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 8220 15892 8248 15932
rect 8389 15929 8401 15963
rect 8435 15960 8447 15963
rect 8435 15932 9812 15960
rect 8435 15929 8447 15932
rect 8389 15923 8447 15929
rect 9398 15892 9404 15904
rect 8220 15864 9404 15892
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 9674 15892 9680 15904
rect 9548 15864 9680 15892
rect 9548 15852 9554 15864
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 9784 15892 9812 15932
rect 9858 15892 9864 15904
rect 9784 15864 9864 15892
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 11572 15864 13369 15892
rect 11572 15852 11578 15864
rect 13357 15861 13369 15864
rect 13403 15861 13415 15895
rect 13357 15855 13415 15861
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 1670 15648 1676 15700
rect 1728 15648 1734 15700
rect 4709 15691 4767 15697
rect 4709 15657 4721 15691
rect 4755 15688 4767 15691
rect 5534 15688 5540 15700
rect 4755 15660 5540 15688
rect 4755 15657 4767 15660
rect 4709 15651 4767 15657
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 6917 15691 6975 15697
rect 6917 15657 6929 15691
rect 6963 15688 6975 15691
rect 7466 15688 7472 15700
rect 6963 15660 7472 15688
rect 6963 15657 6975 15660
rect 6917 15651 6975 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 8110 15648 8116 15700
rect 8168 15688 8174 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8168 15660 9321 15688
rect 8168 15648 8174 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 9309 15651 9367 15657
rect 9968 15660 13277 15688
rect 1688 15620 1716 15648
rect 1949 15623 2007 15629
rect 1949 15620 1961 15623
rect 1688 15592 1961 15620
rect 1949 15589 1961 15592
rect 1995 15589 2007 15623
rect 5166 15620 5172 15632
rect 1949 15583 2007 15589
rect 2608 15592 5172 15620
rect 2608 15561 2636 15592
rect 5166 15580 5172 15592
rect 5224 15580 5230 15632
rect 7837 15623 7895 15629
rect 7837 15589 7849 15623
rect 7883 15620 7895 15623
rect 8754 15620 8760 15632
rect 7883 15592 8760 15620
rect 7883 15589 7895 15592
rect 7837 15583 7895 15589
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 9968 15620 9996 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 9640 15592 9996 15620
rect 10045 15623 10103 15629
rect 9640 15580 9646 15592
rect 10045 15589 10057 15623
rect 10091 15620 10103 15623
rect 13630 15620 13636 15632
rect 10091 15592 13636 15620
rect 10091 15589 10103 15592
rect 10045 15583 10103 15589
rect 13630 15580 13636 15592
rect 13688 15580 13694 15632
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15521 1731 15555
rect 1673 15515 1731 15521
rect 2603 15555 2661 15561
rect 2603 15521 2615 15555
rect 2649 15521 2661 15555
rect 2603 15515 2661 15521
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15552 3939 15555
rect 5350 15552 5356 15564
rect 3927 15524 5356 15552
rect 3927 15521 3939 15524
rect 3881 15515 3939 15521
rect 1688 15416 1716 15515
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 5810 15561 5816 15564
rect 5537 15555 5595 15561
rect 5537 15552 5549 15555
rect 5500 15524 5549 15552
rect 5500 15512 5506 15524
rect 5537 15521 5549 15524
rect 5583 15521 5595 15555
rect 5804 15552 5816 15561
rect 5771 15524 5816 15552
rect 5537 15515 5595 15521
rect 5804 15515 5816 15524
rect 5810 15512 5816 15515
rect 5868 15512 5874 15564
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15552 7803 15555
rect 8202 15552 8208 15564
rect 7791 15524 8208 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8570 15552 8576 15564
rect 8531 15524 8576 15552
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 9490 15552 9496 15564
rect 9451 15524 9496 15552
rect 9490 15512 9496 15524
rect 9548 15512 9554 15564
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10686 15552 10692 15564
rect 10183 15524 10692 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 11422 15552 11428 15564
rect 10919 15524 11428 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 11609 15555 11667 15561
rect 11609 15521 11621 15555
rect 11655 15552 11667 15555
rect 11698 15552 11704 15564
rect 11655 15524 11704 15552
rect 11655 15521 11667 15524
rect 11609 15515 11667 15521
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 12216 15524 12357 15552
rect 12216 15512 12222 15524
rect 12345 15521 12357 15524
rect 12391 15521 12403 15555
rect 13078 15552 13084 15564
rect 13039 15524 13084 15552
rect 12345 15515 12403 15521
rect 13078 15512 13084 15524
rect 13136 15512 13142 15564
rect 2866 15484 2872 15496
rect 2827 15456 2872 15484
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 3844 15456 4813 15484
rect 3844 15444 3850 15456
rect 4801 15453 4813 15456
rect 4847 15453 4859 15487
rect 4982 15484 4988 15496
rect 4943 15456 4988 15484
rect 4801 15447 4859 15453
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 7926 15484 7932 15496
rect 7887 15456 7932 15484
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 9508 15484 9536 15512
rect 8352 15456 9536 15484
rect 8352 15444 8358 15456
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 10008 15456 10241 15484
rect 10008 15444 10014 15456
rect 10229 15453 10241 15456
rect 10275 15484 10287 15487
rect 10502 15484 10508 15496
rect 10275 15456 10508 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 10962 15444 10968 15496
rect 11020 15484 11026 15496
rect 11020 15456 11100 15484
rect 11020 15444 11026 15456
rect 3234 15416 3240 15428
rect 1688 15388 3240 15416
rect 3234 15376 3240 15388
rect 3292 15376 3298 15428
rect 8757 15419 8815 15425
rect 8757 15385 8769 15419
rect 8803 15416 8815 15419
rect 8938 15416 8944 15428
rect 8803 15388 8944 15416
rect 8803 15385 8815 15388
rect 8757 15379 8815 15385
rect 8938 15376 8944 15388
rect 8996 15376 9002 15428
rect 9122 15376 9128 15428
rect 9180 15416 9186 15428
rect 11072 15425 11100 15456
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11330 15484 11336 15496
rect 11204 15456 11336 15484
rect 11204 15444 11210 15456
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 9677 15419 9735 15425
rect 9677 15416 9689 15419
rect 9180 15388 9689 15416
rect 9180 15376 9186 15388
rect 9677 15385 9689 15388
rect 9723 15385 9735 15419
rect 9677 15379 9735 15385
rect 11057 15419 11115 15425
rect 11057 15385 11069 15419
rect 11103 15385 11115 15419
rect 11057 15379 11115 15385
rect 11793 15419 11851 15425
rect 11793 15385 11805 15419
rect 11839 15416 11851 15419
rect 12066 15416 12072 15428
rect 11839 15388 12072 15416
rect 11839 15385 11851 15388
rect 11793 15379 11851 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 15378 15416 15384 15428
rect 12308 15388 15384 15416
rect 12308 15376 12314 15388
rect 15378 15376 15384 15388
rect 15436 15376 15442 15428
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3697 15351 3755 15357
rect 3697 15348 3709 15351
rect 2832 15320 3709 15348
rect 2832 15308 2838 15320
rect 3697 15317 3709 15320
rect 3743 15317 3755 15351
rect 4338 15348 4344 15360
rect 4299 15320 4344 15348
rect 3697 15311 3755 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 6546 15348 6552 15360
rect 5408 15320 6552 15348
rect 5408 15308 5414 15320
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 7374 15348 7380 15360
rect 7335 15320 7380 15348
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 12529 15351 12587 15357
rect 12529 15348 12541 15351
rect 7616 15320 12541 15348
rect 7616 15308 7622 15320
rect 12529 15317 12541 15320
rect 12575 15317 12587 15351
rect 12529 15311 12587 15317
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 16758 15348 16764 15360
rect 12676 15320 16764 15348
rect 12676 15308 12682 15320
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2682 15144 2688 15156
rect 2547 15116 2688 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 3697 15147 3755 15153
rect 3697 15113 3709 15147
rect 3743 15144 3755 15147
rect 3786 15144 3792 15156
rect 3743 15116 3792 15144
rect 3743 15113 3755 15116
rect 3697 15107 3755 15113
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 8665 15147 8723 15153
rect 4172 15116 7779 15144
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 3418 15076 3424 15088
rect 3292 15048 3424 15076
rect 3292 15036 3298 15048
rect 3418 15036 3424 15048
rect 3476 15036 3482 15088
rect 2590 14968 2596 15020
rect 2648 15008 2654 15020
rect 3053 15011 3111 15017
rect 3053 15008 3065 15011
rect 2648 14980 3065 15008
rect 2648 14968 2654 14980
rect 3053 14977 3065 14980
rect 3099 14977 3111 15011
rect 3053 14971 3111 14977
rect 3786 14968 3792 15020
rect 3844 15008 3850 15020
rect 4062 15008 4068 15020
rect 3844 14980 4068 15008
rect 3844 14968 3850 14980
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4172 15017 4200 15116
rect 7751 15076 7779 15116
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 8754 15144 8760 15156
rect 8711 15116 8760 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 9332 15116 9873 15144
rect 9332 15076 9360 15116
rect 9861 15113 9873 15116
rect 9907 15113 9919 15147
rect 11054 15144 11060 15156
rect 11015 15116 11060 15144
rect 9861 15107 9919 15113
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 12253 15147 12311 15153
rect 12253 15144 12265 15147
rect 11256 15116 12265 15144
rect 11256 15076 11284 15116
rect 12253 15113 12265 15116
rect 12299 15113 12311 15147
rect 12253 15107 12311 15113
rect 12621 15147 12679 15153
rect 12621 15113 12633 15147
rect 12667 15113 12679 15147
rect 12621 15107 12679 15113
rect 7751 15048 9360 15076
rect 9692 15048 11284 15076
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4798 15008 4804 15020
rect 4387 14980 4804 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 8570 14968 8576 15020
rect 8628 15008 8634 15020
rect 9122 15008 9128 15020
rect 8628 14980 9128 15008
rect 8628 14968 8634 14980
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9306 15008 9312 15020
rect 9267 14980 9312 15008
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 1578 14940 1584 14952
rect 1539 14912 1584 14940
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 2961 14943 3019 14949
rect 2961 14909 2973 14943
rect 3007 14940 3019 14943
rect 4430 14940 4436 14952
rect 3007 14912 4436 14940
rect 3007 14909 3019 14912
rect 2961 14903 3019 14909
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 4890 14940 4896 14952
rect 4803 14912 4896 14940
rect 4890 14900 4896 14912
rect 4948 14940 4954 14952
rect 5442 14940 5448 14952
rect 4948 14912 5448 14940
rect 4948 14900 4954 14912
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 6914 14940 6920 14952
rect 6871 14912 6920 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 7092 14943 7150 14949
rect 7092 14909 7104 14943
rect 7138 14940 7150 14943
rect 7466 14940 7472 14952
rect 7138 14912 7472 14940
rect 7138 14909 7150 14912
rect 7092 14903 7150 14909
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 9692 14940 9720 15048
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 9824 14980 10425 15008
rect 9824 14968 9830 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 9079 14912 9720 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 11256 14940 11284 15048
rect 11330 15036 11336 15088
rect 11388 15076 11394 15088
rect 12636 15076 12664 15107
rect 12802 15076 12808 15088
rect 11388 15048 12204 15076
rect 12636 15048 12808 15076
rect 11388 15036 11394 15048
rect 11514 15008 11520 15020
rect 11475 14980 11520 15008
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 11609 15011 11667 15017
rect 11609 14977 11621 15011
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 11422 14940 11428 14952
rect 10376 14912 10421 14940
rect 11256 14912 11428 14940
rect 10376 14900 10382 14912
rect 11422 14900 11428 14912
rect 11480 14900 11486 14952
rect 11624 14940 11652 14971
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 12066 15008 12072 15020
rect 11848 14980 12072 15008
rect 11848 14968 11854 14980
rect 12066 14968 12072 14980
rect 12124 14968 12130 15020
rect 12176 15008 12204 15048
rect 12802 15036 12808 15048
rect 12860 15036 12866 15088
rect 13170 15008 13176 15020
rect 12176 14980 13176 15008
rect 13170 14968 13176 14980
rect 13228 15008 13234 15020
rect 14550 15008 14556 15020
rect 13228 14980 14556 15008
rect 13228 14968 13234 14980
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 11532 14912 11652 14940
rect 12253 14943 12311 14949
rect 11532 14884 11560 14912
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12299 14912 12449 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 12802 14940 12808 14952
rect 12676 14912 12808 14940
rect 12676 14900 12682 14912
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 1854 14872 1860 14884
rect 1815 14844 1860 14872
rect 1854 14832 1860 14844
rect 1912 14832 1918 14884
rect 2869 14875 2927 14881
rect 2869 14841 2881 14875
rect 2915 14872 2927 14875
rect 3050 14872 3056 14884
rect 2915 14844 3056 14872
rect 2915 14841 2927 14844
rect 2869 14835 2927 14841
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 4982 14832 4988 14884
rect 5040 14872 5046 14884
rect 5160 14875 5218 14881
rect 5160 14872 5172 14875
rect 5040 14844 5172 14872
rect 5040 14832 5046 14844
rect 5160 14841 5172 14844
rect 5206 14872 5218 14875
rect 8478 14872 8484 14884
rect 5206 14844 8484 14872
rect 5206 14841 5218 14844
rect 5160 14835 5218 14841
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 8754 14872 8760 14884
rect 8588 14844 8760 14872
rect 4065 14807 4123 14813
rect 4065 14773 4077 14807
rect 4111 14804 4123 14807
rect 4246 14804 4252 14816
rect 4111 14776 4252 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 5810 14804 5816 14816
rect 4488 14776 5816 14804
rect 4488 14764 4494 14776
rect 5810 14764 5816 14776
rect 5868 14804 5874 14816
rect 6273 14807 6331 14813
rect 6273 14804 6285 14807
rect 5868 14776 6285 14804
rect 5868 14764 5874 14776
rect 6273 14773 6285 14776
rect 6319 14773 6331 14807
rect 6273 14767 6331 14773
rect 8205 14807 8263 14813
rect 8205 14773 8217 14807
rect 8251 14804 8263 14807
rect 8588 14804 8616 14844
rect 8754 14832 8760 14844
rect 8812 14872 8818 14884
rect 9214 14872 9220 14884
rect 8812 14844 9220 14872
rect 8812 14832 8818 14844
rect 9214 14832 9220 14844
rect 9272 14872 9278 14884
rect 11514 14872 11520 14884
rect 9272 14844 11520 14872
rect 9272 14832 9278 14844
rect 11514 14832 11520 14844
rect 11572 14832 11578 14884
rect 14458 14872 14464 14884
rect 11716 14844 14464 14872
rect 8251 14776 8616 14804
rect 9125 14807 9183 14813
rect 8251 14773 8263 14776
rect 8205 14767 8263 14773
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9582 14804 9588 14816
rect 9171 14776 9588 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 10229 14807 10287 14813
rect 10229 14773 10241 14807
rect 10275 14804 10287 14807
rect 10594 14804 10600 14816
rect 10275 14776 10600 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 11425 14807 11483 14813
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 11716 14804 11744 14844
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 11471 14776 11744 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13173 14807 13231 14813
rect 13173 14804 13185 14807
rect 12676 14776 13185 14804
rect 12676 14764 12682 14776
rect 13173 14773 13185 14776
rect 13219 14773 13231 14807
rect 13173 14767 13231 14773
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 9122 14600 9128 14612
rect 3283 14572 8984 14600
rect 9083 14572 9128 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3145 14535 3203 14541
rect 3145 14501 3157 14535
rect 3191 14532 3203 14535
rect 8570 14532 8576 14544
rect 3191 14504 8576 14532
rect 3191 14501 3203 14504
rect 3145 14495 3203 14501
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 8956 14532 8984 14572
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 9232 14572 10885 14600
rect 9232 14532 9260 14572
rect 10873 14569 10885 14572
rect 10919 14569 10931 14603
rect 10873 14563 10931 14569
rect 11241 14603 11299 14609
rect 11241 14569 11253 14603
rect 11287 14600 11299 14603
rect 11790 14600 11796 14612
rect 11287 14572 11796 14600
rect 11287 14569 11299 14572
rect 11241 14563 11299 14569
rect 11790 14560 11796 14572
rect 11848 14600 11854 14612
rect 12710 14600 12716 14612
rect 11848 14572 12716 14600
rect 11848 14560 11854 14572
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 9766 14532 9772 14544
rect 8956 14504 9260 14532
rect 9600 14504 9772 14532
rect 9600 14476 9628 14504
rect 9766 14492 9772 14504
rect 9824 14492 9830 14544
rect 10134 14532 10140 14544
rect 10095 14504 10140 14532
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14464 1915 14467
rect 3050 14464 3056 14476
rect 1903 14436 3056 14464
rect 1903 14433 1915 14436
rect 1857 14427 1915 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 4430 14464 4436 14476
rect 3344 14436 4436 14464
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2866 14396 2872 14408
rect 2179 14368 2872 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 2498 14288 2504 14340
rect 2556 14328 2562 14340
rect 3344 14328 3372 14436
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 5258 14464 5264 14476
rect 4663 14436 5264 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5442 14464 5448 14476
rect 5403 14436 5448 14464
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5534 14424 5540 14476
rect 5592 14424 5598 14476
rect 5712 14467 5770 14473
rect 5712 14433 5724 14467
rect 5758 14464 5770 14467
rect 5994 14464 6000 14476
rect 5758 14436 6000 14464
rect 5758 14433 5770 14436
rect 5712 14427 5770 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 7541 14467 7599 14473
rect 7541 14464 7553 14467
rect 6880 14436 7553 14464
rect 6880 14424 6886 14436
rect 7541 14433 7553 14436
rect 7587 14433 7599 14467
rect 7541 14427 7599 14433
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 8018 14464 8024 14476
rect 7892 14436 8024 14464
rect 7892 14424 7898 14436
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9309 14467 9367 14473
rect 9309 14464 9321 14467
rect 9272 14436 9321 14464
rect 9272 14424 9278 14436
rect 9309 14433 9321 14436
rect 9355 14433 9367 14467
rect 9309 14427 9367 14433
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9732 14436 10057 14464
rect 9732 14424 9738 14436
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 10502 14424 10508 14476
rect 10560 14464 10566 14476
rect 12069 14467 12127 14473
rect 10560 14436 11468 14464
rect 10560 14424 10566 14436
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 2556 14300 3372 14328
rect 3436 14328 3464 14359
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4580 14368 4721 14396
rect 4580 14356 4586 14368
rect 4709 14365 4721 14368
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5552 14396 5580 14424
rect 4939 14368 5580 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 6972 14368 7297 14396
rect 6972 14356 6978 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 9766 14396 9772 14408
rect 8352 14368 9772 14396
rect 8352 14356 8358 14368
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 9858 14356 9864 14408
rect 9916 14396 9922 14408
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 9916 14368 10241 14396
rect 9916 14356 9922 14368
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 11330 14396 11336 14408
rect 11291 14368 11336 14396
rect 10229 14359 10287 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11440 14405 11468 14436
rect 12069 14433 12081 14467
rect 12115 14464 12127 14467
rect 12250 14464 12256 14476
rect 12115 14436 12256 14464
rect 12115 14433 12127 14436
rect 12069 14427 12127 14433
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 12802 14464 12808 14476
rect 12763 14436 12808 14464
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 14274 14464 14280 14476
rect 13044 14436 14280 14464
rect 13044 14424 13050 14436
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 11425 14399 11483 14405
rect 11425 14365 11437 14399
rect 11471 14365 11483 14399
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 11425 14359 11483 14365
rect 12820 14368 13553 14396
rect 12820 14340 12848 14368
rect 13541 14365 13553 14368
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 14185 14399 14243 14405
rect 14185 14396 14197 14399
rect 14148 14368 14197 14396
rect 14148 14356 14154 14368
rect 14185 14365 14197 14368
rect 14231 14365 14243 14399
rect 14185 14359 14243 14365
rect 4982 14328 4988 14340
rect 3436 14300 4988 14328
rect 2556 14288 2562 14300
rect 4982 14288 4988 14300
rect 5040 14288 5046 14340
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 5442 14328 5448 14340
rect 5132 14300 5448 14328
rect 5132 14288 5138 14300
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 6656 14300 6960 14328
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 4249 14263 4307 14269
rect 2832 14232 2877 14260
rect 2832 14220 2838 14232
rect 4249 14229 4261 14263
rect 4295 14260 4307 14263
rect 6656 14260 6684 14300
rect 4295 14232 6684 14260
rect 4295 14229 4307 14232
rect 4249 14223 4307 14229
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 6825 14263 6883 14269
rect 6825 14260 6837 14263
rect 6788 14232 6837 14260
rect 6788 14220 6794 14232
rect 6825 14229 6837 14232
rect 6871 14229 6883 14263
rect 6932 14260 6960 14300
rect 8478 14288 8484 14340
rect 8536 14328 8542 14340
rect 8665 14331 8723 14337
rect 8665 14328 8677 14331
rect 8536 14300 8677 14328
rect 8536 14288 8542 14300
rect 8665 14297 8677 14300
rect 8711 14297 8723 14331
rect 8665 14291 8723 14297
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14328 9735 14331
rect 9723 14300 12756 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 10502 14260 10508 14272
rect 6932 14232 10508 14260
rect 6825 14223 6883 14229
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 12253 14263 12311 14269
rect 12253 14260 12265 14263
rect 11020 14232 12265 14260
rect 11020 14220 11026 14232
rect 12253 14229 12265 14232
rect 12299 14229 12311 14263
rect 12728 14260 12756 14300
rect 12802 14288 12808 14340
rect 12860 14288 12866 14340
rect 12986 14328 12992 14340
rect 12947 14300 12992 14328
rect 12986 14288 12992 14300
rect 13044 14288 13050 14340
rect 13170 14260 13176 14272
rect 12728 14232 13176 14260
rect 12253 14223 12311 14229
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1636 14028 1869 14056
rect 1636 14016 1642 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 1857 14019 1915 14025
rect 2590 14016 2596 14068
rect 2648 14056 2654 14068
rect 4433 14059 4491 14065
rect 4433 14056 4445 14059
rect 2648 14028 4445 14056
rect 2648 14016 2654 14028
rect 4433 14025 4445 14028
rect 4479 14056 4491 14059
rect 6273 14059 6331 14065
rect 4479 14028 5847 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 5819 13988 5847 14028
rect 6273 14025 6285 14059
rect 6319 14056 6331 14059
rect 9306 14056 9312 14068
rect 6319 14028 9312 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 9306 14016 9312 14028
rect 9364 14056 9370 14068
rect 9582 14056 9588 14068
rect 9364 14028 9588 14056
rect 9364 14016 9370 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9824 14028 10057 14056
rect 9824 14016 9830 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 10410 14016 10416 14068
rect 10468 14056 10474 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 10468 14028 10517 14056
rect 10468 14016 10474 14028
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 10505 14019 10563 14025
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 11112 14028 12449 14056
rect 11112 14016 11118 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 12437 14019 12495 14025
rect 6822 13988 6828 14000
rect 5819 13960 6828 13988
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 8205 13991 8263 13997
rect 8205 13988 8217 13991
rect 7892 13960 8217 13988
rect 7892 13948 7898 13960
rect 8205 13957 8217 13960
rect 8251 13988 8263 13991
rect 8294 13988 8300 14000
rect 8251 13960 8300 13988
rect 8251 13957 8263 13960
rect 8205 13951 8263 13957
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 10594 13948 10600 14000
rect 10652 13988 10658 14000
rect 10962 13988 10968 14000
rect 10652 13960 10968 13988
rect 10652 13948 10658 13960
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 2498 13920 2504 13932
rect 2459 13892 2504 13920
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 4890 13920 4896 13932
rect 4851 13892 4896 13920
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8665 13923 8723 13929
rect 8665 13920 8677 13923
rect 8168 13892 8677 13920
rect 8168 13880 8174 13892
rect 8665 13889 8677 13892
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 3053 13855 3111 13861
rect 2096 13824 3004 13852
rect 2096 13812 2102 13824
rect 2225 13787 2283 13793
rect 2225 13753 2237 13787
rect 2271 13784 2283 13787
rect 2774 13784 2780 13796
rect 2271 13756 2780 13784
rect 2271 13753 2283 13756
rect 2225 13747 2283 13753
rect 2774 13744 2780 13756
rect 2832 13744 2838 13796
rect 2976 13784 3004 13824
rect 3053 13821 3065 13855
rect 3099 13852 3111 13855
rect 4908 13852 4936 13880
rect 3099 13824 4936 13852
rect 5160 13855 5218 13861
rect 3099 13821 3111 13824
rect 3053 13815 3111 13821
rect 5160 13821 5172 13855
rect 5206 13852 5218 13855
rect 5718 13852 5724 13864
rect 5206 13824 5724 13852
rect 5206 13821 5218 13824
rect 5160 13815 5218 13821
rect 5718 13812 5724 13824
rect 5776 13852 5782 13864
rect 6730 13852 6736 13864
rect 5776 13824 6736 13852
rect 5776 13812 5782 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13852 6883 13855
rect 6914 13852 6920 13864
rect 6871 13824 6920 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 6914 13812 6920 13824
rect 6972 13852 6978 13864
rect 7466 13852 7472 13864
rect 6972 13824 7472 13852
rect 6972 13812 6978 13824
rect 7466 13812 7472 13824
rect 7524 13852 7530 13864
rect 8128 13852 8156 13880
rect 7524 13824 8156 13852
rect 7524 13812 7530 13824
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 9858 13852 9864 13864
rect 8352 13824 9864 13852
rect 8352 13812 8358 13824
rect 9858 13812 9864 13824
rect 9916 13852 9922 13864
rect 11164 13852 11192 13883
rect 11514 13880 11520 13932
rect 11572 13920 11578 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 11572 13892 13093 13920
rect 11572 13880 11578 13892
rect 13081 13889 13093 13892
rect 13127 13920 13139 13923
rect 13814 13920 13820 13932
rect 13127 13892 13820 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 12710 13852 12716 13864
rect 9916 13824 12716 13852
rect 9916 13812 9922 13824
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14240 13824 14657 13852
rect 14240 13812 14246 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14918 13852 14924 13864
rect 14879 13824 14924 13852
rect 14645 13815 14703 13821
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 3142 13784 3148 13796
rect 2976 13756 3148 13784
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 3320 13787 3378 13793
rect 3320 13753 3332 13787
rect 3366 13784 3378 13787
rect 4062 13784 4068 13796
rect 3366 13756 4068 13784
rect 3366 13753 3378 13756
rect 3320 13747 3378 13753
rect 4062 13744 4068 13756
rect 4120 13744 4126 13796
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 6270 13784 6276 13796
rect 5592 13756 6276 13784
rect 5592 13744 5598 13756
rect 6270 13744 6276 13756
rect 6328 13784 6334 13796
rect 7098 13793 7104 13796
rect 7092 13784 7104 13793
rect 6328 13756 7104 13784
rect 6328 13744 6334 13756
rect 7092 13747 7104 13756
rect 7098 13744 7104 13747
rect 7156 13744 7162 13796
rect 7742 13744 7748 13796
rect 7800 13784 7806 13796
rect 8570 13784 8576 13796
rect 7800 13756 8576 13784
rect 7800 13744 7806 13756
rect 8570 13744 8576 13756
rect 8628 13744 8634 13796
rect 8754 13744 8760 13796
rect 8812 13784 8818 13796
rect 8910 13787 8968 13793
rect 8910 13784 8922 13787
rect 8812 13756 8922 13784
rect 8812 13744 8818 13756
rect 8910 13753 8922 13756
rect 8956 13753 8968 13787
rect 8910 13747 8968 13753
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 10965 13787 11023 13793
rect 10965 13784 10977 13787
rect 9456 13756 10977 13784
rect 9456 13744 9462 13756
rect 10965 13753 10977 13756
rect 11011 13753 11023 13787
rect 11698 13784 11704 13796
rect 11659 13756 11704 13784
rect 10965 13747 11023 13753
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12897 13787 12955 13793
rect 12897 13784 12909 13787
rect 11808 13756 12909 13784
rect 2317 13719 2375 13725
rect 2317 13685 2329 13719
rect 2363 13716 2375 13719
rect 4338 13716 4344 13728
rect 2363 13688 4344 13716
rect 2363 13685 2375 13688
rect 2317 13679 2375 13685
rect 4338 13676 4344 13688
rect 4396 13676 4402 13728
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 9674 13716 9680 13728
rect 4856 13688 9680 13716
rect 4856 13676 4862 13688
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10560 13688 10885 13716
rect 10560 13676 10566 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 10873 13679 10931 13685
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 11808 13716 11836 13756
rect 12897 13753 12909 13756
rect 12943 13753 12955 13787
rect 13630 13784 13636 13796
rect 13591 13756 13636 13784
rect 12897 13747 12955 13753
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 11204 13688 11836 13716
rect 11204 13676 11210 13688
rect 12342 13676 12348 13728
rect 12400 13716 12406 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 12400 13688 12817 13716
rect 12400 13676 12406 13688
rect 12805 13685 12817 13688
rect 12851 13685 12863 13719
rect 12805 13679 12863 13685
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 2038 13512 2044 13524
rect 1999 13484 2044 13512
rect 2038 13472 2044 13484
rect 2096 13472 2102 13524
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 3050 13512 3056 13524
rect 2823 13484 3056 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3145 13515 3203 13521
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 7374 13512 7380 13524
rect 3191 13484 7380 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 7926 13512 7932 13524
rect 7668 13484 7932 13512
rect 4798 13444 4804 13456
rect 4759 13416 4804 13444
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 7668 13444 7696 13484
rect 7926 13472 7932 13484
rect 7984 13512 7990 13524
rect 8754 13512 8760 13524
rect 7984 13484 8760 13512
rect 7984 13472 7990 13484
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13512 9367 13515
rect 9490 13512 9496 13524
rect 9355 13484 9496 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 10008 13484 10057 13512
rect 10008 13472 10014 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13481 10931 13515
rect 10873 13475 10931 13481
rect 7300 13416 7696 13444
rect 7736 13447 7794 13453
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 4706 13376 4712 13388
rect 1995 13348 4712 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 5902 13385 5908 13388
rect 5896 13376 5908 13385
rect 5863 13348 5908 13376
rect 5896 13339 5908 13348
rect 5960 13376 5966 13388
rect 7300 13376 7328 13416
rect 7736 13413 7748 13447
rect 7782 13444 7794 13447
rect 7834 13444 7840 13456
rect 7782 13416 7840 13444
rect 7782 13413 7794 13416
rect 7736 13407 7794 13413
rect 7834 13404 7840 13416
rect 7892 13404 7898 13456
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 10888 13444 10916 13475
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11204 13484 12081 13512
rect 11204 13472 11210 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 12250 13472 12256 13524
rect 12308 13472 12314 13524
rect 13262 13512 13268 13524
rect 13223 13484 13268 13512
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 13722 13512 13728 13524
rect 13683 13484 13728 13512
rect 13722 13472 13728 13484
rect 13780 13512 13786 13524
rect 14458 13512 14464 13524
rect 13780 13484 14320 13512
rect 14419 13484 14464 13512
rect 13780 13472 13786 13484
rect 8260 13416 10916 13444
rect 11333 13447 11391 13453
rect 8260 13404 8266 13416
rect 11333 13413 11345 13447
rect 11379 13444 11391 13447
rect 11422 13444 11428 13456
rect 11379 13416 11428 13444
rect 11379 13413 11391 13416
rect 11333 13407 11391 13413
rect 11422 13404 11428 13416
rect 11480 13444 11486 13456
rect 12268 13444 12296 13472
rect 11480 13416 12296 13444
rect 11480 13404 11486 13416
rect 13078 13404 13084 13456
rect 13136 13444 13142 13456
rect 13633 13447 13691 13453
rect 13633 13444 13645 13447
rect 13136 13416 13645 13444
rect 13136 13404 13142 13416
rect 13633 13413 13645 13416
rect 13679 13444 13691 13447
rect 14292 13444 14320 13484
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 15286 13444 15292 13456
rect 13679 13416 13768 13444
rect 14292 13416 15292 13444
rect 13679 13413 13691 13416
rect 13633 13407 13691 13413
rect 13740 13388 13768 13416
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 7466 13376 7472 13388
rect 5960 13348 7328 13376
rect 7427 13348 7472 13376
rect 5902 13336 5908 13339
rect 5960 13336 5966 13348
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 7558 13336 7564 13388
rect 7616 13376 7622 13388
rect 8846 13376 8852 13388
rect 7616 13348 8852 13376
rect 7616 13336 7622 13348
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9493 13379 9551 13385
rect 9493 13376 9505 13379
rect 9456 13348 9505 13376
rect 9456 13336 9462 13348
rect 9493 13345 9505 13348
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13376 11299 13379
rect 11698 13376 11704 13388
rect 11287 13348 11704 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 12250 13336 12256 13388
rect 12308 13376 12314 13388
rect 12434 13376 12440 13388
rect 12308 13348 12440 13376
rect 12308 13336 12314 13348
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13722 13336 13728 13388
rect 13780 13336 13786 13388
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 2406 13308 2412 13320
rect 2271 13280 2412 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 2556 13280 3249 13308
rect 2556 13268 2562 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3344 13240 3372 13271
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4893 13311 4951 13317
rect 4396 13280 4660 13308
rect 4396 13268 4402 13280
rect 4632 13240 4660 13280
rect 4893 13277 4905 13311
rect 4939 13277 4951 13311
rect 5074 13308 5080 13320
rect 5035 13280 5080 13308
rect 4893 13271 4951 13277
rect 4908 13240 4936 13271
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 5629 13311 5687 13317
rect 5629 13308 5641 13311
rect 5500 13280 5641 13308
rect 5500 13268 5506 13280
rect 5629 13277 5641 13280
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 10100 13280 10149 13308
rect 10100 13268 10106 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 11146 13308 11152 13320
rect 10367 13280 11152 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13277 12587 13311
rect 12710 13308 12716 13320
rect 12671 13280 12716 13308
rect 12529 13271 12587 13277
rect 3344 13212 4568 13240
rect 4632 13212 4936 13240
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 4154 13172 4160 13184
rect 1627 13144 4160 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 4430 13172 4436 13184
rect 4391 13144 4436 13172
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 4540 13172 4568 13212
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 8849 13243 8907 13249
rect 8849 13240 8861 13243
rect 8628 13212 8861 13240
rect 8628 13200 8634 13212
rect 8849 13209 8861 13212
rect 8895 13209 8907 13243
rect 8849 13203 8907 13209
rect 9416 13212 10916 13240
rect 5166 13172 5172 13184
rect 4540 13144 5172 13172
rect 5166 13132 5172 13144
rect 5224 13172 5230 13184
rect 7009 13175 7067 13181
rect 7009 13172 7021 13175
rect 5224 13144 7021 13172
rect 5224 13132 5230 13144
rect 7009 13141 7021 13144
rect 7055 13141 7067 13175
rect 7009 13135 7067 13141
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 9416 13172 9444 13212
rect 7892 13144 9444 13172
rect 7892 13132 7898 13144
rect 9490 13132 9496 13184
rect 9548 13172 9554 13184
rect 9677 13175 9735 13181
rect 9677 13172 9689 13175
rect 9548 13144 9689 13172
rect 9548 13132 9554 13144
rect 9677 13141 9689 13144
rect 9723 13141 9735 13175
rect 9677 13135 9735 13141
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 10778 13172 10784 13184
rect 10008 13144 10784 13172
rect 10008 13132 10014 13144
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 10888 13172 10916 13212
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 11532 13240 11560 13271
rect 12434 13240 12440 13252
rect 11112 13212 12440 13240
rect 11112 13200 11118 13212
rect 12434 13200 12440 13212
rect 12492 13200 12498 13252
rect 12544 13240 12572 13271
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 13814 13308 13820 13320
rect 13775 13280 13820 13308
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 14366 13240 14372 13252
rect 12544 13212 14372 13240
rect 14366 13200 14372 13212
rect 14424 13240 14430 13252
rect 14642 13240 14648 13252
rect 14424 13212 14648 13240
rect 14424 13200 14430 13212
rect 14642 13200 14648 13212
rect 14700 13200 14706 13252
rect 11974 13172 11980 13184
rect 10888 13144 11980 13172
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 2498 12968 2504 12980
rect 2459 12940 2504 12968
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 4246 12968 4252 12980
rect 3160 12940 4252 12968
rect 3160 12841 3188 12940
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 10410 12968 10416 12980
rect 4764 12940 10416 12968
rect 4764 12928 4770 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 12437 12971 12495 12977
rect 12437 12968 12449 12971
rect 11020 12940 12449 12968
rect 11020 12928 11026 12940
rect 12437 12937 12449 12940
rect 12483 12937 12495 12971
rect 12437 12931 12495 12937
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13906 12968 13912 12980
rect 13044 12940 13912 12968
rect 13044 12928 13050 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 3697 12903 3755 12909
rect 3697 12869 3709 12903
rect 3743 12900 3755 12903
rect 4062 12900 4068 12912
rect 3743 12872 4068 12900
rect 3743 12869 3755 12872
rect 3697 12863 3755 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 4798 12900 4804 12912
rect 4356 12872 4804 12900
rect 4356 12841 4384 12872
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 4890 12860 4896 12912
rect 4948 12860 4954 12912
rect 6270 12900 6276 12912
rect 6231 12872 6276 12900
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 8018 12860 8024 12912
rect 8076 12900 8082 12912
rect 8205 12903 8263 12909
rect 8205 12900 8217 12903
rect 8076 12872 8217 12900
rect 8076 12860 8082 12872
rect 8205 12869 8217 12872
rect 8251 12869 8263 12903
rect 8205 12863 8263 12869
rect 10045 12903 10103 12909
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 10226 12900 10232 12912
rect 10091 12872 10232 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10505 12903 10563 12909
rect 10505 12869 10517 12903
rect 10551 12900 10563 12903
rect 12342 12900 12348 12912
rect 10551 12872 12348 12900
rect 10551 12869 10563 12872
rect 10505 12863 10563 12869
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12764 1639 12767
rect 2590 12764 2596 12776
rect 1627 12736 2596 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 4908 12773 4936 12860
rect 8110 12792 8116 12844
rect 8168 12832 8174 12844
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8168 12804 8677 12832
rect 8168 12792 8174 12804
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 10870 12832 10876 12844
rect 10468 12804 10876 12832
rect 10468 12792 10474 12804
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12801 11115 12835
rect 11698 12832 11704 12844
rect 11659 12804 11704 12832
rect 11057 12795 11115 12801
rect 5166 12773 5172 12776
rect 4065 12767 4123 12773
rect 4065 12733 4077 12767
rect 4111 12764 4123 12767
rect 4893 12767 4951 12773
rect 4111 12736 4844 12764
rect 4111 12733 4123 12736
rect 4065 12727 4123 12733
rect 1394 12656 1400 12708
rect 1452 12696 1458 12708
rect 1857 12699 1915 12705
rect 1857 12696 1869 12699
rect 1452 12668 1869 12696
rect 1452 12656 1458 12668
rect 1857 12665 1869 12668
rect 1903 12665 1915 12699
rect 1857 12659 1915 12665
rect 2869 12699 2927 12705
rect 2869 12665 2881 12699
rect 2915 12696 2927 12699
rect 4157 12699 4215 12705
rect 2915 12668 4108 12696
rect 2915 12665 2927 12668
rect 2869 12659 2927 12665
rect 2958 12628 2964 12640
rect 2919 12600 2964 12628
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 4080 12628 4108 12668
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 4706 12696 4712 12708
rect 4203 12668 4712 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 4706 12656 4712 12668
rect 4764 12656 4770 12708
rect 4816 12696 4844 12736
rect 4893 12733 4905 12767
rect 4939 12733 4951 12767
rect 5160 12764 5172 12773
rect 5127 12736 5172 12764
rect 4893 12727 4951 12733
rect 5160 12727 5172 12736
rect 5166 12724 5172 12727
rect 5224 12724 5230 12776
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 6730 12764 6736 12776
rect 5500 12736 6736 12764
rect 5500 12724 5506 12736
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 6914 12764 6920 12776
rect 6871 12736 6920 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 7024 12736 7963 12764
rect 7024 12696 7052 12736
rect 7098 12705 7104 12708
rect 4816 12668 7052 12696
rect 7092 12659 7104 12705
rect 7156 12696 7162 12708
rect 7156 12668 7192 12696
rect 7098 12656 7104 12659
rect 7156 12656 7162 12668
rect 7834 12628 7840 12640
rect 4080 12600 7840 12628
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 7935 12628 7963 12736
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 11072 12764 11100 12795
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12066 12792 12072 12844
rect 12124 12792 12130 12844
rect 12158 12792 12164 12844
rect 12216 12792 12222 12844
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12768 12804 13001 12832
rect 12768 12792 12774 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 12989 12795 13047 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 11146 12764 11152 12776
rect 8352 12736 11152 12764
rect 8352 12724 8358 12736
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 8932 12699 8990 12705
rect 8932 12665 8944 12699
rect 8978 12696 8990 12699
rect 9306 12696 9312 12708
rect 8978 12668 9312 12696
rect 8978 12665 8990 12668
rect 8932 12659 8990 12665
rect 9306 12656 9312 12668
rect 9364 12656 9370 12708
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 9640 12668 10977 12696
rect 9640 12656 9646 12668
rect 10965 12665 10977 12668
rect 11011 12696 11023 12699
rect 11238 12696 11244 12708
rect 11011 12668 11244 12696
rect 11011 12665 11023 12668
rect 10965 12659 11023 12665
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 12084 12696 12112 12792
rect 12176 12764 12204 12792
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12176 12736 12817 12764
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12764 12955 12767
rect 13170 12764 13176 12776
rect 12943 12736 13176 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 13906 12764 13912 12776
rect 13679 12736 13912 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 13906 12724 13912 12736
rect 13964 12764 13970 12776
rect 14182 12764 14188 12776
rect 13964 12736 14188 12764
rect 13964 12724 13970 12736
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14550 12764 14556 12776
rect 14511 12736 14556 12764
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 12158 12696 12164 12708
rect 12084 12668 12164 12696
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 14826 12696 14832 12708
rect 14787 12668 14832 12696
rect 14826 12656 14832 12668
rect 14884 12656 14890 12708
rect 10226 12628 10232 12640
rect 7935 12600 10232 12628
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 10873 12631 10931 12637
rect 10873 12597 10885 12631
rect 10919 12628 10931 12631
rect 11514 12628 11520 12640
rect 10919 12600 11520 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 1596 12356 1624 12387
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 1949 12427 2007 12433
rect 1949 12424 1961 12427
rect 1912 12396 1961 12424
rect 1912 12384 1918 12396
rect 1949 12393 1961 12396
rect 1995 12393 2007 12427
rect 1949 12387 2007 12393
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 2958 12424 2964 12436
rect 2823 12396 2964 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 4154 12424 4160 12436
rect 3191 12396 4160 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 4982 12424 4988 12436
rect 4724 12396 4988 12424
rect 3878 12356 3884 12368
rect 1596 12328 3884 12356
rect 3878 12316 3884 12328
rect 3936 12316 3942 12368
rect 4522 12316 4528 12368
rect 4580 12356 4586 12368
rect 4724 12365 4752 12396
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 6270 12424 6276 12436
rect 5132 12396 6276 12424
rect 5132 12384 5138 12396
rect 6270 12384 6276 12396
rect 6328 12424 6334 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6328 12396 6929 12424
rect 6328 12384 6334 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 8202 12424 8208 12436
rect 7156 12396 8208 12424
rect 7156 12384 7162 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8754 12424 8760 12436
rect 8715 12396 8760 12424
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 8904 12396 9229 12424
rect 8904 12384 8910 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9217 12387 9275 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 12066 12424 12072 12436
rect 10008 12396 11560 12424
rect 12027 12396 12072 12424
rect 10008 12384 10014 12396
rect 4709 12359 4767 12365
rect 4709 12356 4721 12359
rect 4580 12328 4721 12356
rect 4580 12316 4586 12328
rect 4709 12325 4721 12328
rect 4755 12325 4767 12359
rect 7622 12359 7680 12365
rect 7622 12356 7634 12359
rect 4709 12319 4767 12325
rect 5276 12328 7634 12356
rect 2038 12288 2044 12300
rect 1999 12260 2044 12288
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 5276 12288 5304 12328
rect 7622 12325 7634 12328
rect 7668 12356 7680 12359
rect 8018 12356 8024 12368
rect 7668 12328 8024 12356
rect 7668 12325 7680 12328
rect 7622 12319 7680 12325
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 8128 12328 11008 12356
rect 5804 12291 5862 12297
rect 5804 12288 5816 12291
rect 3436 12260 5304 12288
rect 5368 12260 5816 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2314 12220 2320 12232
rect 2271 12192 2320 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 3436 12229 3464 12260
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3252 12084 3280 12183
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4120 12192 4813 12220
rect 4120 12180 4126 12192
rect 4801 12189 4813 12192
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5368 12220 5396 12260
rect 5804 12257 5816 12260
rect 5850 12288 5862 12291
rect 6730 12288 6736 12300
rect 5850 12260 6736 12288
rect 5850 12257 5862 12260
rect 5804 12251 5862 12257
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7064 12260 7389 12288
rect 7064 12248 7070 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 8128 12288 8156 12328
rect 9398 12288 9404 12300
rect 7377 12251 7435 12257
rect 7484 12260 8156 12288
rect 9359 12260 9404 12288
rect 5534 12220 5540 12232
rect 5031 12192 5396 12220
rect 5495 12192 5540 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 7484 12220 7512 12260
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10042 12288 10048 12300
rect 9732 12260 10048 12288
rect 9732 12248 9738 12260
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 6696 12192 7512 12220
rect 6696 12180 6702 12192
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9364 12192 10149 12220
rect 9364 12180 9370 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10042 12112 10048 12164
rect 10100 12152 10106 12164
rect 10244 12152 10272 12183
rect 10100 12124 10272 12152
rect 10100 12112 10106 12124
rect 10873 12087 10931 12093
rect 10873 12084 10885 12087
rect 3252 12056 10885 12084
rect 10873 12053 10885 12056
rect 10919 12053 10931 12087
rect 10980 12084 11008 12328
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 11532 12356 11560 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12400 12396 12541 12424
rect 12400 12384 12406 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 13262 12424 13268 12436
rect 13223 12396 13268 12424
rect 12529 12387 12587 12393
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12393 14703 12427
rect 14645 12387 14703 12393
rect 14660 12356 14688 12387
rect 11204 12328 11468 12356
rect 11532 12328 14688 12356
rect 11204 12316 11210 12328
rect 11238 12288 11244 12300
rect 11199 12260 11244 12288
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11330 12220 11336 12232
rect 11291 12192 11336 12220
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11440 12229 11468 12328
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 12032 12260 12449 12288
rect 12032 12248 12038 12260
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 13630 12288 13636 12300
rect 13591 12260 13636 12288
rect 12437 12251 12495 12257
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 14182 12248 14188 12300
rect 14240 12288 14246 12300
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 14240 12260 14473 12288
rect 14240 12248 14246 12260
rect 14461 12257 14473 12260
rect 14507 12288 14519 12291
rect 15010 12288 15016 12300
rect 14507 12260 15016 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 12584 12192 12633 12220
rect 12584 12180 12590 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 13722 12220 13728 12232
rect 13683 12192 13728 12220
rect 12621 12183 12679 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 13817 12223 13875 12229
rect 13817 12189 13829 12223
rect 13863 12189 13875 12223
rect 13817 12183 13875 12189
rect 13832 12152 13860 12183
rect 11624 12124 13860 12152
rect 11624 12084 11652 12124
rect 10980 12056 11652 12084
rect 10873 12047 10931 12053
rect 12342 12044 12348 12096
rect 12400 12084 12406 12096
rect 13078 12084 13084 12096
rect 12400 12056 13084 12084
rect 12400 12044 12406 12056
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 1854 11880 1860 11892
rect 1815 11852 1860 11880
rect 1854 11840 1860 11852
rect 1912 11840 1918 11892
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 6362 11880 6368 11892
rect 5592 11852 6368 11880
rect 5592 11840 5598 11852
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 8202 11880 8208 11892
rect 8163 11852 8208 11880
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 9950 11880 9956 11892
rect 8312 11852 9956 11880
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 2958 11744 2964 11756
rect 2547 11716 2964 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 6380 11744 6408 11840
rect 8018 11772 8024 11824
rect 8076 11812 8082 11824
rect 8312 11812 8340 11852
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10502 11880 10508 11892
rect 10463 11852 10508 11880
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 11572 11852 15025 11880
rect 11572 11840 11578 11852
rect 15013 11849 15025 11852
rect 15059 11849 15071 11883
rect 15013 11843 15071 11849
rect 8076 11784 8340 11812
rect 9692 11784 9996 11812
rect 8076 11772 8082 11784
rect 6822 11744 6828 11756
rect 4212 11716 5028 11744
rect 6380 11716 6828 11744
rect 4212 11704 4218 11716
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 2682 11676 2688 11688
rect 2363 11648 2688 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3053 11679 3111 11685
rect 3053 11676 3065 11679
rect 2832 11648 3065 11676
rect 2832 11636 2838 11648
rect 3053 11645 3065 11648
rect 3099 11676 3111 11679
rect 4798 11676 4804 11688
rect 3099 11648 4804 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 4798 11636 4804 11648
rect 4856 11676 4862 11688
rect 4893 11679 4951 11685
rect 4893 11676 4905 11679
rect 4856 11648 4905 11676
rect 4856 11636 4862 11648
rect 4893 11645 4905 11648
rect 4939 11645 4951 11679
rect 5000 11676 5028 11716
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 6638 11676 6644 11688
rect 5000 11648 6644 11676
rect 4893 11639 4951 11645
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 6840 11676 6868 11704
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 6840 11648 8677 11676
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 9692 11676 9720 11784
rect 9968 11756 9996 11784
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 11664 11784 11744 11812
rect 11664 11772 11670 11784
rect 9858 11704 9864 11756
rect 9916 11704 9922 11756
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 11716 11753 11744 11784
rect 12066 11772 12072 11824
rect 12124 11812 12130 11824
rect 12437 11815 12495 11821
rect 12437 11812 12449 11815
rect 12124 11784 12449 11812
rect 12124 11772 12130 11784
rect 12437 11781 12449 11784
rect 12483 11781 12495 11815
rect 12437 11775 12495 11781
rect 13078 11772 13084 11824
rect 13136 11812 13142 11824
rect 13633 11815 13691 11821
rect 13633 11812 13645 11815
rect 13136 11784 13645 11812
rect 13136 11772 13142 11784
rect 13633 11781 13645 11784
rect 13679 11781 13691 11815
rect 13633 11775 13691 11781
rect 13998 11772 14004 11824
rect 14056 11812 14062 11824
rect 14458 11812 14464 11824
rect 14056 11784 14464 11812
rect 14056 11772 14062 11784
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 10100 11716 11069 11744
rect 10100 11704 10106 11716
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12676 11716 13001 11744
rect 12676 11704 12682 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13262 11704 13268 11756
rect 13320 11744 13326 11756
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13320 11716 14197 11744
rect 13320 11704 13326 11716
rect 14185 11713 14197 11716
rect 14231 11744 14243 11747
rect 15102 11744 15108 11756
rect 14231 11716 15108 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 9876 11676 9904 11704
rect 8665 11639 8723 11645
rect 8772 11648 9720 11676
rect 9784 11648 9904 11676
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 3142 11608 3148 11620
rect 2271 11580 3148 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 3320 11611 3378 11617
rect 3320 11608 3332 11611
rect 3252 11580 3332 11608
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 3252 11540 3280 11580
rect 3320 11577 3332 11580
rect 3366 11608 3378 11611
rect 3366 11580 3832 11608
rect 3366 11577 3378 11580
rect 3320 11571 3378 11577
rect 2372 11512 3280 11540
rect 3804 11540 3832 11580
rect 3878 11568 3884 11620
rect 3936 11608 3942 11620
rect 5160 11611 5218 11617
rect 3936 11580 5028 11608
rect 3936 11568 3942 11580
rect 4154 11540 4160 11552
rect 3804 11512 4160 11540
rect 2372 11500 2378 11512
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4433 11543 4491 11549
rect 4433 11509 4445 11543
rect 4479 11540 4491 11543
rect 4614 11540 4620 11552
rect 4479 11512 4620 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 4614 11500 4620 11512
rect 4672 11540 4678 11552
rect 4890 11540 4896 11552
rect 4672 11512 4896 11540
rect 4672 11500 4678 11512
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5000 11540 5028 11580
rect 5160 11577 5172 11611
rect 5206 11608 5218 11611
rect 6178 11608 6184 11620
rect 5206 11580 6184 11608
rect 5206 11577 5218 11580
rect 5160 11571 5218 11577
rect 6178 11568 6184 11580
rect 6236 11568 6242 11620
rect 7070 11611 7128 11617
rect 7070 11608 7082 11611
rect 6288 11580 7082 11608
rect 6288 11552 6316 11580
rect 7070 11577 7082 11580
rect 7116 11577 7128 11611
rect 7070 11571 7128 11577
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 8772 11608 8800 11648
rect 7248 11580 8800 11608
rect 8932 11611 8990 11617
rect 7248 11568 7254 11580
rect 8932 11577 8944 11611
rect 8978 11608 8990 11611
rect 9306 11608 9312 11620
rect 8978 11580 9312 11608
rect 8978 11577 8990 11580
rect 8932 11571 8990 11577
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 9784 11608 9812 11648
rect 10134 11636 10140 11688
rect 10192 11676 10198 11688
rect 10192 11648 11652 11676
rect 10192 11636 10198 11648
rect 9640 11580 9812 11608
rect 9640 11568 9646 11580
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 11514 11608 11520 11620
rect 9916 11580 11520 11608
rect 9916 11568 9922 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 5718 11540 5724 11552
rect 5000 11512 5724 11540
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 6270 11540 6276 11552
rect 6231 11512 6276 11540
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 9490 11540 9496 11552
rect 6696 11512 9496 11540
rect 6696 11500 6702 11512
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 10045 11543 10103 11549
rect 10045 11540 10057 11543
rect 9824 11512 10057 11540
rect 9824 11500 9830 11512
rect 10045 11509 10057 11512
rect 10091 11509 10103 11543
rect 10045 11503 10103 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10376 11512 10885 11540
rect 10376 11500 10382 11512
rect 10873 11509 10885 11512
rect 10919 11509 10931 11543
rect 10873 11503 10931 11509
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 11624 11540 11652 11648
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12492 11648 12817 11676
rect 12492 11636 12498 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 14734 11676 14740 11688
rect 13504 11648 14740 11676
rect 13504 11636 13510 11648
rect 14734 11636 14740 11648
rect 14792 11676 14798 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 14792 11648 14841 11676
rect 14792 11636 14798 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 11698 11568 11704 11620
rect 11756 11608 11762 11620
rect 11882 11608 11888 11620
rect 11756 11580 11888 11608
rect 11756 11568 11762 11580
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12986 11608 12992 11620
rect 12216 11580 12992 11608
rect 12216 11568 12222 11580
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 13078 11568 13084 11620
rect 13136 11608 13142 11620
rect 14001 11611 14059 11617
rect 14001 11608 14013 11611
rect 13136 11580 14013 11608
rect 13136 11568 13142 11580
rect 14001 11577 14013 11580
rect 14047 11577 14059 11611
rect 14001 11571 14059 11577
rect 12710 11540 12716 11552
rect 11011 11512 12716 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13538 11540 13544 11552
rect 12943 11512 13544 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 14093 11543 14151 11549
rect 14093 11540 14105 11543
rect 13964 11512 14105 11540
rect 13964 11500 13970 11512
rect 14093 11509 14105 11512
rect 14139 11509 14151 11543
rect 14093 11503 14151 11509
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1762 11336 1768 11348
rect 1627 11308 1768 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 2041 11339 2099 11345
rect 2041 11305 2053 11339
rect 2087 11336 2099 11339
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2087 11308 2789 11336
rect 2087 11305 2099 11308
rect 2041 11299 2099 11305
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 2777 11299 2835 11305
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3878 11336 3884 11348
rect 3191 11308 3884 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4396 11308 4537 11336
rect 4396 11296 4402 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 6641 11339 6699 11345
rect 6641 11336 6653 11339
rect 4525 11299 4583 11305
rect 4724 11308 6653 11336
rect 2685 11271 2743 11277
rect 2685 11237 2697 11271
rect 2731 11268 2743 11271
rect 3237 11271 3295 11277
rect 3237 11268 3249 11271
rect 2731 11240 3249 11268
rect 2731 11237 2743 11240
rect 2685 11231 2743 11237
rect 3237 11237 3249 11240
rect 3283 11268 3295 11271
rect 4614 11268 4620 11280
rect 3283 11240 4620 11268
rect 3283 11237 3295 11240
rect 3237 11231 3295 11237
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 1946 11200 1952 11212
rect 1907 11172 1952 11200
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4028 11172 4445 11200
rect 4028 11160 4034 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 3142 11132 3148 11144
rect 2271 11104 3148 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 4338 11132 4344 11144
rect 3467 11104 4344 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4724 11141 4752 11308
rect 6641 11305 6653 11308
rect 6687 11305 6699 11339
rect 6641 11299 6699 11305
rect 4890 11228 4896 11280
rect 4948 11268 4954 11280
rect 5506 11271 5564 11277
rect 5506 11268 5518 11271
rect 4948 11240 5518 11268
rect 4948 11228 4954 11240
rect 5506 11237 5518 11240
rect 5552 11237 5564 11271
rect 5506 11231 5564 11237
rect 5718 11228 5724 11280
rect 5776 11228 5782 11280
rect 6656 11268 6684 11299
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 8481 11339 8539 11345
rect 8481 11336 8493 11339
rect 6788 11308 8493 11336
rect 6788 11296 6794 11308
rect 8481 11305 8493 11308
rect 8527 11305 8539 11339
rect 8481 11299 8539 11305
rect 10045 11339 10103 11345
rect 10045 11305 10057 11339
rect 10091 11336 10103 11339
rect 11606 11336 11612 11348
rect 10091 11308 11612 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 7346 11271 7404 11277
rect 7346 11268 7358 11271
rect 6656 11240 7358 11268
rect 7346 11237 7358 11240
rect 7392 11237 7404 11271
rect 7346 11231 7404 11237
rect 5736 11200 5764 11228
rect 5736 11172 6776 11200
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 6748 11132 6776 11172
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6880 11172 7113 11200
rect 6880 11160 6886 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 8496 11200 8524 11299
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 12342 11336 12348 11348
rect 11940 11308 12348 11336
rect 11940 11296 11946 11308
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 12526 11336 12532 11348
rect 12483 11308 12532 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 12710 11296 12716 11348
rect 12768 11296 12774 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13630 11336 13636 11348
rect 13311 11308 13636 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 8628 11240 8953 11268
rect 8628 11228 8634 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 8941 11231 8999 11237
rect 10137 11271 10195 11277
rect 10137 11237 10149 11271
rect 10183 11268 10195 11271
rect 12158 11268 12164 11280
rect 10183 11240 12164 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 12728 11268 12756 11296
rect 14550 11268 14556 11280
rect 12728 11240 14556 11268
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 10042 11200 10048 11212
rect 7101 11163 7159 11169
rect 7208 11172 8432 11200
rect 8496 11172 10048 11200
rect 7208 11132 7236 11172
rect 5316 11104 5361 11132
rect 6748 11104 7236 11132
rect 8404 11132 8432 11172
rect 10042 11160 10048 11172
rect 10100 11200 10106 11212
rect 10100 11172 10272 11200
rect 10100 11160 10106 11172
rect 10244 11141 10272 11172
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11204 11172 11253 11200
rect 11204 11160 11210 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11388 11172 12296 11200
rect 11388 11160 11394 11172
rect 10229 11135 10287 11141
rect 8404 11104 10180 11132
rect 5316 11092 5322 11104
rect 8570 11024 8576 11076
rect 8628 11024 8634 11076
rect 9677 11067 9735 11073
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 10152 11064 10180 11104
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 10376 11104 11437 11132
rect 10376 11092 10382 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 12268 11132 12296 11172
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 12529 11203 12587 11209
rect 12529 11200 12541 11203
rect 12400 11172 12541 11200
rect 12400 11160 12406 11172
rect 12529 11169 12541 11172
rect 12575 11169 12587 11203
rect 12529 11163 12587 11169
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 12768 11172 13645 11200
rect 12768 11160 12774 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 14458 11200 14464 11212
rect 14419 11172 14464 11200
rect 13633 11163 13691 11169
rect 14458 11160 14464 11172
rect 14516 11160 14522 11212
rect 12434 11132 12440 11144
rect 12268 11104 12440 11132
rect 11425 11095 11483 11101
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 12618 11132 12624 11144
rect 12579 11104 12624 11132
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 13725 11135 13783 11141
rect 13725 11132 13737 11135
rect 13596 11104 13737 11132
rect 13596 11092 13602 11104
rect 13725 11101 13737 11104
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11132 13967 11135
rect 14182 11132 14188 11144
rect 13955 11104 14188 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 11974 11064 11980 11076
rect 9723 11036 10088 11064
rect 10152 11036 11980 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 2130 10956 2136 11008
rect 2188 10996 2194 11008
rect 8588 10996 8616 11024
rect 2188 10968 8616 10996
rect 10060 10996 10088 11036
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 12342 11024 12348 11076
rect 12400 11064 12406 11076
rect 14645 11067 14703 11073
rect 14645 11064 14657 11067
rect 12400 11036 14657 11064
rect 12400 11024 12406 11036
rect 14645 11033 14657 11036
rect 14691 11033 14703 11067
rect 14645 11027 14703 11033
rect 10226 10996 10232 11008
rect 10060 10968 10232 10996
rect 2188 10956 2194 10968
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10870 10996 10876 11008
rect 10831 10968 10876 10996
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 12066 10996 12072 11008
rect 12027 10968 12072 10996
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 1857 10795 1915 10801
rect 1857 10761 1869 10795
rect 1903 10792 1915 10795
rect 1946 10792 1952 10804
rect 1903 10764 1952 10792
rect 1903 10761 1915 10764
rect 1857 10755 1915 10761
rect 1946 10752 1952 10764
rect 2004 10752 2010 10804
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 9398 10792 9404 10804
rect 5031 10764 9404 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10502 10792 10508 10804
rect 10091 10764 10508 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11204 10764 12388 10792
rect 11204 10752 11210 10764
rect 4154 10684 4160 10736
rect 4212 10724 4218 10736
rect 4433 10727 4491 10733
rect 4433 10724 4445 10727
rect 4212 10696 4445 10724
rect 4212 10684 4218 10696
rect 4433 10693 4445 10696
rect 4479 10724 4491 10727
rect 5166 10724 5172 10736
rect 4479 10696 5172 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 8662 10724 8668 10736
rect 7892 10696 8668 10724
rect 7892 10684 7898 10696
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 12360 10724 12388 10764
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12492 10764 12940 10792
rect 12492 10752 12498 10764
rect 9692 10696 11652 10724
rect 12360 10696 12848 10724
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 2547 10628 3188 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 2832 10560 3065 10588
rect 2832 10548 2838 10560
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3160 10588 3188 10628
rect 4798 10616 4804 10668
rect 4856 10656 4862 10668
rect 5258 10656 5264 10668
rect 4856 10628 5264 10656
rect 4856 10616 4862 10628
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 4338 10588 4344 10600
rect 3160 10560 4344 10588
rect 3053 10551 3111 10557
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 5169 10591 5227 10597
rect 5169 10557 5181 10591
rect 5215 10557 5227 10591
rect 6840 10588 6868 10616
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 5169 10551 5227 10557
rect 5276 10560 6776 10588
rect 6840 10560 8677 10588
rect 2314 10520 2320 10532
rect 2275 10492 2320 10520
rect 2314 10480 2320 10492
rect 2372 10480 2378 10532
rect 2958 10480 2964 10532
rect 3016 10520 3022 10532
rect 3320 10523 3378 10529
rect 3320 10520 3332 10523
rect 3016 10492 3332 10520
rect 3016 10480 3022 10492
rect 3320 10489 3332 10492
rect 3366 10520 3378 10523
rect 3418 10520 3424 10532
rect 3366 10492 3424 10520
rect 3366 10489 3378 10492
rect 3320 10483 3378 10489
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 2225 10455 2283 10461
rect 2225 10452 2237 10455
rect 1636 10424 2237 10452
rect 1636 10412 1642 10424
rect 2225 10421 2237 10424
rect 2271 10421 2283 10455
rect 5184 10452 5212 10551
rect 5276 10532 5304 10560
rect 5258 10480 5264 10532
rect 5316 10480 5322 10532
rect 5442 10480 5448 10532
rect 5500 10529 5506 10532
rect 5500 10523 5564 10529
rect 5500 10489 5518 10523
rect 5552 10520 5564 10523
rect 5626 10520 5632 10532
rect 5552 10492 5632 10520
rect 5552 10489 5564 10492
rect 5500 10483 5564 10489
rect 5500 10480 5506 10483
rect 5626 10480 5632 10492
rect 5684 10480 5690 10532
rect 6454 10452 6460 10464
rect 5184 10424 6460 10452
rect 2225 10415 2283 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6638 10452 6644 10464
rect 6599 10424 6644 10452
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 6748 10452 6776 10560
rect 8665 10557 8677 10560
rect 8711 10557 8723 10591
rect 9692 10588 9720 10696
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10594 10656 10600 10668
rect 10192 10628 10600 10656
rect 10192 10616 10198 10628
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10928 10628 10977 10656
rect 10928 10616 10934 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 8665 10551 8723 10557
rect 8772 10560 9720 10588
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7070 10523 7128 10529
rect 7070 10520 7082 10523
rect 6972 10492 7082 10520
rect 6972 10480 6978 10492
rect 7070 10489 7082 10492
rect 7116 10489 7128 10523
rect 7070 10483 7128 10489
rect 7190 10480 7196 10532
rect 7248 10520 7254 10532
rect 8772 10520 8800 10560
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 11164 10588 11192 10619
rect 9824 10560 11192 10588
rect 11624 10588 11652 10696
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 12710 10656 12716 10668
rect 11747 10628 12716 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 12820 10597 12848 10696
rect 12912 10665 12940 10764
rect 12986 10752 12992 10804
rect 13044 10792 13050 10804
rect 13633 10795 13691 10801
rect 13044 10764 13584 10792
rect 13044 10752 13050 10764
rect 13556 10736 13584 10764
rect 13633 10761 13645 10795
rect 13679 10792 13691 10795
rect 13722 10792 13728 10804
rect 13679 10764 13728 10792
rect 13679 10761 13691 10764
rect 13633 10755 13691 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 13538 10684 13544 10736
rect 13596 10684 13602 10736
rect 14734 10724 14740 10736
rect 14108 10696 14740 10724
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13262 10656 13268 10668
rect 13127 10628 13268 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 13446 10616 13452 10668
rect 13504 10656 13510 10668
rect 14108 10665 14136 10696
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 14093 10659 14151 10665
rect 14093 10656 14105 10659
rect 13504 10628 14105 10656
rect 13504 10616 13510 10628
rect 14093 10625 14105 10628
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14182 10616 14188 10668
rect 14240 10656 14246 10668
rect 14240 10628 14333 10656
rect 14240 10616 14246 10628
rect 12805 10591 12863 10597
rect 11624 10560 12756 10588
rect 9824 10548 9830 10560
rect 7248 10492 8800 10520
rect 8932 10523 8990 10529
rect 7248 10480 7254 10492
rect 8932 10489 8944 10523
rect 8978 10520 8990 10523
rect 9030 10520 9036 10532
rect 8978 10492 9036 10520
rect 8978 10489 8990 10492
rect 8932 10483 8990 10489
rect 9030 10480 9036 10492
rect 9088 10520 9094 10532
rect 9398 10520 9404 10532
rect 9088 10492 9404 10520
rect 9088 10480 9094 10492
rect 9398 10480 9404 10492
rect 9456 10480 9462 10532
rect 10226 10480 10232 10532
rect 10284 10520 10290 10532
rect 11164 10520 11192 10560
rect 12618 10520 12624 10532
rect 10284 10492 11008 10520
rect 11164 10492 12624 10520
rect 10284 10480 10290 10492
rect 8110 10452 8116 10464
rect 6748 10424 8116 10452
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8205 10455 8263 10461
rect 8205 10421 8217 10455
rect 8251 10452 8263 10455
rect 9306 10452 9312 10464
rect 8251 10424 9312 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 10502 10452 10508 10464
rect 10463 10424 10508 10452
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 10594 10412 10600 10464
rect 10652 10452 10658 10464
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 10652 10424 10885 10452
rect 10652 10412 10658 10424
rect 10873 10421 10885 10424
rect 10919 10421 10931 10455
rect 10980 10452 11008 10492
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 12728 10520 12756 10560
rect 12805 10557 12817 10591
rect 12851 10557 12863 10591
rect 13722 10588 13728 10600
rect 12805 10551 12863 10557
rect 13556 10560 13728 10588
rect 13556 10520 13584 10560
rect 13722 10548 13728 10560
rect 13780 10588 13786 10600
rect 14200 10588 14228 10616
rect 13780 10560 14228 10588
rect 14829 10591 14887 10597
rect 13780 10548 13786 10560
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15286 10588 15292 10600
rect 14875 10560 15292 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 12728 10492 13584 10520
rect 11330 10452 11336 10464
rect 10980 10424 11336 10452
rect 10873 10415 10931 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 13446 10452 13452 10464
rect 12483 10424 13452 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13596 10424 14013 10452
rect 13596 10412 13602 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14001 10415 14059 10421
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14240 10424 15025 10452
rect 14240 10412 14246 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2087 10220 3372 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 1949 10183 2007 10189
rect 1949 10149 1961 10183
rect 1995 10180 2007 10183
rect 2130 10180 2136 10192
rect 1995 10152 2136 10180
rect 1995 10149 2007 10152
rect 1949 10143 2007 10149
rect 2130 10140 2136 10152
rect 2188 10140 2194 10192
rect 3344 10180 3372 10220
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 3476 10220 5825 10248
rect 3476 10208 3482 10220
rect 5813 10217 5825 10220
rect 5859 10248 5871 10251
rect 7190 10248 7196 10260
rect 5859 10220 7196 10248
rect 5859 10217 5871 10220
rect 5813 10211 5871 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 8754 10248 8760 10260
rect 7331 10220 8760 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9398 10248 9404 10260
rect 9079 10220 9404 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9398 10208 9404 10220
rect 9456 10248 9462 10260
rect 10134 10248 10140 10260
rect 9456 10220 9720 10248
rect 10095 10220 10140 10248
rect 9456 10208 9462 10220
rect 4522 10180 4528 10192
rect 3344 10152 4528 10180
rect 4522 10140 4528 10152
rect 4580 10140 4586 10192
rect 4700 10183 4758 10189
rect 4700 10149 4712 10183
rect 4746 10180 4758 10183
rect 6638 10180 6644 10192
rect 4746 10152 6644 10180
rect 4746 10149 4758 10152
rect 4700 10143 4758 10149
rect 6638 10140 6644 10152
rect 6696 10180 6702 10192
rect 9490 10180 9496 10192
rect 6696 10152 9496 10180
rect 6696 10140 6702 10152
rect 9490 10140 9496 10152
rect 9548 10140 9554 10192
rect 9692 10180 9720 10220
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 10468 10220 10548 10248
rect 10468 10208 10474 10220
rect 10520 10180 10548 10220
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10744 10220 10885 10248
rect 10744 10208 10750 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 12066 10248 12072 10260
rect 11287 10220 12072 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12434 10248 12440 10260
rect 12395 10220 12440 10248
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 13504 10220 13737 10248
rect 13504 10208 13510 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 13725 10211 13783 10217
rect 13262 10180 13268 10192
rect 9692 10152 10456 10180
rect 10520 10152 13268 10180
rect 3142 10112 3148 10124
rect 3103 10084 3148 10112
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 6178 10121 6184 10124
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 6172 10112 6184 10121
rect 3283 10084 5672 10112
rect 6139 10084 6184 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10013 2283 10047
rect 2225 10007 2283 10013
rect 2240 9976 2268 10007
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3329 10047 3387 10053
rect 3329 10044 3341 10047
rect 3016 10016 3341 10044
rect 3016 10004 3022 10016
rect 3329 10013 3341 10016
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4154 9976 4160 9988
rect 2240 9948 4160 9976
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 4448 9908 4476 10007
rect 4798 9908 4804 9920
rect 2832 9880 2877 9908
rect 4448 9880 4804 9908
rect 2832 9868 2838 9880
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 5644 9908 5672 10084
rect 6172 10075 6184 10084
rect 6178 10072 6184 10075
rect 6236 10072 6242 10124
rect 7920 10115 7978 10121
rect 7920 10081 7932 10115
rect 7966 10112 7978 10115
rect 9766 10112 9772 10124
rect 7966 10084 9772 10112
rect 7966 10081 7978 10084
rect 7920 10075 7978 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10226 10112 10232 10124
rect 10091 10084 10232 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 10428 10112 10456 10152
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 10428 10084 11468 10112
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5776 10016 5917 10044
rect 5776 10004 5782 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 6972 10016 7665 10044
rect 6972 10004 6978 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 10376 10016 10421 10044
rect 10376 10004 10382 10016
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 11440 10053 11468 10084
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 11572 10084 13645 10112
rect 11572 10072 11578 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 14424 10084 14473 10112
rect 14424 10072 14430 10084
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 14461 10075 14519 10081
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 10744 10016 11345 10044
rect 10744 10004 10750 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 12434 10044 12440 10056
rect 11664 10016 12440 10044
rect 11664 10004 11670 10016
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 12713 10047 12771 10053
rect 12584 10016 12629 10044
rect 12584 10004 12590 10016
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 12802 10044 12808 10056
rect 12759 10016 12808 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13780 10016 13829 10044
rect 13780 10004 13786 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 9677 9979 9735 9985
rect 9677 9945 9689 9979
rect 9723 9976 9735 9979
rect 13630 9976 13636 9988
rect 9723 9948 13636 9976
rect 9723 9945 9735 9948
rect 9677 9939 9735 9945
rect 13630 9936 13636 9948
rect 13688 9936 13694 9988
rect 11054 9908 11060 9920
rect 5644 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 12032 9880 12081 9908
rect 12032 9868 12038 9880
rect 12069 9877 12081 9880
rect 12115 9877 12127 9911
rect 12069 9871 12127 9877
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 13044 9880 13277 9908
rect 13044 9868 13050 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 13265 9871 13323 9877
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 14424 9880 14657 9908
rect 14424 9868 14430 9880
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 14645 9871 14703 9877
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 5534 9704 5540 9716
rect 4816 9676 5540 9704
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 4065 9639 4123 9645
rect 4065 9636 4077 9639
rect 2648 9608 4077 9636
rect 2648 9596 2654 9608
rect 4065 9605 4077 9608
rect 4111 9605 4123 9639
rect 4816 9636 4844 9676
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 5684 9676 6285 9704
rect 5684 9664 5690 9676
rect 6273 9673 6285 9676
rect 6319 9673 6331 9707
rect 8665 9707 8723 9713
rect 6273 9667 6331 9673
rect 6840 9676 7788 9704
rect 6840 9636 6868 9676
rect 4065 9599 4123 9605
rect 4632 9608 4844 9636
rect 5920 9608 6868 9636
rect 7760 9636 7788 9676
rect 8665 9673 8677 9707
rect 8711 9704 8723 9707
rect 10594 9704 10600 9716
rect 8711 9676 10600 9704
rect 8711 9673 8723 9676
rect 8665 9667 8723 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 11054 9704 11060 9716
rect 11015 9676 11060 9704
rect 11054 9664 11060 9676
rect 11112 9664 11118 9716
rect 12158 9704 12164 9716
rect 11348 9676 12164 9704
rect 8570 9636 8576 9648
rect 7760 9608 8576 9636
rect 2958 9568 2964 9580
rect 2919 9540 2964 9568
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 3660 9540 3801 9568
rect 3660 9528 3666 9540
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4488 9540 4537 9568
rect 4488 9528 4494 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 4632 9500 4660 9608
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4755 9540 5028 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4890 9500 4896 9512
rect 2823 9472 4660 9500
rect 4851 9472 4896 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5000 9500 5028 9540
rect 5000 9472 5396 9500
rect 1394 9392 1400 9444
rect 1452 9432 1458 9444
rect 1857 9435 1915 9441
rect 1857 9432 1869 9435
rect 1452 9404 1869 9432
rect 1452 9392 1458 9404
rect 1857 9401 1869 9404
rect 1903 9401 1915 9435
rect 1857 9395 1915 9401
rect 2869 9435 2927 9441
rect 2869 9401 2881 9435
rect 2915 9432 2927 9435
rect 3510 9432 3516 9444
rect 2915 9404 3516 9432
rect 2915 9401 2927 9404
rect 2869 9395 2927 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 4062 9432 4068 9444
rect 3651 9404 4068 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 4062 9392 4068 9404
rect 4120 9392 4126 9444
rect 4246 9392 4252 9444
rect 4304 9432 4310 9444
rect 5166 9441 5172 9444
rect 4433 9435 4491 9441
rect 4433 9432 4445 9435
rect 4304 9404 4445 9432
rect 4304 9392 4310 9404
rect 4433 9401 4445 9404
rect 4479 9401 4491 9435
rect 5160 9432 5172 9441
rect 5127 9404 5172 9432
rect 4433 9395 4491 9401
rect 5160 9395 5172 9404
rect 5166 9392 5172 9395
rect 5224 9392 5230 9444
rect 5368 9432 5396 9472
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5920 9500 5948 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 9861 9639 9919 9645
rect 9861 9605 9873 9639
rect 9907 9636 9919 9639
rect 10686 9636 10692 9648
rect 9907 9608 10692 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 6822 9568 6828 9580
rect 6783 9540 6828 9568
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 9490 9568 9496 9580
rect 9355 9540 9496 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 9824 9540 10425 9568
rect 9824 9528 9830 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 5500 9472 5948 9500
rect 5500 9460 5506 9472
rect 6270 9460 6276 9512
rect 6328 9460 6334 9512
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 8478 9500 8484 9512
rect 6788 9472 8484 9500
rect 6788 9460 6794 9472
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9582 9500 9588 9512
rect 9079 9472 9588 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9500 10287 9503
rect 11348 9500 11376 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12253 9707 12311 9713
rect 12253 9673 12265 9707
rect 12299 9704 12311 9707
rect 14458 9704 14464 9716
rect 12299 9676 14464 9704
rect 12299 9673 12311 9676
rect 12253 9667 12311 9673
rect 14458 9664 14464 9676
rect 14516 9664 14522 9716
rect 11514 9596 11520 9648
rect 11572 9636 11578 9648
rect 11572 9608 13032 9636
rect 11572 9596 11578 9608
rect 13004 9580 13032 9608
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 11790 9568 11796 9580
rect 11747 9540 11796 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 11940 9540 12296 9568
rect 11940 9528 11946 9540
rect 10275 9472 11376 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 11422 9460 11428 9512
rect 11480 9460 11486 9512
rect 12268 9500 12296 9540
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12492 9540 12909 9568
rect 12492 9528 12498 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 13044 9540 13137 9568
rect 13044 9528 13050 9540
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13780 9540 14197 9568
rect 13780 9528 13786 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 14093 9503 14151 9509
rect 12268 9472 12848 9500
rect 6288 9432 6316 9460
rect 7098 9441 7104 9444
rect 5368 9404 6316 9432
rect 7092 9395 7104 9441
rect 7156 9432 7162 9444
rect 11440 9432 11468 9460
rect 12820 9441 12848 9472
rect 14093 9469 14105 9503
rect 14139 9500 14151 9503
rect 14642 9500 14648 9512
rect 14139 9472 14648 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 7156 9404 7192 9432
rect 9048 9404 11468 9432
rect 11517 9435 11575 9441
rect 7098 9392 7104 9395
rect 7156 9392 7162 9404
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 2096 9336 2421 9364
rect 2096 9324 2102 9336
rect 2409 9333 2421 9336
rect 2455 9333 2467 9367
rect 2409 9327 2467 9333
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 3200 9336 3249 9364
rect 3200 9324 3206 9336
rect 3237 9333 3249 9336
rect 3283 9333 3295 9367
rect 3237 9327 3295 9333
rect 3697 9367 3755 9373
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 4706 9364 4712 9376
rect 3743 9336 4712 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 7834 9364 7840 9376
rect 6420 9336 7840 9364
rect 6420 9324 6426 9336
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8202 9364 8208 9376
rect 8115 9336 8208 9364
rect 8202 9324 8208 9336
rect 8260 9364 8266 9376
rect 9048 9364 9076 9404
rect 11517 9401 11529 9435
rect 11563 9432 11575 9435
rect 12253 9435 12311 9441
rect 12253 9432 12265 9435
rect 11563 9404 12265 9432
rect 11563 9401 11575 9404
rect 11517 9395 11575 9401
rect 12253 9401 12265 9404
rect 12299 9401 12311 9435
rect 12253 9395 12311 9401
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 14182 9432 14188 9444
rect 12851 9404 14188 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 14182 9392 14188 9404
rect 14240 9432 14246 9444
rect 14844 9432 14872 9463
rect 14240 9404 14872 9432
rect 14240 9392 14246 9404
rect 8260 9336 9076 9364
rect 9125 9367 9183 9373
rect 8260 9324 8266 9336
rect 9125 9333 9137 9367
rect 9171 9364 9183 9367
rect 9306 9364 9312 9376
rect 9171 9336 9312 9364
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 10318 9364 10324 9376
rect 10279 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11425 9367 11483 9373
rect 11425 9364 11437 9367
rect 11388 9336 11437 9364
rect 11388 9324 11394 9336
rect 11425 9333 11437 9336
rect 11471 9333 11483 9367
rect 11425 9327 11483 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12526 9364 12532 9376
rect 12483 9336 12532 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13633 9367 13691 9373
rect 13633 9364 13645 9367
rect 13136 9336 13645 9364
rect 13136 9324 13142 9336
rect 13633 9333 13645 9336
rect 13679 9333 13691 9367
rect 13633 9327 13691 9333
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13872 9336 14013 9364
rect 13872 9324 13878 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 14001 9327 14059 9333
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 14332 9336 15025 9364
rect 14332 9324 14338 9336
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 15013 9327 15071 9333
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 1854 9160 1860 9172
rect 1627 9132 1860 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 5166 9160 5172 9172
rect 4396 9132 5172 9160
rect 4396 9120 4402 9132
rect 5166 9120 5172 9132
rect 5224 9160 5230 9172
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 5224 9132 5457 9160
rect 5224 9120 5230 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 6512 9132 7696 9160
rect 6512 9120 6518 9132
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 2774 9092 2780 9104
rect 1995 9064 2780 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 2774 9052 2780 9064
rect 2832 9052 2838 9104
rect 4890 9092 4896 9104
rect 4080 9064 4896 9092
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 3602 9024 3608 9036
rect 2648 8996 3608 9024
rect 2648 8984 2654 8996
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 4080 9033 4108 9064
rect 4890 9052 4896 9064
rect 4948 9052 4954 9104
rect 7098 9092 7104 9104
rect 5000 9064 7104 9092
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4321 9027 4379 9033
rect 4321 9024 4333 9027
rect 4212 8996 4333 9024
rect 4212 8984 4218 8996
rect 4321 8993 4333 8996
rect 4367 8993 4379 9027
rect 4321 8987 4379 8993
rect 4614 8984 4620 9036
rect 4672 9024 4678 9036
rect 5000 9024 5028 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 7668 9101 7696 9132
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9674 9160 9680 9172
rect 9272 9132 9680 9160
rect 9272 9120 9278 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 10008 9132 10057 9160
rect 10008 9120 10014 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 11882 9160 11888 9172
rect 10744 9132 11888 9160
rect 10744 9120 10750 9132
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 12115 9132 13737 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 7653 9095 7711 9101
rect 7653 9061 7665 9095
rect 7699 9092 7711 9095
rect 7834 9092 7840 9104
rect 7699 9064 7840 9092
rect 7699 9061 7711 9064
rect 7653 9055 7711 9061
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 8012 9095 8070 9101
rect 8012 9061 8024 9095
rect 8058 9092 8070 9095
rect 8202 9092 8208 9104
rect 8058 9064 8208 9092
rect 8058 9061 8070 9064
rect 8012 9055 8070 9061
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 13906 9092 13912 9104
rect 8720 9064 13912 9092
rect 8720 9052 8726 9064
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 4672 8996 5028 9024
rect 5905 9027 5963 9033
rect 4672 8984 4678 8996
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 9950 9024 9956 9036
rect 5951 8996 9956 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 11241 9027 11299 9033
rect 11241 8993 11253 9027
rect 11287 9024 11299 9027
rect 12158 9024 12164 9036
rect 11287 8996 12164 9024
rect 11287 8993 11299 8996
rect 11241 8987 11299 8993
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12437 9027 12495 9033
rect 12437 9024 12449 9027
rect 12400 8996 12449 9024
rect 12400 8984 12406 8996
rect 12437 8993 12449 8996
rect 12483 8993 12495 9027
rect 13630 9024 13636 9036
rect 13591 8996 13636 9024
rect 12437 8987 12495 8993
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 14458 9024 14464 9036
rect 14419 8996 14464 9024
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2240 8820 2268 8919
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 2924 8928 3249 8956
rect 2924 8916 2930 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 7742 8956 7748 8968
rect 7703 8928 7748 8956
rect 3421 8919 3479 8925
rect 2777 8891 2835 8897
rect 2777 8857 2789 8891
rect 2823 8888 2835 8891
rect 3326 8888 3332 8900
rect 2823 8860 3332 8888
rect 2823 8857 2835 8860
rect 2777 8851 2835 8857
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 3142 8820 3148 8832
rect 2240 8792 3148 8820
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3436 8820 3464 8919
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 10137 8959 10195 8965
rect 8904 8928 9996 8956
rect 8904 8916 8910 8928
rect 3786 8848 3792 8900
rect 3844 8888 3850 8900
rect 4062 8888 4068 8900
rect 3844 8860 4068 8888
rect 3844 8848 3850 8860
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 6270 8888 6276 8900
rect 5368 8860 6276 8888
rect 5368 8820 5396 8860
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 9766 8888 9772 8900
rect 9140 8860 9772 8888
rect 3436 8792 5396 8820
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 9140 8829 9168 8860
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 5684 8792 9137 8820
rect 5684 8780 5690 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 9674 8820 9680 8832
rect 9635 8792 9680 8820
rect 9125 8783 9183 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9968 8820 9996 8928
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10410 8956 10416 8968
rect 10367 8928 10416 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10042 8848 10048 8900
rect 10100 8888 10106 8900
rect 10152 8888 10180 8919
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 11330 8956 11336 8968
rect 10652 8928 11336 8956
rect 10652 8916 10658 8928
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 12526 8956 12532 8968
rect 11572 8928 11617 8956
rect 12487 8928 12532 8956
rect 11572 8916 11578 8928
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 12986 8956 12992 8968
rect 12759 8928 12992 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13780 8928 13829 8956
rect 13780 8916 13786 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 10778 8888 10784 8900
rect 10100 8860 10784 8888
rect 10100 8848 10106 8860
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8888 10931 8891
rect 12158 8888 12164 8900
rect 10919 8860 12164 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12342 8820 12348 8832
rect 9968 8792 12348 8820
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 13078 8780 13084 8832
rect 13136 8820 13142 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 13136 8792 13277 8820
rect 13136 8780 13142 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 13964 8792 14657 8820
rect 13964 8780 13970 8792
rect 14645 8789 14657 8792
rect 14691 8789 14703 8823
rect 14645 8783 14703 8789
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 4614 8616 4620 8628
rect 3200 8588 4620 8616
rect 3200 8576 3206 8588
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 6270 8616 6276 8628
rect 4764 8588 6132 8616
rect 6231 8588 6276 8616
rect 4764 8576 4770 8588
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 6104 8548 6132 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 8662 8616 8668 8628
rect 8623 8588 8668 8616
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 10042 8616 10048 8628
rect 8904 8588 10048 8616
rect 8904 8576 8910 8588
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 11057 8619 11115 8625
rect 11057 8616 11069 8619
rect 10192 8588 11069 8616
rect 10192 8576 10198 8588
rect 11057 8585 11069 8588
rect 11103 8585 11115 8619
rect 11057 8579 11115 8585
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 12437 8619 12495 8625
rect 12437 8616 12449 8619
rect 11204 8588 12449 8616
rect 11204 8576 11210 8588
rect 12437 8585 12449 8588
rect 12483 8585 12495 8619
rect 12437 8579 12495 8585
rect 12986 8576 12992 8628
rect 13044 8616 13050 8628
rect 13630 8616 13636 8628
rect 13044 8588 13400 8616
rect 13591 8588 13636 8616
rect 13044 8576 13050 8588
rect 6638 8548 6644 8560
rect 2648 8520 4844 8548
rect 6104 8520 6644 8548
rect 2648 8508 2654 8520
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 4246 8480 4252 8492
rect 3191 8452 4252 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4522 8480 4528 8492
rect 4387 8452 4528 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8412 1639 8415
rect 1762 8412 1768 8424
rect 1627 8384 1768 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 2774 8412 2780 8424
rect 1903 8384 2780 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8412 4123 8415
rect 4111 8384 4752 8412
rect 4111 8381 4123 8384
rect 4065 8375 4123 8381
rect 2866 8344 2872 8356
rect 2827 8316 2872 8344
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 3050 8304 3056 8356
rect 3108 8344 3114 8356
rect 4157 8347 4215 8353
rect 4157 8344 4169 8347
rect 3108 8316 4169 8344
rect 3108 8304 3114 8316
rect 4157 8313 4169 8316
rect 4203 8313 4215 8347
rect 4157 8307 4215 8313
rect 2498 8276 2504 8288
rect 2459 8248 2504 8276
rect 2498 8236 2504 8248
rect 2556 8236 2562 8288
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3697 8279 3755 8285
rect 3697 8245 3709 8279
rect 3743 8276 3755 8279
rect 3878 8276 3884 8288
rect 3743 8248 3884 8276
rect 3743 8245 3755 8248
rect 3697 8239 3755 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4724 8276 4752 8384
rect 4816 8344 4844 8520
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 8202 8548 8208 8560
rect 8115 8520 8208 8548
rect 8202 8508 8208 8520
rect 8260 8548 8266 8560
rect 8260 8520 11744 8548
rect 8260 8508 8266 8520
rect 9030 8440 9036 8492
rect 9088 8480 9094 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 9088 8452 9229 8480
rect 9088 8440 9094 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 10410 8480 10416 8492
rect 10371 8452 10416 8480
rect 9217 8443 9275 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11716 8489 11744 8520
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 11848 8520 13124 8548
rect 11848 8508 11854 8520
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11112 8452 11529 8480
rect 11112 8440 11118 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 11747 8452 11836 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8412 4951 8415
rect 5626 8412 5632 8424
rect 4939 8384 5632 8412
rect 4939 8381 4951 8384
rect 4893 8375 4951 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 9125 8415 9183 8421
rect 7024 8384 9076 8412
rect 5166 8353 5172 8356
rect 5160 8344 5172 8353
rect 4816 8316 5172 8344
rect 5160 8307 5172 8316
rect 5166 8304 5172 8307
rect 5224 8304 5230 8356
rect 7024 8344 7052 8384
rect 5276 8316 7052 8344
rect 7092 8347 7150 8353
rect 5276 8276 5304 8316
rect 7092 8313 7104 8347
rect 7138 8344 7150 8347
rect 8846 8344 8852 8356
rect 7138 8316 8852 8344
rect 7138 8313 7150 8316
rect 7092 8307 7150 8313
rect 8846 8304 8852 8316
rect 8904 8304 8910 8356
rect 9048 8344 9076 8384
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 10502 8412 10508 8424
rect 9171 8384 10508 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11808 8412 11836 8452
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 12342 8480 12348 8492
rect 11940 8452 12348 8480
rect 11940 8440 11946 8452
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13096 8489 13124 8520
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13262 8480 13268 8492
rect 13127 8452 13268 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13372 8480 13400 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 14458 8508 14464 8560
rect 14516 8548 14522 8560
rect 15013 8551 15071 8557
rect 15013 8548 15025 8551
rect 14516 8520 15025 8548
rect 14516 8508 14522 8520
rect 15013 8517 15025 8520
rect 15059 8517 15071 8551
rect 15013 8511 15071 8517
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 13372 8452 14197 8480
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 10836 8384 11560 8412
rect 11808 8384 12265 8412
rect 10836 8372 10842 8384
rect 9582 8344 9588 8356
rect 9048 8316 9588 8344
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 9766 8344 9772 8356
rect 9692 8316 9772 8344
rect 4724 8248 5304 8276
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 8662 8276 8668 8288
rect 5592 8248 8668 8276
rect 5592 8236 5598 8248
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 9033 8279 9091 8285
rect 9033 8245 9045 8279
rect 9079 8276 9091 8279
rect 9692 8276 9720 8316
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 10318 8344 10324 8356
rect 10279 8316 10324 8344
rect 10318 8304 10324 8316
rect 10376 8304 10382 8356
rect 11238 8344 11244 8356
rect 11072 8316 11244 8344
rect 9858 8276 9864 8288
rect 9079 8248 9720 8276
rect 9819 8248 9864 8276
rect 9079 8245 9091 8248
rect 9033 8239 9091 8245
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10229 8279 10287 8285
rect 10229 8245 10241 8279
rect 10275 8276 10287 8279
rect 11072 8276 11100 8316
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 11422 8344 11428 8356
rect 11383 8316 11428 8344
rect 11422 8304 11428 8316
rect 11480 8304 11486 8356
rect 11532 8344 11560 8384
rect 12253 8381 12265 8384
rect 12299 8381 12311 8415
rect 12360 8412 12388 8440
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12360 8384 12817 8412
rect 12253 8375 12311 8381
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 13170 8372 13176 8424
rect 13228 8412 13234 8424
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 13228 8384 14105 8412
rect 13228 8372 13234 8384
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14608 8384 14841 8412
rect 14608 8372 14614 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 13722 8344 13728 8356
rect 11532 8316 13728 8344
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 10275 8248 11100 8276
rect 12253 8279 12311 8285
rect 10275 8245 10287 8248
rect 10229 8239 10287 8245
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12710 8276 12716 8288
rect 12299 8248 12716 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14001 8279 14059 8285
rect 14001 8276 14013 8279
rect 13872 8248 14013 8276
rect 13872 8236 13878 8248
rect 14001 8245 14013 8248
rect 14047 8245 14059 8279
rect 14001 8239 14059 8245
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2682 8072 2688 8084
rect 1627 8044 2688 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2958 8072 2964 8084
rect 2823 8044 2964 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 9674 8072 9680 8084
rect 3068 8044 9680 8072
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 3068 8004 3096 8044
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10318 8072 10324 8084
rect 10091 8044 10324 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10318 8032 10324 8044
rect 10376 8072 10382 8084
rect 10502 8072 10508 8084
rect 10376 8044 10508 8072
rect 10376 8032 10382 8044
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 11238 8072 11244 8084
rect 11199 8044 11244 8072
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 12526 8072 12532 8084
rect 11379 8044 12532 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 2280 7976 3096 8004
rect 3145 8007 3203 8013
rect 2280 7964 2286 7976
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 9766 8004 9772 8016
rect 3191 7976 9772 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10137 8007 10195 8013
rect 10137 7973 10149 8007
rect 10183 8004 10195 8007
rect 10686 8004 10692 8016
rect 10183 7976 10692 8004
rect 10183 7973 10195 7976
rect 10137 7967 10195 7973
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 4430 7936 4436 7948
rect 1995 7908 4436 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4724 7908 4813 7936
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2590 7868 2596 7880
rect 2271 7840 2596 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 3234 7868 3240 7880
rect 3195 7840 3240 7868
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3786 7868 3792 7880
rect 3467 7840 3792 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 4724 7812 4752 7908
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 5626 7936 5632 7948
rect 5587 7908 5632 7936
rect 4801 7899 4859 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5896 7939 5954 7945
rect 5896 7936 5908 7939
rect 5736 7908 5908 7936
rect 4890 7868 4896 7880
rect 4851 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5736 7868 5764 7908
rect 5896 7905 5908 7908
rect 5942 7936 5954 7939
rect 6270 7936 6276 7948
rect 5942 7908 6276 7936
rect 5942 7905 5954 7908
rect 5896 7899 5954 7905
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 7558 7936 7564 7948
rect 7515 7908 7564 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 7736 7939 7794 7945
rect 7736 7905 7748 7939
rect 7782 7936 7794 7939
rect 8202 7936 8208 7948
rect 7782 7908 8208 7936
rect 7782 7905 7794 7908
rect 7736 7899 7794 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9214 7936 9220 7948
rect 8904 7908 9220 7936
rect 8904 7896 8910 7908
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9490 7936 9496 7948
rect 9451 7908 9496 7936
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 10870 7936 10876 7948
rect 10336 7908 10876 7936
rect 5123 7840 5764 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9180 7840 10241 7868
rect 9180 7828 9186 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 3016 7772 4568 7800
rect 3016 7760 3022 7772
rect 4430 7732 4436 7744
rect 4391 7704 4436 7732
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 4540 7732 4568 7772
rect 4706 7760 4712 7812
rect 4764 7760 4770 7812
rect 4982 7760 4988 7812
rect 5040 7800 5046 7812
rect 5442 7800 5448 7812
rect 5040 7772 5448 7800
rect 5040 7760 5046 7772
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 6564 7772 7135 7800
rect 5074 7732 5080 7744
rect 4540 7704 5080 7732
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5166 7692 5172 7744
rect 5224 7732 5230 7744
rect 6564 7732 6592 7772
rect 5224 7704 6592 7732
rect 5224 7692 5230 7704
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7009 7735 7067 7741
rect 7009 7732 7021 7735
rect 6972 7704 7021 7732
rect 6972 7692 6978 7704
rect 7009 7701 7021 7704
rect 7055 7701 7067 7735
rect 7107 7732 7135 7772
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 10336 7800 10364 7908
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11348 7936 11376 8035
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 12860 8044 13277 8072
rect 12860 8032 12866 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13722 8072 13728 8084
rect 13683 8044 13728 8072
rect 13265 8035 13323 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 11514 7964 11520 8016
rect 11572 8004 11578 8016
rect 12618 8004 12624 8016
rect 11572 7976 12624 8004
rect 11572 7964 11578 7976
rect 11296 7908 11376 7936
rect 11296 7896 11302 7908
rect 12158 7896 12164 7948
rect 12216 7936 12222 7948
rect 12544 7945 12572 7976
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 12437 7939 12495 7945
rect 12437 7936 12449 7939
rect 12216 7908 12449 7936
rect 12216 7896 12222 7908
rect 12437 7905 12449 7908
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7905 12587 7939
rect 12529 7899 12587 7905
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 12952 7908 13645 7936
rect 12952 7896 12958 7908
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 14461 7939 14519 7945
rect 14461 7905 14473 7939
rect 14507 7936 14519 7939
rect 14734 7936 14740 7948
rect 14507 7908 14740 7936
rect 14507 7905 14519 7908
rect 14461 7899 14519 7905
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 10744 7840 11437 7868
rect 10744 7828 10750 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 11664 7840 12725 7868
rect 11664 7828 11670 7840
rect 12713 7837 12725 7840
rect 12759 7868 12771 7871
rect 12759 7840 13216 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 8720 7772 10364 7800
rect 10873 7803 10931 7809
rect 8720 7760 8726 7772
rect 10873 7769 10885 7803
rect 10919 7800 10931 7803
rect 12802 7800 12808 7812
rect 10919 7772 11100 7800
rect 10919 7769 10931 7772
rect 10873 7763 10931 7769
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 7107 7704 8861 7732
rect 7009 7695 7067 7701
rect 8849 7701 8861 7704
rect 8895 7701 8907 7735
rect 9306 7732 9312 7744
rect 9267 7704 9312 7732
rect 8849 7695 8907 7701
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7732 9735 7735
rect 10962 7732 10968 7744
rect 9723 7704 10968 7732
rect 9723 7701 9735 7704
rect 9677 7695 9735 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11072 7732 11100 7772
rect 11624 7772 12808 7800
rect 11624 7732 11652 7772
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 13188 7800 13216 7840
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 13909 7871 13967 7877
rect 13909 7868 13921 7871
rect 13320 7840 13921 7868
rect 13320 7828 13326 7840
rect 13909 7837 13921 7840
rect 13955 7868 13967 7871
rect 14182 7868 14188 7880
rect 13955 7840 14188 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14458 7800 14464 7812
rect 13188 7772 14464 7800
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 11072 7704 11652 7732
rect 12069 7735 12127 7741
rect 12069 7701 12081 7735
rect 12115 7732 12127 7735
rect 13170 7732 13176 7744
rect 12115 7704 13176 7732
rect 12115 7701 12127 7704
rect 12069 7695 12127 7701
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 14642 7732 14648 7744
rect 14603 7704 14648 7732
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 2866 7528 2872 7540
rect 1903 7500 2872 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 9030 7528 9036 7540
rect 3292 7500 9036 7528
rect 3292 7488 3298 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11330 7528 11336 7540
rect 10928 7500 11336 7528
rect 10928 7488 10934 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 12434 7528 12440 7540
rect 12395 7500 12440 7528
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14826 7528 14832 7540
rect 14056 7500 14832 7528
rect 14056 7488 14062 7500
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 2314 7420 2320 7472
rect 2372 7460 2378 7472
rect 2958 7460 2964 7472
rect 2372 7432 2964 7460
rect 2372 7420 2378 7432
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 4433 7463 4491 7469
rect 4433 7429 4445 7463
rect 4479 7460 4491 7463
rect 4614 7460 4620 7472
rect 4479 7432 4620 7460
rect 4479 7429 4491 7432
rect 4433 7423 4491 7429
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 8202 7460 8208 7472
rect 8163 7432 8208 7460
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 10505 7463 10563 7469
rect 10505 7429 10517 7463
rect 10551 7429 10563 7463
rect 10505 7423 10563 7429
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 6822 7392 6828 7404
rect 2547 7364 3188 7392
rect 6783 7364 6828 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 3016 7296 3065 7324
rect 3016 7284 3022 7296
rect 3053 7293 3065 7296
rect 3099 7293 3111 7327
rect 3160 7324 3188 7364
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 8662 7392 8668 7404
rect 7892 7364 8668 7392
rect 7892 7352 7898 7364
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 10520 7392 10548 7423
rect 12710 7420 12716 7472
rect 12768 7460 12774 7472
rect 13262 7460 13268 7472
rect 12768 7432 13268 7460
rect 12768 7420 12774 7432
rect 10428 7364 10548 7392
rect 3786 7324 3792 7336
rect 3160 7296 3792 7324
rect 3053 7287 3111 7293
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4856 7296 4905 7324
rect 4856 7284 4862 7296
rect 4893 7293 4905 7296
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 5000 7296 8248 7324
rect 3326 7265 3332 7268
rect 3320 7256 3332 7265
rect 3287 7228 3332 7256
rect 3320 7219 3332 7228
rect 3326 7216 3332 7219
rect 3384 7216 3390 7268
rect 5000 7256 5028 7296
rect 5166 7265 5172 7268
rect 5160 7256 5172 7265
rect 3436 7228 5028 7256
rect 5079 7228 5172 7256
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 3436 7188 3464 7228
rect 5160 7219 5172 7228
rect 5224 7256 5230 7268
rect 5224 7228 6960 7256
rect 5166 7216 5172 7219
rect 5224 7216 5230 7228
rect 6932 7200 6960 7228
rect 7006 7216 7012 7268
rect 7064 7265 7070 7268
rect 7064 7259 7128 7265
rect 7064 7225 7082 7259
rect 7116 7225 7128 7259
rect 7064 7219 7128 7225
rect 7064 7216 7070 7219
rect 2363 7160 3464 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3786 7188 3792 7200
rect 3568 7160 3792 7188
rect 3568 7148 3574 7160
rect 3786 7148 3792 7160
rect 3844 7148 3850 7200
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 5442 7188 5448 7200
rect 4580 7160 5448 7188
rect 4580 7148 4586 7160
rect 5442 7148 5448 7160
rect 5500 7188 5506 7200
rect 6273 7191 6331 7197
rect 6273 7188 6285 7191
rect 5500 7160 6285 7188
rect 5500 7148 5506 7160
rect 6273 7157 6285 7160
rect 6319 7157 6331 7191
rect 6273 7151 6331 7157
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 8110 7188 8116 7200
rect 6972 7160 8116 7188
rect 6972 7148 6978 7160
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8220 7188 8248 7296
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 8921 7327 8979 7333
rect 8921 7324 8933 7327
rect 8812 7296 8933 7324
rect 8812 7284 8818 7296
rect 8921 7293 8933 7296
rect 8967 7293 8979 7327
rect 8921 7287 8979 7293
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10428 7324 10456 7364
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10778 7392 10784 7404
rect 10652 7364 10784 7392
rect 10652 7352 10658 7364
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11146 7392 11152 7404
rect 11107 7364 11152 7392
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12894 7392 12900 7404
rect 11747 7364 12900 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13004 7401 13032 7432
rect 13262 7420 13268 7432
rect 13320 7420 13326 7472
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 13228 7364 14105 7392
rect 13228 7352 13234 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14240 7364 14285 7392
rect 14240 7352 14246 7364
rect 9732 7296 10456 7324
rect 10873 7327 10931 7333
rect 9732 7284 9738 7296
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 12434 7324 12440 7336
rect 10919 7296 12440 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 15010 7324 15016 7336
rect 14875 7296 15016 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 11146 7256 11152 7268
rect 10612 7228 11152 7256
rect 9858 7188 9864 7200
rect 8220 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 10134 7188 10140 7200
rect 10091 7160 10140 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10612 7188 10640 7228
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 12710 7256 12716 7268
rect 12400 7228 12716 7256
rect 12400 7216 12406 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 12805 7259 12863 7265
rect 12805 7225 12817 7259
rect 12851 7256 12863 7259
rect 13170 7256 13176 7268
rect 12851 7228 13176 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 13170 7216 13176 7228
rect 13228 7256 13234 7268
rect 13538 7256 13544 7268
rect 13228 7228 13544 7256
rect 13228 7216 13234 7228
rect 13538 7216 13544 7228
rect 13596 7216 13602 7268
rect 10284 7160 10640 7188
rect 10284 7148 10290 7160
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 11756 7160 12909 7188
rect 11756 7148 11762 7160
rect 12897 7157 12909 7160
rect 12943 7188 12955 7191
rect 12986 7188 12992 7200
rect 12943 7160 12992 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 13630 7188 13636 7200
rect 13591 7160 13636 7188
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13998 7188 14004 7200
rect 13959 7160 14004 7188
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 14240 7160 15025 7188
rect 14240 7148 14246 7160
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 1946 6984 1952 6996
rect 1907 6956 1952 6984
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 2096 6956 7880 6984
rect 2096 6944 2102 6956
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 2682 6916 2688 6928
rect 2464 6888 2688 6916
rect 2464 6876 2470 6888
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 3145 6919 3203 6925
rect 3145 6885 3157 6919
rect 3191 6916 3203 6919
rect 3234 6916 3240 6928
rect 3191 6888 3240 6916
rect 3191 6885 3203 6888
rect 3145 6879 3203 6885
rect 3234 6876 3240 6888
rect 3292 6876 3298 6928
rect 4985 6919 5043 6925
rect 4985 6885 4997 6919
rect 5031 6916 5043 6919
rect 5534 6916 5540 6928
rect 5031 6888 5540 6916
rect 5031 6885 5043 6888
rect 4985 6879 5043 6885
rect 5534 6876 5540 6888
rect 5592 6876 5598 6928
rect 6086 6925 6092 6928
rect 6080 6879 6092 6925
rect 6144 6916 6150 6928
rect 6144 6888 6180 6916
rect 6086 6876 6092 6879
rect 6144 6876 6150 6888
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2087 6820 2728 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2700 6780 2728 6820
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 7558 6848 7564 6860
rect 2832 6820 7564 6848
rect 2832 6808 2838 6820
rect 3234 6780 3240 6792
rect 2700 6752 3096 6780
rect 3195 6752 3240 6780
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 3068 6712 3096 6752
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3344 6789 3372 6820
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 7742 6848 7748 6860
rect 7699 6820 7748 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 7852 6848 7880 6956
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 10226 6984 10232 6996
rect 8168 6956 10232 6984
rect 8168 6944 8174 6956
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 12526 6984 12532 6996
rect 10560 6956 12532 6984
rect 10560 6944 10566 6956
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 12860 6956 13185 6984
rect 12860 6944 12866 6956
rect 13173 6953 13185 6956
rect 13219 6953 13231 6987
rect 13173 6947 13231 6953
rect 13909 6987 13967 6993
rect 13909 6953 13921 6987
rect 13955 6984 13967 6987
rect 13998 6984 14004 6996
rect 13955 6956 14004 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 7920 6919 7978 6925
rect 7920 6885 7932 6919
rect 7966 6916 7978 6919
rect 8202 6916 8208 6928
rect 7966 6888 8208 6916
rect 7966 6885 7978 6888
rect 7920 6879 7978 6885
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 8662 6876 8668 6928
rect 8720 6916 8726 6928
rect 9944 6919 10002 6925
rect 8720 6888 9720 6916
rect 8720 6876 8726 6888
rect 9692 6857 9720 6888
rect 9944 6885 9956 6919
rect 9990 6916 10002 6919
rect 10134 6916 10140 6928
rect 9990 6888 10140 6916
rect 9990 6885 10002 6888
rect 9944 6879 10002 6885
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 10778 6876 10784 6928
rect 10836 6916 10842 6928
rect 11698 6916 11704 6928
rect 10836 6888 11704 6916
rect 10836 6876 10842 6888
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 11885 6919 11943 6925
rect 11885 6885 11897 6919
rect 11931 6916 11943 6919
rect 12158 6916 12164 6928
rect 11931 6888 12164 6916
rect 11931 6885 11943 6888
rect 11885 6879 11943 6885
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 13078 6916 13084 6928
rect 13039 6888 13084 6916
rect 13078 6876 13084 6888
rect 13136 6876 13142 6928
rect 9677 6851 9735 6857
rect 7852 6820 9168 6848
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 5074 6780 5080 6792
rect 3568 6752 4752 6780
rect 5035 6752 5080 6780
rect 3568 6740 3574 6752
rect 4430 6712 4436 6724
rect 1627 6684 3004 6712
rect 3068 6684 4436 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2096 6616 2789 6644
rect 2096 6604 2102 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2976 6644 3004 6684
rect 4430 6672 4436 6684
rect 4488 6672 4494 6724
rect 3050 6644 3056 6656
rect 2976 6616 3056 6644
rect 2777 6607 2835 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 3200 6616 4629 6644
rect 3200 6604 3206 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 4724 6644 4752 6752
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5534 6780 5540 6792
rect 5307 6752 5540 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 5626 6712 5632 6724
rect 4856 6684 5632 6712
rect 4856 6672 4862 6684
rect 5626 6672 5632 6684
rect 5684 6712 5690 6724
rect 5828 6712 5856 6743
rect 5684 6684 5856 6712
rect 6748 6684 7328 6712
rect 5684 6672 5690 6684
rect 6748 6644 6776 6684
rect 7190 6644 7196 6656
rect 4724 6616 6776 6644
rect 7151 6616 7196 6644
rect 4617 6607 4675 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7300 6644 7328 6684
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 7300 6616 9045 6644
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9140 6644 9168 6820
rect 9677 6817 9689 6851
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 9784 6820 12112 6848
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9784 6780 9812 6820
rect 9456 6752 9812 6780
rect 9456 6740 9462 6752
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 12084 6789 12112 6820
rect 12434 6808 12440 6860
rect 12492 6808 12498 6860
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 12676 6820 13492 6848
rect 12676 6808 12682 6820
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11664 6752 11989 6780
rect 11664 6740 11670 6752
rect 11977 6749 11989 6752
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6749 12127 6783
rect 12452 6780 12480 6808
rect 12986 6780 12992 6792
rect 12452 6752 12992 6780
rect 12069 6743 12127 6749
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13464 6780 13492 6820
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14056 6820 14289 6848
rect 14056 6808 14062 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 13464 6752 14381 6780
rect 13357 6743 13415 6749
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 10980 6684 12725 6712
rect 10980 6644 11008 6684
rect 12713 6681 12725 6684
rect 12759 6681 12771 6715
rect 12713 6675 12771 6681
rect 13262 6672 13268 6724
rect 13320 6712 13326 6724
rect 13372 6712 13400 6743
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 14516 6752 14561 6780
rect 14516 6740 14522 6752
rect 13722 6712 13728 6724
rect 13320 6684 13728 6712
rect 13320 6672 13326 6684
rect 13722 6672 13728 6684
rect 13780 6672 13786 6724
rect 9140 6616 11008 6644
rect 11057 6647 11115 6653
rect 9033 6607 9091 6613
rect 11057 6613 11069 6647
rect 11103 6644 11115 6647
rect 11330 6644 11336 6656
rect 11103 6616 11336 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 11517 6647 11575 6653
rect 11517 6613 11529 6647
rect 11563 6644 11575 6647
rect 12894 6644 12900 6656
rect 11563 6616 12900 6644
rect 11563 6613 11575 6616
rect 11517 6607 11575 6613
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 1854 6440 1860 6452
rect 1815 6412 1860 6440
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 5166 6440 5172 6452
rect 2280 6412 5172 6440
rect 2280 6400 2286 6412
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 7248 6412 7788 6440
rect 7248 6400 7254 6412
rect 4246 6332 4252 6384
rect 4304 6372 4310 6384
rect 4433 6375 4491 6381
rect 4433 6372 4445 6375
rect 4304 6344 4445 6372
rect 4304 6332 4310 6344
rect 4433 6341 4445 6344
rect 4479 6341 4491 6375
rect 7760 6372 7788 6412
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 10042 6440 10048 6452
rect 8260 6412 9904 6440
rect 10003 6412 10048 6440
rect 8260 6400 8266 6412
rect 8478 6372 8484 6384
rect 7760 6344 8484 6372
rect 4433 6335 4491 6341
rect 2222 6264 2228 6316
rect 2280 6304 2286 6316
rect 2409 6307 2467 6313
rect 2409 6304 2421 6307
rect 2280 6276 2421 6304
rect 2280 6264 2286 6276
rect 2409 6273 2421 6276
rect 2455 6273 2467 6307
rect 4448 6304 4476 6335
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 9876 6372 9904 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10505 6443 10563 6449
rect 10505 6409 10517 6443
rect 10551 6440 10563 6443
rect 10962 6440 10968 6452
rect 10551 6412 10968 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 12437 6443 12495 6449
rect 11072 6412 11836 6440
rect 10410 6372 10416 6384
rect 8588 6344 8708 6372
rect 9876 6344 10416 6372
rect 2409 6267 2467 6273
rect 2884 6276 3188 6304
rect 4448 6276 5028 6304
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 2884 6236 2912 6276
rect 2363 6208 2912 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 3016 6208 3065 6236
rect 3016 6196 3022 6208
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3160 6236 3188 6276
rect 3786 6236 3792 6248
rect 3160 6208 3792 6236
rect 3053 6199 3111 6205
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 2225 6103 2283 6109
rect 2225 6100 2237 6103
rect 2188 6072 2237 6100
rect 2188 6060 2194 6072
rect 2225 6069 2237 6072
rect 2271 6069 2283 6103
rect 3068 6100 3096 6199
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4856 6208 4905 6236
rect 4856 6196 4862 6208
rect 4893 6205 4905 6208
rect 4939 6205 4951 6239
rect 5000 6236 5028 6276
rect 8588 6248 8616 6344
rect 8680 6313 8708 6344
rect 10410 6332 10416 6344
rect 10468 6372 10474 6384
rect 11072 6372 11100 6412
rect 10468 6344 11100 6372
rect 10468 6332 10474 6344
rect 8672 6307 8730 6313
rect 8672 6273 8684 6307
rect 8718 6273 8730 6307
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 8672 6267 8730 6273
rect 10336 6276 11069 6304
rect 10336 6248 10364 6276
rect 11057 6273 11069 6276
rect 11103 6304 11115 6307
rect 11698 6304 11704 6316
rect 11103 6276 11704 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11808 6304 11836 6412
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 12526 6440 12532 6452
rect 12483 6412 12532 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 13722 6332 13728 6384
rect 13780 6372 13786 6384
rect 13780 6344 14228 6372
rect 13780 6332 13786 6344
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 11808 6276 13093 6304
rect 13081 6273 13093 6276
rect 13127 6304 13139 6307
rect 13354 6304 13360 6316
rect 13127 6276 13360 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 14200 6313 14228 6344
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 15010 6304 15016 6316
rect 14516 6276 15016 6304
rect 14516 6264 14522 6276
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 6822 6236 6828 6248
rect 5000 6208 6408 6236
rect 6735 6208 6828 6236
rect 4893 6199 4951 6205
rect 3326 6177 3332 6180
rect 3320 6168 3332 6177
rect 3287 6140 3332 6168
rect 3320 6131 3332 6140
rect 3326 6128 3332 6131
rect 3384 6128 3390 6180
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 5166 6177 5172 6180
rect 5160 6168 5172 6177
rect 4028 6140 5028 6168
rect 5127 6140 5172 6168
rect 4028 6128 4034 6140
rect 4798 6100 4804 6112
rect 3068 6072 4804 6100
rect 2225 6063 2283 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5000 6100 5028 6140
rect 5160 6131 5172 6140
rect 5166 6128 5172 6131
rect 5224 6128 5230 6180
rect 6086 6128 6092 6180
rect 6144 6128 6150 6180
rect 6104 6100 6132 6128
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 5000 6072 6285 6100
rect 6273 6069 6285 6072
rect 6319 6069 6331 6103
rect 6380 6100 6408 6208
rect 6822 6196 6828 6208
rect 6880 6236 6886 6248
rect 8570 6236 8576 6248
rect 6880 6208 8576 6236
rect 6880 6196 6886 6208
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 10318 6236 10324 6248
rect 8812 6208 10324 6236
rect 8812 6196 8818 6208
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 10870 6236 10876 6248
rect 10831 6208 10876 6236
rect 10870 6196 10876 6208
rect 10928 6236 10934 6248
rect 13722 6236 13728 6248
rect 10928 6208 13728 6236
rect 10928 6196 10934 6208
rect 13722 6196 13728 6208
rect 13780 6236 13786 6248
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 13780 6208 14841 6236
rect 13780 6196 13786 6208
rect 14829 6205 14841 6208
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 7098 6177 7104 6180
rect 7092 6168 7104 6177
rect 7059 6140 7104 6168
rect 7092 6131 7104 6140
rect 7098 6128 7104 6131
rect 7156 6128 7162 6180
rect 8910 6171 8968 6177
rect 8910 6168 8922 6171
rect 7208 6140 8922 6168
rect 7208 6100 7236 6140
rect 8910 6137 8922 6140
rect 8956 6137 8968 6171
rect 10778 6168 10784 6180
rect 8910 6131 8968 6137
rect 9784 6140 10784 6168
rect 6380 6072 7236 6100
rect 6273 6063 6331 6069
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 7800 6072 8217 6100
rect 7800 6060 7806 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8205 6063 8263 6069
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 9784 6100 9812 6140
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 10980 6140 11836 6168
rect 8720 6072 9812 6100
rect 8720 6060 8726 6072
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10980 6109 11008 6140
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 9916 6072 10977 6100
rect 9916 6060 9922 6072
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 10965 6063 11023 6069
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11296 6072 11713 6100
rect 11296 6060 11302 6072
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11808 6100 11836 6140
rect 12618 6128 12624 6180
rect 12676 6128 12682 6180
rect 12894 6168 12900 6180
rect 12855 6140 12900 6168
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 13262 6128 13268 6180
rect 13320 6168 13326 6180
rect 14001 6171 14059 6177
rect 14001 6168 14013 6171
rect 13320 6140 14013 6168
rect 13320 6128 13326 6140
rect 14001 6137 14013 6140
rect 14047 6137 14059 6171
rect 14001 6131 14059 6137
rect 12636 6100 12664 6128
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 11808 6072 12817 6100
rect 11701 6063 11759 6069
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13170 6100 13176 6112
rect 13044 6072 13176 6100
rect 13044 6060 13050 6072
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 13633 6103 13691 6109
rect 13633 6100 13645 6103
rect 13504 6072 13645 6100
rect 13504 6060 13510 6072
rect 13633 6069 13645 6072
rect 13679 6069 13691 6103
rect 13633 6063 13691 6069
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 13872 6072 14105 6100
rect 13872 6060 13878 6072
rect 14093 6069 14105 6072
rect 14139 6069 14151 6103
rect 15010 6100 15016 6112
rect 14971 6072 15016 6100
rect 14093 6063 14151 6069
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 2038 5896 2044 5908
rect 1999 5868 2044 5896
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 5166 5896 5172 5908
rect 3476 5868 5172 5896
rect 3476 5856 3482 5868
rect 5166 5856 5172 5868
rect 5224 5896 5230 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 5224 5868 8493 5896
rect 5224 5856 5230 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 8941 5899 8999 5905
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 10226 5896 10232 5908
rect 8987 5868 10232 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 12342 5896 12348 5908
rect 11624 5868 12020 5896
rect 12303 5868 12348 5896
rect 1949 5831 2007 5837
rect 1949 5797 1961 5831
rect 1995 5828 2007 5831
rect 11330 5828 11336 5840
rect 1995 5800 11336 5828
rect 1995 5797 2007 5800
rect 1949 5791 2007 5797
rect 11330 5788 11336 5800
rect 11388 5788 11394 5840
rect 11624 5828 11652 5868
rect 11992 5828 12020 5868
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 12860 5868 13553 5896
rect 12860 5856 12866 5868
rect 13541 5865 13553 5868
rect 13587 5865 13599 5899
rect 13541 5859 13599 5865
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 13998 5896 14004 5908
rect 13780 5868 14004 5896
rect 13780 5856 13786 5868
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 11440 5800 11652 5828
rect 11716 5800 11928 5828
rect 11992 5800 12296 5828
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 4479 5732 4660 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 3234 5692 3240 5704
rect 3195 5664 3240 5692
rect 2225 5655 2283 5661
rect 1946 5584 1952 5636
rect 2004 5624 2010 5636
rect 2130 5624 2136 5636
rect 2004 5596 2136 5624
rect 2004 5584 2010 5596
rect 2130 5584 2136 5596
rect 2188 5584 2194 5636
rect 2240 5624 2268 5655
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 3418 5692 3424 5704
rect 3379 5664 3424 5692
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 4522 5692 4528 5704
rect 4483 5664 4528 5692
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4430 5624 4436 5636
rect 2240 5596 4436 5624
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 2958 5556 2964 5568
rect 2823 5528 2964 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4632 5556 4660 5732
rect 4798 5720 4804 5772
rect 4856 5760 4862 5772
rect 5528 5763 5586 5769
rect 4856 5732 5304 5760
rect 4856 5720 4862 5732
rect 5276 5704 5304 5732
rect 5528 5729 5540 5763
rect 5574 5760 5586 5763
rect 6270 5760 6276 5772
rect 5574 5732 6276 5760
rect 5574 5729 5586 5732
rect 5528 5723 5586 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 7098 5760 7104 5772
rect 7059 5732 7104 5760
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7374 5769 7380 5772
rect 7357 5763 7380 5769
rect 7357 5760 7369 5763
rect 7208 5732 7369 5760
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 5166 5692 5172 5704
rect 4755 5664 5172 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 5316 5664 5361 5692
rect 5316 5652 5322 5664
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 7208 5692 7236 5732
rect 7357 5729 7369 5732
rect 7432 5760 7438 5772
rect 7432 5732 7505 5760
rect 7357 5723 7380 5729
rect 7374 5720 7380 5723
rect 7432 5720 7438 5732
rect 7650 5720 7656 5772
rect 7708 5760 7714 5772
rect 7708 5732 8156 5760
rect 7708 5720 7714 5732
rect 8128 5704 8156 5732
rect 8202 5720 8208 5772
rect 8260 5760 8266 5772
rect 9490 5760 9496 5772
rect 8260 5732 9496 5760
rect 8260 5720 8266 5732
rect 9490 5720 9496 5732
rect 9548 5760 9554 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9548 5732 9689 5760
rect 9548 5720 9554 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 11440 5760 11468 5800
rect 9677 5723 9735 5729
rect 9876 5732 11468 5760
rect 11517 5763 11575 5769
rect 6696 5664 7236 5692
rect 6696 5652 6702 5664
rect 8110 5652 8116 5704
rect 8168 5692 8174 5704
rect 9876 5692 9904 5732
rect 11517 5729 11529 5763
rect 11563 5760 11575 5763
rect 11716 5760 11744 5800
rect 11563 5732 11744 5760
rect 11900 5760 11928 5800
rect 12158 5760 12164 5772
rect 11900 5732 12164 5760
rect 11563 5729 11575 5732
rect 11517 5723 11575 5729
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 8168 5664 9904 5692
rect 8168 5652 8174 5664
rect 9950 5652 9956 5704
rect 10008 5692 10014 5704
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 10008 5664 10057 5692
rect 10008 5652 10014 5664
rect 10045 5661 10057 5664
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11606 5692 11612 5704
rect 11020 5664 11612 5692
rect 11020 5652 11026 5664
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11716 5664 11805 5692
rect 11716 5636 11744 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 12268 5692 12296 5800
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 12952 5800 14964 5828
rect 12952 5788 12958 5800
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 12584 5732 12725 5760
rect 12584 5720 12590 5732
rect 12713 5729 12725 5732
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 12860 5732 12905 5760
rect 12860 5720 12866 5732
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 14936 5769 14964 5800
rect 13909 5763 13967 5769
rect 13909 5760 13921 5763
rect 13044 5732 13921 5760
rect 13044 5720 13050 5732
rect 13909 5729 13921 5732
rect 13955 5729 13967 5763
rect 13909 5723 13967 5729
rect 14921 5763 14979 5769
rect 14921 5729 14933 5763
rect 14967 5729 14979 5763
rect 14921 5723 14979 5729
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12268 5664 12909 5692
rect 11793 5655 11851 5661
rect 12897 5661 12909 5664
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 13354 5652 13360 5704
rect 13412 5692 13418 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13412 5664 14105 5692
rect 13412 5652 13418 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 6564 5596 7144 5624
rect 6564 5556 6592 5596
rect 4632 5528 6592 5556
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 6914 5556 6920 5568
rect 6687 5528 6920 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7116 5556 7144 5596
rect 8202 5584 8208 5636
rect 8260 5624 8266 5636
rect 10870 5624 10876 5636
rect 8260 5596 10876 5624
rect 8260 5584 8266 5596
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 11698 5584 11704 5636
rect 11756 5584 11762 5636
rect 10410 5556 10416 5568
rect 7116 5528 10416 5556
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 11238 5556 11244 5568
rect 11195 5528 11244 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 14737 5559 14795 5565
rect 14737 5556 14749 5559
rect 12400 5528 14749 5556
rect 12400 5516 12406 5528
rect 14737 5525 14749 5528
rect 14783 5525 14795 5559
rect 14737 5519 14795 5525
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 3326 5352 3332 5364
rect 2516 5324 3332 5352
rect 2516 5225 2544 5324
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 4430 5352 4436 5364
rect 4343 5324 4436 5352
rect 4430 5312 4436 5324
rect 4488 5352 4494 5364
rect 9766 5352 9772 5364
rect 4488 5324 7880 5352
rect 4488 5312 4494 5324
rect 2590 5244 2596 5296
rect 2648 5284 2654 5296
rect 2648 5256 3096 5284
rect 2648 5244 2654 5256
rect 3068 5225 3096 5256
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5185 2559 5219
rect 2501 5179 2559 5185
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5185 3111 5219
rect 7852 5216 7880 5324
rect 8220 5324 9772 5352
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 8220 5293 8248 5324
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10134 5352 10140 5364
rect 9876 5324 10140 5352
rect 8205 5287 8263 5293
rect 8205 5284 8217 5287
rect 8076 5256 8217 5284
rect 8076 5244 8082 5256
rect 8205 5253 8217 5256
rect 8251 5253 8263 5287
rect 8205 5247 8263 5253
rect 8386 5244 8392 5296
rect 8444 5284 8450 5296
rect 8444 5256 8708 5284
rect 8444 5244 8450 5256
rect 8680 5225 8708 5256
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9876 5284 9904 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 12342 5352 12348 5364
rect 10928 5324 12348 5352
rect 10928 5312 10934 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13228 5324 13645 5352
rect 13228 5312 13234 5324
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 13633 5315 13691 5321
rect 9732 5256 9904 5284
rect 9732 5244 9738 5256
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 10045 5287 10103 5293
rect 10045 5284 10057 5287
rect 10008 5256 10057 5284
rect 10008 5244 10014 5256
rect 10045 5253 10057 5256
rect 10091 5253 10103 5287
rect 12437 5287 12495 5293
rect 10045 5247 10103 5253
rect 10428 5256 11376 5284
rect 8665 5219 8723 5225
rect 7852 5188 8616 5216
rect 3053 5179 3111 5185
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 3309 5151 3367 5157
rect 3309 5148 3321 5151
rect 2832 5120 3321 5148
rect 2832 5108 2838 5120
rect 3309 5117 3321 5120
rect 3355 5117 3367 5151
rect 3309 5111 3367 5117
rect 3602 5108 3608 5160
rect 3660 5148 3666 5160
rect 4798 5148 4804 5160
rect 3660 5120 4804 5148
rect 3660 5108 3666 5120
rect 4798 5108 4804 5120
rect 4856 5148 4862 5160
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 4856 5120 4905 5148
rect 4856 5108 4862 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 6454 5148 6460 5160
rect 4893 5111 4951 5117
rect 5000 5120 6460 5148
rect 2225 5083 2283 5089
rect 2225 5049 2237 5083
rect 2271 5080 2283 5083
rect 3786 5080 3792 5092
rect 2271 5052 3792 5080
rect 2271 5049 2283 5052
rect 2225 5043 2283 5049
rect 3786 5040 3792 5052
rect 3844 5040 3850 5092
rect 4430 5040 4436 5092
rect 4488 5080 4494 5092
rect 5000 5080 5028 5120
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 8386 5148 8392 5160
rect 6871 5120 8392 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 5166 5089 5172 5092
rect 5160 5080 5172 5089
rect 4488 5052 5028 5080
rect 5127 5052 5172 5080
rect 4488 5040 4494 5052
rect 5160 5043 5172 5052
rect 5166 5040 5172 5043
rect 5224 5040 5230 5092
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 6638 5080 6644 5092
rect 5592 5052 6644 5080
rect 5592 5040 5598 5052
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 2317 5015 2375 5021
rect 2317 4981 2329 5015
rect 2363 5012 2375 5015
rect 5718 5012 5724 5024
rect 2363 4984 5724 5012
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6840 5012 6868 5111
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8588 5148 8616 5188
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 10134 5216 10140 5228
rect 8665 5179 8723 5185
rect 9692 5188 10140 5216
rect 8921 5151 8979 5157
rect 8921 5148 8933 5151
rect 8588 5120 8933 5148
rect 8921 5117 8933 5120
rect 8967 5117 8979 5151
rect 8921 5111 8979 5117
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 7092 5083 7150 5089
rect 7092 5080 7104 5083
rect 6972 5052 7104 5080
rect 6972 5040 6978 5052
rect 7092 5049 7104 5052
rect 7138 5080 7150 5083
rect 9692 5080 9720 5188
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10428 5148 10456 5256
rect 11146 5216 11152 5228
rect 11107 5188 11152 5216
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 7138 5052 9720 5080
rect 9968 5120 10456 5148
rect 7138 5049 7150 5052
rect 7092 5043 7150 5049
rect 7190 5012 7196 5024
rect 6840 4984 7196 5012
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 9968 5012 9996 5120
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 11348 5148 11376 5256
rect 12437 5253 12449 5287
rect 12483 5284 12495 5287
rect 12618 5284 12624 5296
rect 12483 5256 12624 5284
rect 12483 5253 12495 5256
rect 12437 5247 12495 5253
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 13872 5256 14872 5284
rect 13872 5244 13878 5256
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 11480 5188 12909 5216
rect 11480 5176 11486 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 11606 5148 11612 5160
rect 11020 5120 11065 5148
rect 11348 5120 11612 5148
rect 11020 5108 11026 5120
rect 11606 5108 11612 5120
rect 11664 5148 11670 5160
rect 11664 5120 12940 5148
rect 11664 5108 11670 5120
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 10873 5083 10931 5089
rect 10873 5080 10885 5083
rect 10284 5052 10885 5080
rect 10284 5040 10290 5052
rect 10873 5049 10885 5052
rect 10919 5080 10931 5083
rect 11330 5080 11336 5092
rect 10919 5052 11336 5080
rect 10919 5049 10931 5052
rect 10873 5043 10931 5049
rect 11330 5040 11336 5052
rect 11388 5040 11394 5092
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 12492 5052 12817 5080
rect 12492 5040 12498 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12912 5080 12940 5120
rect 12986 5080 12992 5092
rect 12899 5052 12992 5080
rect 12805 5043 12863 5049
rect 12986 5040 12992 5052
rect 13044 5080 13050 5092
rect 13096 5080 13124 5179
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13228 5188 14197 5216
rect 13228 5176 13234 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14090 5148 14096 5160
rect 14047 5120 14096 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 14844 5157 14872 5256
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 13044 5052 13124 5080
rect 13044 5040 13050 5052
rect 13538 5040 13544 5092
rect 13596 5080 13602 5092
rect 14550 5080 14556 5092
rect 13596 5052 14556 5080
rect 13596 5040 13602 5052
rect 14550 5040 14556 5052
rect 14608 5040 14614 5092
rect 10502 5012 10508 5024
rect 7800 4984 9996 5012
rect 10463 4984 10508 5012
rect 7800 4972 7806 4984
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 11146 4972 11152 5024
rect 11204 5012 11210 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11204 4984 11713 5012
rect 11204 4972 11210 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 14090 5012 14096 5024
rect 14051 4984 14096 5012
rect 11701 4975 11759 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 15010 5012 15016 5024
rect 14971 4984 15016 5012
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 6638 4808 6644 4820
rect 2087 4780 6644 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 6972 4780 8677 4808
rect 6972 4768 6978 4780
rect 8665 4777 8677 4780
rect 8711 4808 8723 4811
rect 9674 4808 9680 4820
rect 8711 4780 9680 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10091 4780 11376 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 11348 4740 11376 4780
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 11480 4780 12081 4808
rect 11480 4768 11486 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 12069 4771 12127 4777
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 12860 4780 13277 4808
rect 12860 4768 12866 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13630 4808 13636 4820
rect 13543 4780 13636 4808
rect 13265 4771 13323 4777
rect 13630 4768 13636 4780
rect 13688 4808 13694 4820
rect 14182 4808 14188 4820
rect 13688 4780 14188 4808
rect 13688 4768 13694 4780
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 3344 4712 10916 4740
rect 11348 4712 12204 4740
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 2038 4672 2044 4684
rect 1995 4644 2044 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 3145 4675 3203 4681
rect 3145 4672 3157 4675
rect 3108 4644 3157 4672
rect 3108 4632 3114 4644
rect 3145 4641 3157 4644
rect 3191 4641 3203 4675
rect 3145 4635 3203 4641
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3344 4672 3372 4712
rect 4614 4672 4620 4684
rect 3283 4644 3372 4672
rect 4575 4644 4620 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 4755 4644 5212 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4604 2283 4607
rect 2271 4576 3372 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 1581 4539 1639 4545
rect 1581 4505 1593 4539
rect 1627 4536 1639 4539
rect 3234 4536 3240 4548
rect 1627 4508 3240 4536
rect 1627 4505 1639 4508
rect 1581 4499 1639 4505
rect 3234 4496 3240 4508
rect 3292 4496 3298 4548
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3344 4468 3372 4576
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 3476 4576 3521 4604
rect 3476 4564 3482 4576
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 4724 4604 4752 4635
rect 4890 4604 4896 4616
rect 3752 4576 4752 4604
rect 4803 4576 4896 4604
rect 3752 4564 3758 4576
rect 4890 4564 4896 4576
rect 4948 4604 4954 4616
rect 5184 4604 5212 4644
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5316 4644 5457 4672
rect 5316 4632 5322 4644
rect 5445 4641 5457 4644
rect 5491 4641 5503 4675
rect 5445 4635 5503 4641
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 5701 4675 5759 4681
rect 5701 4672 5713 4675
rect 5592 4644 5713 4672
rect 5592 4632 5598 4644
rect 5701 4641 5713 4644
rect 5747 4641 5759 4675
rect 5701 4635 5759 4641
rect 7552 4675 7610 4681
rect 7552 4641 7564 4675
rect 7598 4672 7610 4675
rect 8294 4672 8300 4684
rect 7598 4644 8300 4672
rect 7598 4641 7610 4644
rect 7552 4635 7610 4641
rect 8294 4632 8300 4644
rect 8352 4672 8358 4684
rect 9306 4672 9312 4684
rect 8352 4644 8616 4672
rect 9267 4644 9312 4672
rect 8352 4632 8358 4644
rect 4948 4576 5120 4604
rect 5184 4576 5304 4604
rect 4948 4564 4954 4576
rect 4154 4468 4160 4480
rect 2832 4440 2877 4468
rect 3344 4440 4160 4468
rect 2832 4428 2838 4440
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 4614 4468 4620 4480
rect 4295 4440 4620 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 5092 4468 5120 4576
rect 5276 4548 5304 4576
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 7248 4576 7297 4604
rect 7248 4564 7254 4576
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 5258 4496 5264 4548
rect 5316 4496 5322 4548
rect 8588 4536 8616 4644
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 10686 4672 10692 4684
rect 9824 4644 10692 4672
rect 9824 4632 9830 4644
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9582 4604 9588 4616
rect 8812 4576 9588 4604
rect 8812 4564 8818 4576
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9640 4576 10149 4604
rect 9640 4564 9646 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 8588 4508 9260 4536
rect 5626 4468 5632 4480
rect 5092 4440 5632 4468
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 6822 4468 6828 4480
rect 6144 4440 6828 4468
rect 6144 4428 6150 4440
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 9122 4468 9128 4480
rect 9083 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9232 4468 9260 4508
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 9732 4508 9777 4536
rect 9732 4496 9738 4508
rect 10244 4468 10272 4567
rect 10888 4545 10916 4712
rect 12176 4684 12204 4712
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 12437 4743 12495 4749
rect 12437 4740 12449 4743
rect 12400 4712 12449 4740
rect 12400 4700 12406 4712
rect 12437 4709 12449 4712
rect 12483 4709 12495 4743
rect 12437 4703 12495 4709
rect 12529 4743 12587 4749
rect 12529 4709 12541 4743
rect 12575 4740 12587 4743
rect 13538 4740 13544 4752
rect 12575 4712 13544 4740
rect 12575 4709 12587 4712
rect 12529 4703 12587 4709
rect 13538 4700 13544 4712
rect 13596 4700 13602 4752
rect 13722 4740 13728 4752
rect 13683 4712 13728 4740
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 11020 4644 11253 4672
rect 11020 4632 11026 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 11379 4644 12112 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 11112 4576 11437 4604
rect 11112 4564 11118 4576
rect 11425 4573 11437 4576
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 10873 4539 10931 4545
rect 10873 4505 10885 4539
rect 10919 4505 10931 4539
rect 12084 4536 12112 4644
rect 12158 4632 12164 4684
rect 12216 4672 12222 4684
rect 14461 4675 14519 4681
rect 14461 4672 14473 4675
rect 12216 4644 14473 4672
rect 12216 4632 12222 4644
rect 14461 4641 14473 4644
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 12618 4604 12624 4616
rect 12579 4576 12624 4604
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 13044 4576 13829 4604
rect 13044 4564 13050 4576
rect 13817 4573 13829 4576
rect 13863 4573 13875 4607
rect 14734 4604 14740 4616
rect 13817 4567 13875 4573
rect 14476 4576 14740 4604
rect 14476 4536 14504 4576
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 14642 4536 14648 4548
rect 12084 4508 14504 4536
rect 14603 4508 14648 4536
rect 10873 4499 10931 4505
rect 14642 4496 14648 4508
rect 14700 4496 14706 4548
rect 9232 4440 10272 4468
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 12618 4468 12624 4480
rect 11388 4440 12624 4468
rect 11388 4428 11394 4440
rect 12618 4428 12624 4440
rect 12676 4428 12682 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 4062 4264 4068 4276
rect 3292 4236 4068 4264
rect 3292 4224 3298 4236
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 8202 4264 8208 4276
rect 4172 4236 7779 4264
rect 8163 4236 8208 4264
rect 1854 4156 1860 4208
rect 1912 4196 1918 4208
rect 2866 4196 2872 4208
rect 1912 4168 2872 4196
rect 1912 4156 1918 4168
rect 2866 4156 2872 4168
rect 2924 4156 2930 4208
rect 4172 4196 4200 4236
rect 4890 4196 4896 4208
rect 2976 4168 4200 4196
rect 4356 4168 4896 4196
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2314 4128 2320 4140
rect 2188 4100 2320 4128
rect 2188 4088 2194 4100
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2976 4137 3004 4168
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 4246 4128 4252 4140
rect 3191 4100 4252 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4356 4137 4384 4168
rect 4890 4156 4896 4168
rect 4948 4156 4954 4208
rect 6178 4156 6184 4208
rect 6236 4196 6242 4208
rect 6273 4199 6331 4205
rect 6273 4196 6285 4199
rect 6236 4168 6285 4196
rect 6236 4156 6242 4168
rect 6273 4165 6285 4168
rect 6319 4165 6331 4199
rect 7751 4196 7779 4236
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 9674 4264 9680 4276
rect 8680 4236 9680 4264
rect 8680 4196 8708 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 10045 4267 10103 4273
rect 10045 4264 10057 4267
rect 9916 4236 10057 4264
rect 9916 4224 9922 4236
rect 10045 4233 10057 4236
rect 10091 4233 10103 4267
rect 10045 4227 10103 4233
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 10468 4236 10517 4264
rect 10468 4224 10474 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 10505 4227 10563 4233
rect 10686 4224 10692 4276
rect 10744 4264 10750 4276
rect 13170 4264 13176 4276
rect 10744 4236 13176 4264
rect 10744 4224 10750 4236
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 7751 4168 8708 4196
rect 10152 4168 11192 4196
rect 6273 4159 6331 4165
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4488 4100 5028 4128
rect 4488 4088 4494 4100
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 2406 4060 2412 4072
rect 1627 4032 2412 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 4890 4060 4896 4072
rect 4851 4032 4896 4060
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5000 4060 5028 4100
rect 5160 4063 5218 4069
rect 5160 4060 5172 4063
rect 5000 4032 5172 4060
rect 5160 4029 5172 4032
rect 5206 4060 5218 4063
rect 6086 4060 6092 4072
rect 5206 4032 6092 4060
rect 5206 4029 5218 4032
rect 5160 4023 5218 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6288 4060 6316 4159
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 10152 4128 10180 4168
rect 9732 4100 10180 4128
rect 9732 4088 9738 4100
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 11054 4128 11060 4140
rect 10284 4100 11060 4128
rect 10284 4088 10290 4100
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11164 4128 11192 4168
rect 11164 4100 11836 4128
rect 6825 4063 6883 4069
rect 6288 4032 6408 4060
rect 1394 3952 1400 4004
rect 1452 3992 1458 4004
rect 1857 3995 1915 4001
rect 1857 3992 1869 3995
rect 1452 3964 1869 3992
rect 1452 3952 1458 3964
rect 1857 3961 1869 3964
rect 1903 3961 1915 3995
rect 4522 3992 4528 4004
rect 1857 3955 1915 3961
rect 2516 3964 4528 3992
rect 2516 3933 2544 3964
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 6270 3992 6276 4004
rect 5316 3964 6276 3992
rect 5316 3952 5322 3964
rect 6270 3952 6276 3964
rect 6328 3952 6334 4004
rect 6380 3992 6408 4032
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 8202 4060 8208 4072
rect 6871 4032 8208 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7208 4004 7236 4032
rect 8202 4020 8208 4032
rect 8260 4060 8266 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8260 4032 8677 4060
rect 8260 4020 8266 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 11808 4060 11836 4100
rect 12158 4088 12164 4140
rect 12216 4128 12222 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12216 4100 12909 4128
rect 12216 4088 12222 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 14734 4128 14740 4140
rect 13044 4100 13089 4128
rect 14695 4100 14740 4128
rect 13044 4088 13050 4100
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 16758 4128 16764 4140
rect 14976 4100 16764 4128
rect 14976 4088 14982 4100
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 13262 4060 13268 4072
rect 8665 4023 8723 4029
rect 8772 4032 11008 4060
rect 11808 4032 13268 4060
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 6380 3964 7082 3992
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7070 3955 7128 3961
rect 7190 3952 7196 4004
rect 7248 3952 7254 4004
rect 7282 3952 7288 4004
rect 7340 3992 7346 4004
rect 8772 3992 8800 4032
rect 7340 3964 8800 3992
rect 8932 3995 8990 4001
rect 7340 3952 7346 3964
rect 8932 3961 8944 3995
rect 8978 3961 8990 3995
rect 8932 3955 8990 3961
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 2869 3927 2927 3933
rect 2869 3893 2881 3927
rect 2915 3924 2927 3927
rect 3050 3924 3056 3936
rect 2915 3896 3056 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 3694 3924 3700 3936
rect 3655 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 4062 3924 4068 3936
rect 4023 3896 4068 3924
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 7558 3924 7564 3936
rect 4212 3896 7564 3924
rect 4212 3884 4218 3896
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8956 3924 8984 3955
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9490 3992 9496 4004
rect 9088 3964 9496 3992
rect 9088 3952 9094 3964
rect 9490 3952 9496 3964
rect 9548 3992 9554 4004
rect 10873 3995 10931 4001
rect 10873 3992 10885 3995
rect 9548 3964 10885 3992
rect 9548 3952 9554 3964
rect 10873 3961 10885 3964
rect 10919 3961 10931 3995
rect 10980 3992 11008 4032
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 13998 4060 14004 4072
rect 13679 4032 14004 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 13538 3992 13544 4004
rect 10980 3964 13544 3992
rect 10873 3955 10931 3961
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 13906 3992 13912 4004
rect 13867 3964 13912 3992
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 10042 3924 10048 3936
rect 7984 3896 10048 3924
rect 7984 3884 7990 3896
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10965 3927 11023 3933
rect 10965 3924 10977 3927
rect 10192 3896 10977 3924
rect 10192 3884 10198 3896
rect 10965 3893 10977 3896
rect 11011 3893 11023 3927
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 10965 3887 11023 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 12124 3896 12449 3924
rect 12124 3884 12130 3896
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 12802 3924 12808 3936
rect 12763 3896 12808 3924
rect 12437 3887 12495 3893
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 14090 3924 14096 3936
rect 13044 3896 14096 3924
rect 13044 3884 13050 3896
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 2038 3720 2044 3732
rect 1999 3692 2044 3720
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 2832 3692 3157 3720
rect 2832 3680 2838 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3145 3683 3203 3689
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3292 3692 3337 3720
rect 3292 3680 3298 3692
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 3752 3692 4537 3720
rect 3752 3680 3758 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 4525 3683 4583 3689
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 5224 3692 8585 3720
rect 5224 3680 5230 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 9033 3723 9091 3729
rect 9033 3689 9045 3723
rect 9079 3720 9091 3723
rect 9214 3720 9220 3732
rect 9079 3692 9220 3720
rect 9079 3689 9091 3692
rect 9033 3683 9091 3689
rect 9214 3680 9220 3692
rect 9272 3720 9278 3732
rect 9858 3720 9864 3732
rect 9272 3692 9864 3720
rect 9272 3680 9278 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 11238 3720 11244 3732
rect 10008 3692 10548 3720
rect 11199 3692 11244 3720
rect 10008 3680 10014 3692
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 5258 3652 5264 3664
rect 3476 3624 5264 3652
rect 3476 3612 3482 3624
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 6086 3612 6092 3664
rect 6144 3652 6150 3664
rect 6362 3652 6368 3664
rect 6144 3624 6368 3652
rect 6144 3612 6150 3624
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 6822 3612 6828 3664
rect 6880 3652 6886 3664
rect 6880 3624 10272 3652
rect 6880 3612 6886 3624
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 4062 3584 4068 3596
rect 1995 3556 4068 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4614 3584 4620 3596
rect 4575 3556 4620 3584
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4890 3544 4896 3596
rect 4948 3584 4954 3596
rect 5626 3593 5632 3596
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 4948 3556 5365 3584
rect 4948 3544 4954 3556
rect 5353 3553 5365 3556
rect 5399 3553 5411 3587
rect 5620 3584 5632 3593
rect 5539 3556 5632 3584
rect 5353 3547 5411 3553
rect 5620 3547 5632 3556
rect 5684 3584 5690 3596
rect 6730 3584 6736 3596
rect 5684 3556 6736 3584
rect 5626 3544 5632 3547
rect 5684 3544 5690 3556
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7449 3587 7507 3593
rect 7449 3584 7461 3587
rect 6972 3556 7461 3584
rect 6972 3544 6978 3556
rect 7449 3553 7461 3556
rect 7495 3553 7507 3587
rect 7449 3547 7507 3553
rect 9217 3587 9275 3593
rect 9217 3553 9229 3587
rect 9263 3584 9275 3587
rect 9306 3584 9312 3596
rect 9263 3556 9312 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9456 3556 10057 3584
rect 9456 3544 9462 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 2222 3516 2228 3528
rect 2183 3488 2228 3516
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3516 3387 3519
rect 4706 3516 4712 3528
rect 3375 3488 3464 3516
rect 3375 3485 3387 3488
rect 3329 3479 3387 3485
rect 3436 3460 3464 3488
rect 3528 3488 4712 3516
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 2777 3451 2835 3457
rect 2777 3448 2789 3451
rect 2464 3420 2789 3448
rect 2464 3408 2470 3420
rect 2777 3417 2789 3420
rect 2823 3417 2835 3451
rect 2777 3411 2835 3417
rect 3418 3408 3424 3460
rect 3476 3408 3482 3460
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 3528 3380 3556 3488
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 4847 3488 5396 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 4982 3448 4988 3460
rect 4304 3420 4988 3448
rect 4304 3408 4310 3420
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 4154 3380 4160 3392
rect 1627 3352 3556 3380
rect 4115 3352 4160 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 5074 3380 5080 3392
rect 4488 3352 5080 3380
rect 4488 3340 4494 3352
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5368 3380 5396 3488
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6638 3516 6644 3528
rect 6420 3488 6644 3516
rect 6420 3476 6426 3488
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7190 3516 7196 3528
rect 7151 3488 7196 3516
rect 7190 3476 7196 3488
rect 7248 3476 7254 3528
rect 9122 3476 9128 3528
rect 9180 3516 9186 3528
rect 10244 3525 10272 3624
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 9180 3488 10149 3516
rect 9180 3476 9186 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 10520 3516 10548 3692
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 12986 3720 12992 3732
rect 11379 3692 12992 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 14458 3720 14464 3732
rect 13096 3692 14464 3720
rect 10594 3612 10600 3664
rect 10652 3652 10658 3664
rect 12710 3652 12716 3664
rect 10652 3624 12716 3652
rect 10652 3612 10658 3624
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 10778 3544 10784 3596
rect 10836 3584 10842 3596
rect 12437 3587 12495 3593
rect 10836 3556 11560 3584
rect 10836 3544 10842 3556
rect 11330 3516 11336 3528
rect 10520 3488 11336 3516
rect 10229 3479 10287 3485
rect 11330 3476 11336 3488
rect 11388 3516 11394 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 11388 3488 11437 3516
rect 11388 3476 11394 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11532 3516 11560 3556
rect 12437 3553 12449 3587
rect 12483 3584 12495 3587
rect 12802 3584 12808 3596
rect 12483 3556 12808 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 12802 3544 12808 3556
rect 12860 3584 12866 3596
rect 13096 3584 13124 3692
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 13538 3652 13544 3664
rect 13499 3624 13544 3652
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13262 3584 13268 3596
rect 12860 3556 13124 3584
rect 13223 3556 13268 3584
rect 12860 3544 12866 3556
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 14277 3587 14335 3593
rect 14277 3553 14289 3587
rect 14323 3584 14335 3587
rect 14550 3584 14556 3596
rect 14323 3556 14556 3584
rect 14323 3553 14335 3556
rect 14277 3547 14335 3553
rect 14550 3544 14556 3556
rect 14608 3584 14614 3596
rect 14734 3584 14740 3596
rect 14608 3556 14740 3584
rect 14608 3544 14614 3556
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 11532 3488 12541 3516
rect 11425 3479 11483 3485
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 16390 3516 16396 3528
rect 14507 3488 16396 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 9677 3451 9735 3457
rect 9677 3448 9689 3451
rect 8128 3420 9689 3448
rect 5534 3380 5540 3392
rect 5368 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3380 5598 3392
rect 6638 3380 6644 3392
rect 5592 3352 6644 3380
rect 5592 3340 5598 3352
rect 6638 3340 6644 3352
rect 6696 3380 6702 3392
rect 6733 3383 6791 3389
rect 6733 3380 6745 3383
rect 6696 3352 6745 3380
rect 6696 3340 6702 3352
rect 6733 3349 6745 3352
rect 6779 3349 6791 3383
rect 6733 3343 6791 3349
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 8128 3380 8156 3420
rect 9677 3417 9689 3420
rect 9723 3417 9735 3451
rect 9677 3411 9735 3417
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 12636 3448 12664 3479
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 10100 3420 12664 3448
rect 10100 3408 10106 3420
rect 10870 3380 10876 3392
rect 6880 3352 8156 3380
rect 10831 3352 10876 3380
rect 6880 3340 6886 3352
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 12066 3380 12072 3392
rect 12027 3352 12072 3380
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 2501 3179 2559 3185
rect 2501 3176 2513 3179
rect 1820 3148 2513 3176
rect 1820 3136 1826 3148
rect 2501 3145 2513 3148
rect 2547 3145 2559 3179
rect 4430 3176 4436 3188
rect 2501 3139 2559 3145
rect 3620 3148 4436 3176
rect 2222 3068 2228 3120
rect 2280 3108 2286 3120
rect 3620 3108 3648 3148
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 5166 3176 5172 3188
rect 4580 3148 5172 3176
rect 4580 3136 4586 3148
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 6086 3176 6092 3188
rect 5592 3148 6092 3176
rect 5592 3136 5598 3148
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 6512 3148 7779 3176
rect 6512 3136 6518 3148
rect 2280 3080 3648 3108
rect 3697 3111 3755 3117
rect 2280 3068 2286 3080
rect 3697 3077 3709 3111
rect 3743 3108 3755 3111
rect 4890 3108 4896 3120
rect 3743 3080 4896 3108
rect 3743 3077 3755 3080
rect 3697 3071 3755 3077
rect 4890 3068 4896 3080
rect 4948 3068 4954 3120
rect 7751 3108 7779 3148
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8168 3148 8217 3176
rect 8168 3136 8174 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 9398 3176 9404 3188
rect 8711 3148 9404 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10778 3176 10784 3188
rect 10100 3148 10784 3176
rect 10100 3136 10106 3148
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11057 3179 11115 3185
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 12434 3176 12440 3188
rect 11103 3148 12440 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 9861 3111 9919 3117
rect 9861 3108 9873 3111
rect 7751 3080 9873 3108
rect 9861 3077 9873 3080
rect 9907 3077 9919 3111
rect 9861 3071 9919 3077
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 12253 3111 12311 3117
rect 12253 3108 12265 3111
rect 10192 3080 12265 3108
rect 10192 3068 10198 3080
rect 12253 3077 12265 3080
rect 12299 3077 12311 3111
rect 12253 3071 12311 3077
rect 2958 3040 2964 3052
rect 2919 3012 2964 3040
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3970 3040 3976 3052
rect 3191 3012 3976 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4614 3040 4620 3052
rect 4387 3012 4620 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 10226 3000 10232 3052
rect 10284 3040 10290 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10284 3012 10425 3040
rect 10284 3000 10290 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 11606 3040 11612 3052
rect 11567 3012 11612 3040
rect 10413 3003 10471 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 13538 3040 13544 3052
rect 12268 3012 13544 3040
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2972 1639 2975
rect 4430 2972 4436 2984
rect 1627 2944 4436 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 4982 2972 4988 2984
rect 4939 2944 4988 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5160 2975 5218 2981
rect 5160 2941 5172 2975
rect 5206 2972 5218 2975
rect 5442 2972 5448 2984
rect 5206 2944 5448 2972
rect 5206 2941 5218 2944
rect 5160 2935 5218 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 8202 2972 8208 2984
rect 6871 2944 8208 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8996 2944 9137 2972
rect 8996 2932 9002 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2972 10379 2975
rect 12268 2972 12296 3012
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 16022 3040 16028 3052
rect 13679 3012 16028 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 12434 2972 12440 2984
rect 10367 2944 12296 2972
rect 12395 2944 12440 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 12584 2944 13369 2972
rect 12584 2932 12590 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 14277 2975 14335 2981
rect 14277 2941 14289 2975
rect 14323 2972 14335 2975
rect 14366 2972 14372 2984
rect 14323 2944 14372 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 1854 2904 1860 2916
rect 1815 2876 1860 2904
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 2866 2904 2872 2916
rect 2827 2876 2872 2904
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 7092 2907 7150 2913
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 7742 2904 7748 2916
rect 7138 2876 7748 2904
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 9033 2907 9091 2913
rect 9033 2873 9045 2907
rect 9079 2904 9091 2907
rect 11698 2904 11704 2916
rect 9079 2876 11704 2904
rect 9079 2873 9091 2876
rect 9033 2867 9091 2873
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 12253 2907 12311 2913
rect 12253 2873 12265 2907
rect 12299 2904 12311 2907
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 12299 2876 12725 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 12713 2867 12771 2873
rect 14553 2907 14611 2913
rect 14553 2873 14565 2907
rect 14599 2904 14611 2907
rect 15746 2904 15752 2916
rect 14599 2876 15752 2904
rect 14599 2873 14611 2876
rect 14553 2867 14611 2873
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 4065 2839 4123 2845
rect 4065 2805 4077 2839
rect 4111 2836 4123 2839
rect 5626 2836 5632 2848
rect 4111 2808 5632 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 6273 2839 6331 2845
rect 6273 2805 6285 2839
rect 6319 2836 6331 2839
rect 7006 2836 7012 2848
rect 6319 2808 7012 2836
rect 6319 2805 6331 2808
rect 6273 2799 6331 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 10042 2836 10048 2848
rect 7892 2808 10048 2836
rect 7892 2796 7898 2808
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 11146 2836 11152 2848
rect 10275 2808 11152 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 11425 2839 11483 2845
rect 11425 2836 11437 2839
rect 11388 2808 11437 2836
rect 11388 2796 11394 2808
rect 11425 2805 11437 2808
rect 11471 2805 11483 2839
rect 11425 2799 11483 2805
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 11974 2836 11980 2848
rect 11563 2808 11980 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 4430 2632 4436 2644
rect 4391 2604 4436 2632
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 4890 2632 4896 2644
rect 4851 2604 4896 2632
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6917 2635 6975 2641
rect 6917 2632 6929 2635
rect 6135 2604 6929 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6917 2601 6929 2604
rect 6963 2601 6975 2635
rect 6917 2595 6975 2601
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 9122 2632 9128 2644
rect 8159 2604 9128 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 10134 2632 10140 2644
rect 10095 2604 10140 2632
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10410 2632 10416 2644
rect 10275 2604 10416 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 4801 2567 4859 2573
rect 4801 2533 4813 2567
rect 4847 2564 4859 2567
rect 6822 2564 6828 2576
rect 4847 2536 6828 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 6932 2536 8800 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1946 2496 1952 2508
rect 1443 2468 1952 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2400 2499 2458 2505
rect 2400 2465 2412 2499
rect 2446 2496 2458 2499
rect 2866 2496 2872 2508
rect 2446 2468 2872 2496
rect 2446 2465 2458 2468
rect 2400 2459 2458 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5994 2496 6000 2508
rect 5955 2468 6000 2496
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6638 2496 6644 2508
rect 6288 2468 6644 2496
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5718 2428 5724 2440
rect 5123 2400 5724 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 106 2252 112 2304
rect 164 2292 170 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 164 2264 1593 2292
rect 164 2252 170 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 2148 2292 2176 2391
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6288 2437 6316 2468
rect 6638 2456 6644 2468
rect 6696 2496 6702 2508
rect 6932 2496 6960 2536
rect 7282 2496 7288 2508
rect 6696 2468 6960 2496
rect 7243 2468 7288 2496
rect 6696 2456 6702 2468
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2496 7435 2499
rect 7834 2496 7840 2508
rect 7423 2468 7840 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 8662 2496 8668 2508
rect 8527 2468 8668 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8662 2456 8668 2468
rect 8720 2456 8726 2508
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 6788 2400 7481 2428
rect 6788 2388 6794 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 8570 2428 8576 2440
rect 8531 2400 8576 2428
rect 7469 2391 7527 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8772 2437 8800 2536
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 10244 2564 10272 2595
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10502 2592 10508 2644
rect 10560 2632 10566 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10560 2604 10977 2632
rect 10560 2592 10566 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 10965 2595 11023 2601
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 12066 2632 12072 2644
rect 11471 2604 12072 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 14366 2632 14372 2644
rect 12492 2604 14372 2632
rect 12492 2592 12498 2604
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 9456 2536 10272 2564
rect 9456 2524 9462 2536
rect 10778 2524 10784 2576
rect 10836 2564 10842 2576
rect 12158 2564 12164 2576
rect 10836 2536 12164 2564
rect 10836 2524 10842 2536
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 9306 2456 9312 2508
rect 9364 2496 9370 2508
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 9364 2468 9505 2496
rect 9364 2456 9370 2468
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 11330 2496 11336 2508
rect 11291 2468 11336 2496
rect 9493 2459 9551 2465
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 12345 2499 12403 2505
rect 12345 2465 12357 2499
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9214 2428 9220 2440
rect 8803 2400 9220 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10686 2388 10692 2440
rect 10744 2428 10750 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 10744 2400 11529 2428
rect 10744 2388 10750 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 3513 2363 3571 2369
rect 3513 2329 3525 2363
rect 3559 2360 3571 2363
rect 6748 2360 6776 2388
rect 3559 2332 6776 2360
rect 3559 2329 3571 2332
rect 3513 2323 3571 2329
rect 9950 2320 9956 2372
rect 10008 2360 10014 2372
rect 12360 2360 12388 2459
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2496 13967 2499
rect 13998 2496 14004 2508
rect 13955 2468 14004 2496
rect 13955 2465 13967 2468
rect 13909 2459 13967 2465
rect 13998 2456 14004 2468
rect 14056 2456 14062 2508
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12768 2400 12817 2428
rect 12768 2388 12774 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 14185 2431 14243 2437
rect 14185 2397 14197 2431
rect 14231 2428 14243 2431
rect 15378 2428 15384 2440
rect 14231 2400 15384 2428
rect 14231 2397 14243 2400
rect 14185 2391 14243 2397
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 10008 2332 12388 2360
rect 10008 2320 10014 2332
rect 4982 2292 4988 2304
rect 2148 2264 4988 2292
rect 1581 2255 1639 2261
rect 4982 2252 4988 2264
rect 5040 2292 5046 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 5040 2264 9321 2292
rect 5040 2252 5046 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2292 9827 2295
rect 10778 2292 10784 2304
rect 9815 2264 10784 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 12158 2292 12164 2304
rect 12119 2264 12164 2292
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 10318 2088 10324 2100
rect 6052 2060 10324 2088
rect 6052 2048 6058 2060
rect 10318 2048 10324 2060
rect 10376 2088 10382 2100
rect 10870 2088 10876 2100
rect 10376 2060 10876 2088
rect 10376 2048 10382 2060
rect 10870 2048 10876 2060
rect 10928 2048 10934 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 11882 2088 11888 2100
rect 11020 2060 11888 2088
rect 11020 2048 11026 2060
rect 11882 2048 11888 2060
rect 11940 2048 11946 2100
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 7926 2020 7932 2032
rect 3108 1992 7932 2020
rect 3108 1980 3114 1992
rect 7926 1980 7932 1992
rect 7984 1980 7990 2032
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 12158 2020 12164 2032
rect 8260 1992 12164 2020
rect 8260 1980 8266 1992
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 13354 1980 13360 2032
rect 13412 2020 13418 2032
rect 14182 2020 14188 2032
rect 13412 1992 14188 2020
rect 13412 1980 13418 1992
rect 14182 1980 14188 1992
rect 14240 1980 14246 2032
rect 3786 1912 3792 1964
rect 3844 1952 3850 1964
rect 7466 1952 7472 1964
rect 3844 1924 7472 1952
rect 3844 1912 3850 1924
rect 7466 1912 7472 1924
rect 7524 1912 7530 1964
rect 8662 1912 8668 1964
rect 8720 1912 8726 1964
rect 5810 1844 5816 1896
rect 5868 1884 5874 1896
rect 6362 1884 6368 1896
rect 5868 1856 6368 1884
rect 5868 1844 5874 1856
rect 6362 1844 6368 1856
rect 6420 1844 6426 1896
rect 8680 1884 8708 1912
rect 11974 1884 11980 1896
rect 8680 1856 11980 1884
rect 11974 1844 11980 1856
rect 12032 1884 12038 1896
rect 12250 1884 12256 1896
rect 12032 1856 12256 1884
rect 12032 1844 12038 1856
rect 12250 1844 12256 1856
rect 12308 1844 12314 1896
rect 12345 1887 12403 1893
rect 12345 1853 12357 1887
rect 12391 1884 12403 1887
rect 12710 1884 12716 1896
rect 12391 1856 12716 1884
rect 12391 1853 12403 1856
rect 12345 1847 12403 1853
rect 12710 1844 12716 1856
rect 12768 1844 12774 1896
rect 2498 1776 2504 1828
rect 2556 1816 2562 1828
rect 12526 1816 12532 1828
rect 2556 1788 12532 1816
rect 2556 1776 2562 1788
rect 12526 1776 12532 1788
rect 12584 1776 12590 1828
rect 7834 1708 7840 1760
rect 7892 1748 7898 1760
rect 8202 1748 8208 1760
rect 7892 1720 8208 1748
rect 7892 1708 7898 1720
rect 8202 1708 8208 1720
rect 8260 1708 8266 1760
rect 11606 1708 11612 1760
rect 11664 1748 11670 1760
rect 12342 1748 12348 1760
rect 11664 1720 12348 1748
rect 11664 1708 11670 1720
rect 12342 1708 12348 1720
rect 12400 1708 12406 1760
rect 7282 1640 7288 1692
rect 7340 1680 7346 1692
rect 12802 1680 12808 1692
rect 7340 1652 12808 1680
rect 7340 1640 7346 1652
rect 12802 1640 12808 1652
rect 12860 1640 12866 1692
rect 7190 1572 7196 1624
rect 7248 1612 7254 1624
rect 8754 1612 8760 1624
rect 7248 1584 8760 1612
rect 7248 1572 7254 1584
rect 8754 1572 8760 1584
rect 8812 1572 8818 1624
rect 9582 1572 9588 1624
rect 9640 1612 9646 1624
rect 11330 1612 11336 1624
rect 9640 1584 11336 1612
rect 9640 1572 9646 1584
rect 11330 1572 11336 1584
rect 11388 1572 11394 1624
rect 1302 1436 1308 1488
rect 1360 1476 1366 1488
rect 12345 1479 12403 1485
rect 12345 1476 12357 1479
rect 1360 1448 12357 1476
rect 1360 1436 1366 1448
rect 12345 1445 12357 1448
rect 12391 1445 12403 1479
rect 12345 1439 12403 1445
rect 8570 1232 8576 1284
rect 8628 1272 8634 1284
rect 9030 1272 9036 1284
rect 8628 1244 9036 1272
rect 8628 1232 8634 1244
rect 9030 1232 9036 1244
rect 9088 1232 9094 1284
<< via1 >>
rect 4804 18028 4856 18080
rect 9404 18028 9456 18080
rect 5172 17960 5224 18012
rect 9496 17960 9548 18012
rect 7196 17892 7248 17944
rect 12072 17892 12124 17944
rect 3516 17824 3568 17876
rect 9036 17824 9088 17876
rect 6000 17756 6052 17808
rect 11152 17756 11204 17808
rect 4528 17688 4580 17740
rect 10232 17688 10284 17740
rect 6920 17620 6972 17672
rect 11336 17620 11388 17672
rect 4160 17552 4212 17604
rect 9864 17552 9916 17604
rect 10508 17552 10560 17604
rect 12440 17552 12492 17604
rect 5540 17484 5592 17536
rect 10692 17484 10744 17536
rect 11428 17484 11480 17536
rect 16028 17484 16080 17536
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 3056 17280 3108 17332
rect 6184 17280 6236 17332
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 8024 17280 8076 17332
rect 10508 17280 10560 17332
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 2136 17212 2188 17264
rect 2780 17144 2832 17196
rect 3240 17144 3292 17196
rect 6276 17187 6328 17196
rect 6276 17153 6285 17187
rect 6285 17153 6319 17187
rect 6319 17153 6328 17187
rect 6276 17144 6328 17153
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 2964 17119 3016 17128
rect 2964 17085 2973 17119
rect 2973 17085 3007 17119
rect 3007 17085 3016 17119
rect 2964 17076 3016 17085
rect 3976 17076 4028 17128
rect 3884 17008 3936 17060
rect 7104 17076 7156 17128
rect 7196 17076 7248 17128
rect 6000 17051 6052 17060
rect 6000 17017 6009 17051
rect 6009 17017 6043 17051
rect 6043 17017 6052 17051
rect 6000 17008 6052 17017
rect 7380 17051 7432 17060
rect 7380 17017 7389 17051
rect 7389 17017 7423 17051
rect 7423 17017 7432 17051
rect 8392 17144 8444 17196
rect 12808 17144 12860 17196
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 9772 17076 9824 17085
rect 10140 17076 10192 17128
rect 11888 17076 11940 17128
rect 12532 17076 12584 17128
rect 7380 17008 7432 17017
rect 8760 17008 8812 17060
rect 9220 17008 9272 17060
rect 13544 17008 13596 17060
rect 7932 16940 7984 16992
rect 8668 16940 8720 16992
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9680 16940 9732 16992
rect 10508 16940 10560 16992
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 4436 16736 4488 16788
rect 5540 16736 5592 16788
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 9312 16736 9364 16788
rect 11428 16736 11480 16788
rect 12072 16779 12124 16788
rect 12072 16745 12081 16779
rect 12081 16745 12115 16779
rect 12115 16745 12124 16779
rect 12072 16736 12124 16745
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 13544 16779 13596 16788
rect 13544 16745 13553 16779
rect 13553 16745 13587 16779
rect 13587 16745 13596 16779
rect 13544 16736 13596 16745
rect 3332 16668 3384 16720
rect 7840 16668 7892 16720
rect 10048 16668 10100 16720
rect 11244 16668 11296 16720
rect 1952 16600 2004 16652
rect 2136 16600 2188 16652
rect 3976 16600 4028 16652
rect 5356 16600 5408 16652
rect 6644 16600 6696 16652
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 3148 16532 3200 16584
rect 3240 16532 3292 16584
rect 5908 16532 5960 16584
rect 6736 16532 6788 16584
rect 7748 16600 7800 16652
rect 8300 16600 8352 16652
rect 8392 16600 8444 16652
rect 6276 16464 6328 16516
rect 8024 16532 8076 16584
rect 8576 16532 8628 16584
rect 10324 16600 10376 16652
rect 10416 16643 10468 16652
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 11796 16600 11848 16652
rect 12072 16600 12124 16652
rect 12348 16600 12400 16652
rect 12716 16600 12768 16652
rect 9128 16532 9180 16584
rect 10508 16532 10560 16584
rect 7656 16464 7708 16516
rect 9036 16507 9088 16516
rect 9036 16473 9045 16507
rect 9045 16473 9079 16507
rect 9079 16473 9088 16507
rect 9036 16464 9088 16473
rect 9404 16464 9456 16516
rect 9680 16464 9732 16516
rect 5448 16396 5500 16448
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 6736 16396 6788 16448
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 10232 16396 10284 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 3332 16192 3384 16244
rect 6828 16192 6880 16244
rect 4252 16124 4304 16176
rect 4620 16099 4672 16108
rect 4620 16065 4629 16099
rect 4629 16065 4663 16099
rect 4663 16065 4672 16099
rect 4620 16056 4672 16065
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 6920 16056 6972 16108
rect 7840 16056 7892 16108
rect 9956 16192 10008 16244
rect 10784 16124 10836 16176
rect 12624 16167 12676 16176
rect 12624 16133 12633 16167
rect 12633 16133 12667 16167
rect 12667 16133 12676 16167
rect 12624 16124 12676 16133
rect 8852 16056 8904 16108
rect 10876 16056 10928 16108
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 2688 16031 2740 16040
rect 2688 15997 2697 16031
rect 2697 15997 2731 16031
rect 2731 15997 2740 16031
rect 2688 15988 2740 15997
rect 4344 16031 4396 16040
rect 4344 15997 4353 16031
rect 4353 15997 4387 16031
rect 4387 15997 4396 16031
rect 4344 15988 4396 15997
rect 6460 15988 6512 16040
rect 8300 15988 8352 16040
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 9220 15988 9272 16040
rect 9312 15988 9364 16040
rect 9864 15988 9916 16040
rect 10508 15988 10560 16040
rect 11244 15988 11296 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 12900 15988 12952 16040
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 2044 15963 2096 15972
rect 2044 15929 2053 15963
rect 2053 15929 2087 15963
rect 2087 15929 2096 15963
rect 2044 15920 2096 15929
rect 2964 15963 3016 15972
rect 2964 15929 2973 15963
rect 2973 15929 3007 15963
rect 3007 15929 3016 15963
rect 2964 15920 3016 15929
rect 3884 15920 3936 15972
rect 1400 15852 1452 15904
rect 2320 15852 2372 15904
rect 4160 15852 4212 15904
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6368 15852 6420 15904
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 7380 15852 7432 15904
rect 9404 15852 9456 15904
rect 9496 15852 9548 15904
rect 9680 15852 9732 15904
rect 9864 15852 9916 15904
rect 11520 15852 11572 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 1676 15648 1728 15700
rect 5540 15648 5592 15700
rect 7472 15648 7524 15700
rect 8116 15648 8168 15700
rect 5172 15580 5224 15632
rect 8760 15580 8812 15632
rect 9588 15580 9640 15632
rect 13636 15580 13688 15632
rect 5356 15512 5408 15564
rect 5448 15512 5500 15564
rect 5816 15555 5868 15564
rect 5816 15521 5850 15555
rect 5850 15521 5868 15555
rect 5816 15512 5868 15521
rect 8208 15512 8260 15564
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 9496 15555 9548 15564
rect 9496 15521 9505 15555
rect 9505 15521 9539 15555
rect 9539 15521 9548 15555
rect 9496 15512 9548 15521
rect 10692 15512 10744 15564
rect 11428 15512 11480 15564
rect 11704 15512 11756 15564
rect 12164 15512 12216 15564
rect 13084 15555 13136 15564
rect 13084 15521 13093 15555
rect 13093 15521 13127 15555
rect 13127 15521 13136 15555
rect 13084 15512 13136 15521
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 3792 15444 3844 15496
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 7932 15487 7984 15496
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 7932 15444 7984 15453
rect 8300 15444 8352 15496
rect 9956 15444 10008 15496
rect 10508 15444 10560 15496
rect 10968 15444 11020 15496
rect 3240 15376 3292 15428
rect 8944 15376 8996 15428
rect 9128 15376 9180 15428
rect 11152 15444 11204 15496
rect 11336 15444 11388 15496
rect 12072 15376 12124 15428
rect 12256 15376 12308 15428
rect 15384 15376 15436 15428
rect 2780 15308 2832 15360
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 5356 15308 5408 15360
rect 6552 15308 6604 15360
rect 7380 15351 7432 15360
rect 7380 15317 7389 15351
rect 7389 15317 7423 15351
rect 7423 15317 7432 15351
rect 7380 15308 7432 15317
rect 7564 15308 7616 15360
rect 12624 15308 12676 15360
rect 16764 15308 16816 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 2688 15104 2740 15156
rect 3792 15104 3844 15156
rect 3240 15036 3292 15088
rect 3424 15036 3476 15088
rect 2596 14968 2648 15020
rect 3792 14968 3844 15020
rect 4068 14968 4120 15020
rect 8760 15104 8812 15156
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 4804 14968 4856 15020
rect 8576 14968 8628 15020
rect 9128 14968 9180 15020
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 1584 14943 1636 14952
rect 1584 14909 1593 14943
rect 1593 14909 1627 14943
rect 1627 14909 1636 14943
rect 1584 14900 1636 14909
rect 4436 14900 4488 14952
rect 4896 14943 4948 14952
rect 4896 14909 4905 14943
rect 4905 14909 4939 14943
rect 4939 14909 4948 14943
rect 4896 14900 4948 14909
rect 5448 14900 5500 14952
rect 6920 14900 6972 14952
rect 7472 14900 7524 14952
rect 9772 14968 9824 15020
rect 10324 14943 10376 14952
rect 10324 14909 10333 14943
rect 10333 14909 10367 14943
rect 10367 14909 10376 14943
rect 11336 15036 11388 15088
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 10324 14900 10376 14909
rect 11428 14900 11480 14952
rect 11796 14968 11848 15020
rect 12072 14968 12124 15020
rect 12808 15036 12860 15088
rect 13176 14968 13228 15020
rect 14556 14968 14608 15020
rect 12624 14900 12676 14952
rect 12808 14900 12860 14952
rect 1860 14875 1912 14884
rect 1860 14841 1869 14875
rect 1869 14841 1903 14875
rect 1903 14841 1912 14875
rect 1860 14832 1912 14841
rect 3056 14832 3108 14884
rect 4988 14832 5040 14884
rect 8484 14832 8536 14884
rect 4252 14764 4304 14816
rect 4436 14764 4488 14816
rect 5816 14764 5868 14816
rect 8760 14832 8812 14884
rect 9220 14832 9272 14884
rect 11520 14832 11572 14884
rect 9588 14764 9640 14816
rect 10600 14764 10652 14816
rect 14464 14832 14516 14884
rect 12624 14764 12676 14816
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 9128 14603 9180 14612
rect 8576 14492 8628 14544
rect 9128 14569 9137 14603
rect 9137 14569 9171 14603
rect 9171 14569 9180 14603
rect 9128 14560 9180 14569
rect 11796 14560 11848 14612
rect 12716 14560 12768 14612
rect 9772 14492 9824 14544
rect 10140 14535 10192 14544
rect 10140 14501 10149 14535
rect 10149 14501 10183 14535
rect 10183 14501 10192 14535
rect 10140 14492 10192 14501
rect 3056 14424 3108 14476
rect 2872 14356 2924 14408
rect 2504 14288 2556 14340
rect 4436 14424 4488 14476
rect 5264 14424 5316 14476
rect 5448 14467 5500 14476
rect 5448 14433 5457 14467
rect 5457 14433 5491 14467
rect 5491 14433 5500 14467
rect 5448 14424 5500 14433
rect 5540 14424 5592 14476
rect 6000 14424 6052 14476
rect 6828 14424 6880 14476
rect 7840 14424 7892 14476
rect 8024 14424 8076 14476
rect 9220 14424 9272 14476
rect 9588 14424 9640 14476
rect 9680 14424 9732 14476
rect 10508 14424 10560 14476
rect 4528 14356 4580 14408
rect 6920 14356 6972 14408
rect 8300 14356 8352 14408
rect 9772 14356 9824 14408
rect 9864 14356 9916 14408
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 12256 14424 12308 14476
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 12992 14424 13044 14476
rect 14280 14424 14332 14476
rect 14096 14356 14148 14408
rect 4988 14288 5040 14340
rect 5080 14288 5132 14340
rect 5448 14288 5500 14340
rect 2780 14263 2832 14272
rect 2780 14229 2789 14263
rect 2789 14229 2823 14263
rect 2823 14229 2832 14263
rect 2780 14220 2832 14229
rect 6736 14220 6788 14272
rect 8484 14288 8536 14340
rect 10508 14220 10560 14272
rect 10968 14220 11020 14272
rect 12808 14288 12860 14340
rect 12992 14331 13044 14340
rect 12992 14297 13001 14331
rect 13001 14297 13035 14331
rect 13035 14297 13044 14331
rect 12992 14288 13044 14297
rect 13176 14220 13228 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 1584 14016 1636 14068
rect 2596 14016 2648 14068
rect 9312 14016 9364 14068
rect 9588 14016 9640 14068
rect 9772 14016 9824 14068
rect 10416 14016 10468 14068
rect 11060 14016 11112 14068
rect 6828 13948 6880 14000
rect 7840 13948 7892 14000
rect 8300 13948 8352 14000
rect 10600 13948 10652 14000
rect 10968 13948 11020 14000
rect 2504 13923 2556 13932
rect 2504 13889 2513 13923
rect 2513 13889 2547 13923
rect 2547 13889 2556 13923
rect 2504 13880 2556 13889
rect 4896 13923 4948 13932
rect 4896 13889 4905 13923
rect 4905 13889 4939 13923
rect 4939 13889 4948 13923
rect 4896 13880 4948 13889
rect 8116 13880 8168 13932
rect 2044 13812 2096 13864
rect 2780 13744 2832 13796
rect 5724 13812 5776 13864
rect 6736 13812 6788 13864
rect 6920 13812 6972 13864
rect 7472 13812 7524 13864
rect 8300 13812 8352 13864
rect 9864 13812 9916 13864
rect 11520 13880 11572 13932
rect 13820 13880 13872 13932
rect 12716 13812 12768 13864
rect 14188 13812 14240 13864
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 3148 13744 3200 13796
rect 4068 13744 4120 13796
rect 5540 13744 5592 13796
rect 6276 13744 6328 13796
rect 7104 13787 7156 13796
rect 7104 13753 7138 13787
rect 7138 13753 7156 13787
rect 7104 13744 7156 13753
rect 7748 13744 7800 13796
rect 8576 13744 8628 13796
rect 8760 13744 8812 13796
rect 9404 13744 9456 13796
rect 11704 13787 11756 13796
rect 11704 13753 11713 13787
rect 11713 13753 11747 13787
rect 11747 13753 11756 13787
rect 11704 13744 11756 13753
rect 4344 13676 4396 13728
rect 4804 13676 4856 13728
rect 9680 13676 9732 13728
rect 10508 13676 10560 13728
rect 11152 13676 11204 13728
rect 13636 13787 13688 13796
rect 13636 13753 13645 13787
rect 13645 13753 13679 13787
rect 13679 13753 13688 13787
rect 13636 13744 13688 13753
rect 12348 13676 12400 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 2044 13515 2096 13524
rect 2044 13481 2053 13515
rect 2053 13481 2087 13515
rect 2087 13481 2096 13515
rect 2044 13472 2096 13481
rect 3056 13472 3108 13524
rect 7380 13472 7432 13524
rect 4804 13447 4856 13456
rect 4804 13413 4813 13447
rect 4813 13413 4847 13447
rect 4847 13413 4856 13447
rect 4804 13404 4856 13413
rect 7932 13472 7984 13524
rect 8760 13472 8812 13524
rect 9496 13472 9548 13524
rect 9956 13472 10008 13524
rect 4712 13336 4764 13388
rect 5908 13379 5960 13388
rect 5908 13345 5942 13379
rect 5942 13345 5960 13379
rect 7840 13404 7892 13456
rect 8208 13404 8260 13456
rect 11152 13472 11204 13524
rect 12256 13472 12308 13524
rect 13268 13515 13320 13524
rect 13268 13481 13277 13515
rect 13277 13481 13311 13515
rect 13311 13481 13320 13515
rect 13268 13472 13320 13481
rect 13728 13515 13780 13524
rect 13728 13481 13737 13515
rect 13737 13481 13771 13515
rect 13771 13481 13780 13515
rect 14464 13515 14516 13524
rect 13728 13472 13780 13481
rect 11428 13404 11480 13456
rect 13084 13404 13136 13456
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 15292 13404 15344 13456
rect 7472 13379 7524 13388
rect 5908 13336 5960 13345
rect 7472 13345 7481 13379
rect 7481 13345 7515 13379
rect 7515 13345 7524 13379
rect 7472 13336 7524 13345
rect 7564 13336 7616 13388
rect 8852 13336 8904 13388
rect 9404 13336 9456 13388
rect 11704 13336 11756 13388
rect 12256 13336 12308 13388
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 13728 13336 13780 13388
rect 2412 13268 2464 13320
rect 2504 13268 2556 13320
rect 4344 13268 4396 13320
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 5448 13268 5500 13320
rect 10048 13268 10100 13320
rect 11152 13268 11204 13320
rect 12716 13311 12768 13320
rect 4160 13132 4212 13184
rect 4436 13175 4488 13184
rect 4436 13141 4445 13175
rect 4445 13141 4479 13175
rect 4479 13141 4488 13175
rect 4436 13132 4488 13141
rect 8576 13200 8628 13252
rect 5172 13132 5224 13184
rect 7840 13132 7892 13184
rect 9496 13132 9548 13184
rect 9956 13132 10008 13184
rect 10784 13132 10836 13184
rect 11060 13200 11112 13252
rect 12440 13200 12492 13252
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 13820 13311 13872 13320
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 13820 13268 13872 13277
rect 14372 13200 14424 13252
rect 14648 13200 14700 13252
rect 11980 13132 12032 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 2504 12971 2556 12980
rect 2504 12937 2513 12971
rect 2513 12937 2547 12971
rect 2547 12937 2556 12971
rect 2504 12928 2556 12937
rect 4252 12928 4304 12980
rect 4712 12928 4764 12980
rect 10416 12928 10468 12980
rect 10968 12928 11020 12980
rect 12992 12928 13044 12980
rect 13912 12928 13964 12980
rect 4068 12860 4120 12912
rect 4804 12860 4856 12912
rect 4896 12860 4948 12912
rect 6276 12903 6328 12912
rect 6276 12869 6285 12903
rect 6285 12869 6319 12903
rect 6319 12869 6328 12903
rect 6276 12860 6328 12869
rect 8024 12860 8076 12912
rect 10232 12860 10284 12912
rect 12348 12860 12400 12912
rect 2596 12724 2648 12776
rect 8116 12792 8168 12844
rect 10416 12792 10468 12844
rect 10876 12792 10928 12844
rect 11704 12835 11756 12844
rect 1400 12656 1452 12708
rect 2964 12631 3016 12640
rect 2964 12597 2973 12631
rect 2973 12597 3007 12631
rect 3007 12597 3016 12631
rect 2964 12588 3016 12597
rect 4712 12656 4764 12708
rect 5172 12767 5224 12776
rect 5172 12733 5206 12767
rect 5206 12733 5224 12767
rect 5172 12724 5224 12733
rect 5448 12724 5500 12776
rect 6736 12724 6788 12776
rect 6920 12724 6972 12776
rect 7104 12699 7156 12708
rect 7104 12665 7138 12699
rect 7138 12665 7156 12699
rect 7104 12656 7156 12665
rect 7840 12588 7892 12640
rect 8300 12724 8352 12776
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12072 12792 12124 12844
rect 12164 12792 12216 12844
rect 12716 12792 12768 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 11152 12724 11204 12776
rect 9312 12656 9364 12708
rect 9588 12656 9640 12708
rect 11244 12656 11296 12708
rect 13176 12724 13228 12776
rect 13912 12724 13964 12776
rect 14188 12724 14240 12776
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 12164 12656 12216 12708
rect 14832 12699 14884 12708
rect 14832 12665 14841 12699
rect 14841 12665 14875 12699
rect 14875 12665 14884 12699
rect 14832 12656 14884 12665
rect 10232 12588 10284 12640
rect 11520 12588 11572 12640
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 1860 12384 1912 12436
rect 2964 12384 3016 12436
rect 4160 12384 4212 12436
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 3884 12316 3936 12368
rect 4528 12316 4580 12368
rect 4988 12384 5040 12436
rect 5080 12384 5132 12436
rect 6276 12384 6328 12436
rect 7104 12384 7156 12436
rect 8208 12384 8260 12436
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 8852 12384 8904 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 9956 12384 10008 12436
rect 12072 12427 12124 12436
rect 2044 12291 2096 12300
rect 2044 12257 2053 12291
rect 2053 12257 2087 12291
rect 2087 12257 2096 12291
rect 2044 12248 2096 12257
rect 8024 12316 8076 12368
rect 2320 12180 2372 12232
rect 4068 12180 4120 12232
rect 6736 12248 6788 12300
rect 7012 12248 7064 12300
rect 9404 12291 9456 12300
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 6644 12180 6696 12232
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 9680 12248 9732 12300
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 9312 12180 9364 12232
rect 10048 12112 10100 12164
rect 11152 12316 11204 12368
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 12072 12384 12124 12393
rect 12348 12384 12400 12436
rect 13268 12427 13320 12436
rect 13268 12393 13277 12427
rect 13277 12393 13311 12427
rect 13311 12393 13320 12427
rect 13268 12384 13320 12393
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 11980 12248 12032 12300
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 14188 12248 14240 12300
rect 15016 12248 15068 12300
rect 12532 12180 12584 12232
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 12348 12044 12400 12096
rect 13084 12044 13136 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 1860 11883 1912 11892
rect 1860 11849 1869 11883
rect 1869 11849 1903 11883
rect 1903 11849 1912 11883
rect 1860 11840 1912 11849
rect 5540 11840 5592 11892
rect 6368 11840 6420 11892
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 2964 11704 3016 11756
rect 4160 11704 4212 11756
rect 8024 11772 8076 11824
rect 9956 11840 10008 11892
rect 10508 11883 10560 11892
rect 10508 11849 10517 11883
rect 10517 11849 10551 11883
rect 10551 11849 10560 11883
rect 10508 11840 10560 11849
rect 11520 11840 11572 11892
rect 6828 11747 6880 11756
rect 2688 11636 2740 11688
rect 2780 11636 2832 11688
rect 4804 11636 4856 11688
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 6644 11636 6696 11688
rect 11612 11772 11664 11824
rect 9864 11704 9916 11756
rect 9956 11704 10008 11756
rect 10048 11704 10100 11756
rect 12072 11772 12124 11824
rect 13084 11772 13136 11824
rect 14004 11772 14056 11824
rect 14464 11772 14516 11824
rect 12624 11704 12676 11756
rect 13268 11704 13320 11756
rect 15108 11704 15160 11756
rect 3148 11568 3200 11620
rect 2320 11500 2372 11552
rect 3884 11568 3936 11620
rect 4160 11500 4212 11552
rect 4620 11500 4672 11552
rect 4896 11500 4948 11552
rect 6184 11568 6236 11620
rect 7196 11568 7248 11620
rect 9312 11568 9364 11620
rect 9588 11568 9640 11620
rect 10140 11636 10192 11688
rect 9864 11568 9916 11620
rect 11520 11568 11572 11620
rect 5724 11500 5776 11552
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 6644 11500 6696 11552
rect 9496 11500 9548 11552
rect 9772 11500 9824 11552
rect 10324 11500 10376 11552
rect 12440 11636 12492 11688
rect 13452 11636 13504 11688
rect 14740 11636 14792 11688
rect 11704 11568 11756 11620
rect 11888 11568 11940 11620
rect 12164 11568 12216 11620
rect 12992 11568 13044 11620
rect 13084 11568 13136 11620
rect 12716 11500 12768 11552
rect 13544 11500 13596 11552
rect 13912 11500 13964 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 1768 11296 1820 11348
rect 3884 11296 3936 11348
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 4344 11296 4396 11348
rect 4620 11228 4672 11280
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 3976 11160 4028 11212
rect 3148 11092 3200 11144
rect 4344 11092 4396 11144
rect 4896 11228 4948 11280
rect 5724 11228 5776 11280
rect 6736 11296 6788 11348
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 6828 11160 6880 11212
rect 11612 11296 11664 11348
rect 11888 11296 11940 11348
rect 12348 11296 12400 11348
rect 12532 11296 12584 11348
rect 12716 11296 12768 11348
rect 13636 11296 13688 11348
rect 8576 11228 8628 11280
rect 12164 11228 12216 11280
rect 14556 11228 14608 11280
rect 10048 11160 10100 11212
rect 11152 11160 11204 11212
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 5264 11092 5316 11101
rect 8576 11024 8628 11076
rect 10324 11092 10376 11144
rect 12348 11160 12400 11212
rect 12716 11160 12768 11212
rect 14464 11203 14516 11212
rect 14464 11169 14473 11203
rect 14473 11169 14507 11203
rect 14507 11169 14516 11203
rect 14464 11160 14516 11169
rect 12440 11092 12492 11144
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 13544 11092 13596 11144
rect 14188 11092 14240 11144
rect 2136 10956 2188 11008
rect 11980 11024 12032 11076
rect 12348 11024 12400 11076
rect 10232 10956 10284 11008
rect 10876 10999 10928 11008
rect 10876 10965 10885 10999
rect 10885 10965 10919 10999
rect 10919 10965 10928 10999
rect 10876 10956 10928 10965
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 12072 10956 12124 10965
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 1952 10752 2004 10804
rect 9404 10752 9456 10804
rect 10508 10752 10560 10804
rect 11152 10752 11204 10804
rect 4160 10684 4212 10736
rect 5172 10684 5224 10736
rect 7840 10684 7892 10736
rect 8668 10684 8720 10736
rect 12440 10752 12492 10804
rect 2780 10548 2832 10600
rect 4804 10616 4856 10668
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 4344 10548 4396 10600
rect 2320 10523 2372 10532
rect 2320 10489 2329 10523
rect 2329 10489 2363 10523
rect 2363 10489 2372 10523
rect 2320 10480 2372 10489
rect 2964 10480 3016 10532
rect 3424 10480 3476 10532
rect 1584 10412 1636 10464
rect 5264 10480 5316 10532
rect 5448 10480 5500 10532
rect 5632 10480 5684 10532
rect 6460 10412 6512 10464
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 10140 10616 10192 10668
rect 10600 10616 10652 10668
rect 10876 10616 10928 10668
rect 6920 10480 6972 10532
rect 7196 10480 7248 10532
rect 9772 10548 9824 10600
rect 12716 10616 12768 10668
rect 12992 10752 13044 10804
rect 13728 10752 13780 10804
rect 13544 10684 13596 10736
rect 13268 10616 13320 10668
rect 13452 10616 13504 10668
rect 14740 10684 14792 10736
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 9036 10480 9088 10532
rect 9404 10480 9456 10532
rect 10232 10480 10284 10532
rect 8116 10412 8168 10464
rect 9312 10412 9364 10464
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 10508 10412 10560 10421
rect 10600 10412 10652 10464
rect 12624 10480 12676 10532
rect 13728 10548 13780 10600
rect 15292 10548 15344 10600
rect 11336 10412 11388 10464
rect 13452 10412 13504 10464
rect 13544 10412 13596 10464
rect 14188 10412 14240 10464
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2136 10140 2188 10192
rect 3424 10208 3476 10260
rect 7196 10208 7248 10260
rect 8760 10208 8812 10260
rect 9404 10208 9456 10260
rect 10140 10251 10192 10260
rect 4528 10140 4580 10192
rect 6644 10140 6696 10192
rect 9496 10140 9548 10192
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 10416 10208 10468 10260
rect 10692 10208 10744 10260
rect 12072 10208 12124 10260
rect 12440 10251 12492 10260
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 13452 10208 13504 10260
rect 3148 10115 3200 10124
rect 3148 10081 3157 10115
rect 3157 10081 3191 10115
rect 3191 10081 3200 10115
rect 3148 10072 3200 10081
rect 6184 10115 6236 10124
rect 2964 10004 3016 10056
rect 4160 9936 4212 9988
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2780 9868 2832 9877
rect 4804 9868 4856 9920
rect 6184 10081 6218 10115
rect 6218 10081 6236 10115
rect 6184 10072 6236 10081
rect 9772 10072 9824 10124
rect 10232 10072 10284 10124
rect 13268 10140 13320 10192
rect 5724 10004 5776 10056
rect 6920 10004 6972 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10692 10004 10744 10056
rect 11520 10072 11572 10124
rect 14372 10072 14424 10124
rect 11612 10004 11664 10056
rect 12440 10004 12492 10056
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 12808 10004 12860 10056
rect 13728 10004 13780 10056
rect 13636 9936 13688 9988
rect 11060 9868 11112 9920
rect 11980 9868 12032 9920
rect 12992 9868 13044 9920
rect 14372 9868 14424 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 2596 9596 2648 9648
rect 5540 9664 5592 9716
rect 5632 9664 5684 9716
rect 10600 9664 10652 9716
rect 11060 9707 11112 9716
rect 11060 9673 11069 9707
rect 11069 9673 11103 9707
rect 11103 9673 11112 9707
rect 11060 9664 11112 9673
rect 2964 9571 3016 9580
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 3608 9528 3660 9580
rect 4436 9528 4488 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 1400 9392 1452 9444
rect 3516 9392 3568 9444
rect 4068 9392 4120 9444
rect 4252 9392 4304 9444
rect 5172 9435 5224 9444
rect 5172 9401 5206 9435
rect 5206 9401 5224 9435
rect 5172 9392 5224 9401
rect 5448 9460 5500 9512
rect 8576 9596 8628 9648
rect 10692 9596 10744 9648
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 9496 9528 9548 9580
rect 9772 9528 9824 9580
rect 6276 9460 6328 9512
rect 6736 9460 6788 9512
rect 8484 9460 8536 9512
rect 9588 9460 9640 9512
rect 12164 9664 12216 9716
rect 14464 9664 14516 9716
rect 11520 9596 11572 9648
rect 11796 9528 11848 9580
rect 11888 9528 11940 9580
rect 11428 9460 11480 9512
rect 12440 9528 12492 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 13728 9528 13780 9580
rect 7104 9435 7156 9444
rect 7104 9401 7138 9435
rect 7138 9401 7156 9435
rect 14648 9460 14700 9512
rect 7104 9392 7156 9401
rect 2044 9324 2096 9376
rect 3148 9324 3200 9376
rect 4712 9324 4764 9376
rect 6368 9324 6420 9376
rect 7840 9324 7892 9376
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 14188 9392 14240 9444
rect 8208 9324 8260 9333
rect 9312 9324 9364 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 11336 9324 11388 9376
rect 12532 9324 12584 9376
rect 13084 9324 13136 9376
rect 13820 9324 13872 9376
rect 14280 9324 14332 9376
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 1860 9120 1912 9172
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 4344 9120 4396 9172
rect 5172 9120 5224 9172
rect 6460 9120 6512 9172
rect 2780 9052 2832 9104
rect 2596 8984 2648 9036
rect 3608 8984 3660 9036
rect 4896 9052 4948 9104
rect 4160 8984 4212 9036
rect 4620 8984 4672 9036
rect 7104 9052 7156 9104
rect 9220 9120 9272 9172
rect 9680 9120 9732 9172
rect 9956 9120 10008 9172
rect 10692 9120 10744 9172
rect 11888 9120 11940 9172
rect 7840 9052 7892 9104
rect 8208 9052 8260 9104
rect 8668 9052 8720 9104
rect 13912 9052 13964 9104
rect 9956 8984 10008 9036
rect 12164 8984 12216 9036
rect 12348 8984 12400 9036
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 14464 9027 14516 9036
rect 14464 8993 14473 9027
rect 14473 8993 14507 9027
rect 14507 8993 14516 9027
rect 14464 8984 14516 8993
rect 2872 8916 2924 8968
rect 7748 8959 7800 8968
rect 3332 8848 3384 8900
rect 3148 8780 3200 8832
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 8852 8916 8904 8968
rect 3792 8848 3844 8900
rect 4068 8848 4120 8900
rect 6276 8848 6328 8900
rect 5632 8780 5684 8832
rect 9772 8848 9824 8900
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 10048 8848 10100 8900
rect 10416 8916 10468 8968
rect 10600 8916 10652 8968
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 12532 8959 12584 8968
rect 11520 8916 11572 8925
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 12992 8916 13044 8968
rect 13728 8916 13780 8968
rect 10784 8848 10836 8900
rect 12164 8848 12216 8900
rect 12348 8780 12400 8832
rect 13084 8780 13136 8832
rect 13912 8780 13964 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 3148 8576 3200 8628
rect 4620 8576 4672 8628
rect 4712 8576 4764 8628
rect 6276 8619 6328 8628
rect 2596 8508 2648 8560
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 8852 8576 8904 8628
rect 10048 8576 10100 8628
rect 10140 8576 10192 8628
rect 11152 8576 11204 8628
rect 12992 8576 13044 8628
rect 13636 8619 13688 8628
rect 4252 8440 4304 8492
rect 4528 8440 4580 8492
rect 1768 8372 1820 8424
rect 2780 8372 2832 8424
rect 2872 8347 2924 8356
rect 2872 8313 2881 8347
rect 2881 8313 2915 8347
rect 2915 8313 2924 8347
rect 2872 8304 2924 8313
rect 3056 8304 3108 8356
rect 2504 8279 2556 8288
rect 2504 8245 2513 8279
rect 2513 8245 2547 8279
rect 2547 8245 2556 8279
rect 2504 8236 2556 8245
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 3884 8236 3936 8288
rect 6644 8508 6696 8560
rect 8208 8551 8260 8560
rect 8208 8517 8217 8551
rect 8217 8517 8251 8551
rect 8251 8517 8260 8551
rect 8208 8508 8260 8517
rect 9036 8440 9088 8492
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 11060 8440 11112 8492
rect 11796 8508 11848 8560
rect 5632 8372 5684 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 5172 8347 5224 8356
rect 5172 8313 5206 8347
rect 5206 8313 5224 8347
rect 5172 8304 5224 8313
rect 8852 8304 8904 8356
rect 10508 8372 10560 8424
rect 10784 8372 10836 8424
rect 11888 8440 11940 8492
rect 12348 8440 12400 8492
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 13268 8440 13320 8492
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 14464 8508 14516 8560
rect 9588 8304 9640 8356
rect 5540 8236 5592 8288
rect 8668 8236 8720 8288
rect 9772 8304 9824 8356
rect 10324 8347 10376 8356
rect 10324 8313 10333 8347
rect 10333 8313 10367 8347
rect 10367 8313 10376 8347
rect 10324 8304 10376 8313
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 11244 8304 11296 8356
rect 11428 8347 11480 8356
rect 11428 8313 11437 8347
rect 11437 8313 11471 8347
rect 11471 8313 11480 8347
rect 11428 8304 11480 8313
rect 13176 8372 13228 8424
rect 14556 8372 14608 8424
rect 13728 8304 13780 8356
rect 12716 8236 12768 8288
rect 13820 8236 13872 8288
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 2688 8032 2740 8084
rect 2964 8032 3016 8084
rect 2228 7964 2280 8016
rect 9680 8032 9732 8084
rect 10324 8032 10376 8084
rect 10508 8032 10560 8084
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 9772 7964 9824 8016
rect 10692 7964 10744 8016
rect 4436 7896 4488 7948
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2596 7828 2648 7880
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 3792 7828 3844 7880
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 6276 7896 6328 7948
rect 7564 7896 7616 7948
rect 8208 7896 8260 7948
rect 8852 7896 8904 7948
rect 9220 7896 9272 7948
rect 9496 7939 9548 7948
rect 9496 7905 9505 7939
rect 9505 7905 9539 7939
rect 9539 7905 9548 7939
rect 9496 7896 9548 7905
rect 9128 7828 9180 7880
rect 2964 7760 3016 7812
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 4712 7760 4764 7812
rect 4988 7760 5040 7812
rect 5448 7760 5500 7812
rect 5080 7692 5132 7744
rect 5172 7692 5224 7744
rect 6920 7692 6972 7744
rect 8668 7760 8720 7812
rect 10876 7896 10928 7948
rect 11244 7896 11296 7948
rect 12532 8032 12584 8084
rect 12808 8032 12860 8084
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 11520 7964 11572 8016
rect 12164 7896 12216 7948
rect 12624 7964 12676 8016
rect 12900 7896 12952 7948
rect 14740 7896 14792 7948
rect 10692 7828 10744 7880
rect 11612 7828 11664 7880
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 10968 7692 11020 7744
rect 12808 7760 12860 7812
rect 13268 7828 13320 7880
rect 14188 7828 14240 7880
rect 14464 7760 14516 7812
rect 13176 7692 13228 7744
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 2872 7488 2924 7540
rect 3240 7488 3292 7540
rect 9036 7488 9088 7540
rect 10876 7488 10928 7540
rect 11336 7488 11388 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 14004 7488 14056 7540
rect 14832 7488 14884 7540
rect 2320 7420 2372 7472
rect 2964 7420 3016 7472
rect 4620 7420 4672 7472
rect 8208 7463 8260 7472
rect 8208 7429 8217 7463
rect 8217 7429 8251 7463
rect 8251 7429 8260 7463
rect 8208 7420 8260 7429
rect 6828 7395 6880 7404
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 2964 7284 3016 7336
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 7840 7352 7892 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 12716 7420 12768 7472
rect 3792 7284 3844 7336
rect 4804 7284 4856 7336
rect 3332 7259 3384 7268
rect 3332 7225 3366 7259
rect 3366 7225 3384 7259
rect 3332 7216 3384 7225
rect 5172 7259 5224 7268
rect 5172 7225 5206 7259
rect 5206 7225 5224 7259
rect 5172 7216 5224 7225
rect 7012 7216 7064 7268
rect 3516 7148 3568 7200
rect 3792 7148 3844 7200
rect 4528 7148 4580 7200
rect 5448 7148 5500 7200
rect 6920 7148 6972 7200
rect 8116 7148 8168 7200
rect 8760 7284 8812 7336
rect 9680 7284 9732 7336
rect 10600 7352 10652 7404
rect 10784 7352 10836 7404
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 12900 7352 12952 7404
rect 13268 7420 13320 7472
rect 13176 7352 13228 7404
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 12440 7284 12492 7336
rect 15016 7284 15068 7336
rect 9864 7148 9916 7200
rect 10140 7148 10192 7200
rect 10232 7148 10284 7200
rect 11152 7216 11204 7268
rect 12348 7216 12400 7268
rect 12716 7216 12768 7268
rect 13176 7216 13228 7268
rect 13544 7216 13596 7268
rect 11704 7148 11756 7200
rect 12992 7148 13044 7200
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 14188 7148 14240 7200
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 2044 6944 2096 6996
rect 2412 6876 2464 6928
rect 2688 6876 2740 6928
rect 3240 6876 3292 6928
rect 5540 6876 5592 6928
rect 6092 6919 6144 6928
rect 6092 6885 6126 6919
rect 6126 6885 6144 6919
rect 6092 6876 6144 6885
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2780 6808 2832 6860
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 7564 6808 7616 6860
rect 7748 6808 7800 6860
rect 8116 6944 8168 6996
rect 10232 6944 10284 6996
rect 10508 6944 10560 6996
rect 12532 6944 12584 6996
rect 12808 6944 12860 6996
rect 14004 6944 14056 6996
rect 8208 6876 8260 6928
rect 8668 6876 8720 6928
rect 10140 6876 10192 6928
rect 10784 6876 10836 6928
rect 11704 6876 11756 6928
rect 12164 6876 12216 6928
rect 13084 6919 13136 6928
rect 13084 6885 13093 6919
rect 13093 6885 13127 6919
rect 13127 6885 13136 6919
rect 13084 6876 13136 6885
rect 3516 6740 3568 6792
rect 5080 6783 5132 6792
rect 2044 6604 2096 6656
rect 4436 6672 4488 6724
rect 3056 6604 3108 6656
rect 3148 6604 3200 6656
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5540 6740 5592 6792
rect 4804 6672 4856 6724
rect 5632 6672 5684 6724
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 9404 6740 9456 6792
rect 11612 6740 11664 6792
rect 12440 6808 12492 6860
rect 12624 6808 12676 6860
rect 12992 6740 13044 6792
rect 14004 6808 14056 6860
rect 13268 6672 13320 6724
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 13728 6672 13780 6724
rect 11336 6604 11388 6656
rect 12900 6604 12952 6656
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 1860 6443 1912 6452
rect 1860 6409 1869 6443
rect 1869 6409 1903 6443
rect 1903 6409 1912 6443
rect 1860 6400 1912 6409
rect 2228 6400 2280 6452
rect 5172 6400 5224 6452
rect 7196 6400 7248 6452
rect 4252 6332 4304 6384
rect 8208 6400 8260 6452
rect 10048 6443 10100 6452
rect 2228 6264 2280 6316
rect 8484 6332 8536 6384
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 10968 6400 11020 6452
rect 2964 6196 3016 6248
rect 2136 6060 2188 6112
rect 3792 6196 3844 6248
rect 4804 6196 4856 6248
rect 10416 6332 10468 6384
rect 11704 6264 11756 6316
rect 12532 6400 12584 6452
rect 13728 6332 13780 6384
rect 13360 6264 13412 6316
rect 14464 6264 14516 6316
rect 15016 6264 15068 6316
rect 6828 6239 6880 6248
rect 3332 6171 3384 6180
rect 3332 6137 3366 6171
rect 3366 6137 3384 6171
rect 3332 6128 3384 6137
rect 3976 6128 4028 6180
rect 5172 6171 5224 6180
rect 4804 6060 4856 6112
rect 5172 6137 5206 6171
rect 5206 6137 5224 6171
rect 5172 6128 5224 6137
rect 6092 6128 6144 6180
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 8576 6196 8628 6248
rect 8760 6196 8812 6248
rect 10324 6196 10376 6248
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 13728 6196 13780 6248
rect 7104 6171 7156 6180
rect 7104 6137 7138 6171
rect 7138 6137 7156 6171
rect 7104 6128 7156 6137
rect 7748 6060 7800 6112
rect 8668 6060 8720 6112
rect 10784 6128 10836 6180
rect 9864 6060 9916 6112
rect 11244 6060 11296 6112
rect 12624 6128 12676 6180
rect 12900 6171 12952 6180
rect 12900 6137 12909 6171
rect 12909 6137 12943 6171
rect 12943 6137 12952 6171
rect 12900 6128 12952 6137
rect 13268 6128 13320 6180
rect 12992 6060 13044 6112
rect 13176 6060 13228 6112
rect 13452 6060 13504 6112
rect 13820 6060 13872 6112
rect 15016 6103 15068 6112
rect 15016 6069 15025 6103
rect 15025 6069 15059 6103
rect 15059 6069 15068 6103
rect 15016 6060 15068 6069
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 2044 5899 2096 5908
rect 2044 5865 2053 5899
rect 2053 5865 2087 5899
rect 2087 5865 2096 5899
rect 2044 5856 2096 5865
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3424 5856 3476 5908
rect 5172 5856 5224 5908
rect 10232 5856 10284 5908
rect 12348 5899 12400 5908
rect 11336 5788 11388 5840
rect 12348 5865 12357 5899
rect 12357 5865 12391 5899
rect 12391 5865 12400 5899
rect 12348 5856 12400 5865
rect 12808 5856 12860 5908
rect 13728 5856 13780 5908
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 3240 5695 3292 5704
rect 1952 5584 2004 5636
rect 2136 5584 2188 5636
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 4436 5584 4488 5636
rect 2964 5516 3016 5568
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 4804 5720 4856 5772
rect 6276 5720 6328 5772
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 7380 5763 7432 5772
rect 5172 5652 5224 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 6644 5652 6696 5704
rect 7380 5729 7403 5763
rect 7403 5729 7432 5763
rect 7380 5720 7432 5729
rect 7656 5720 7708 5772
rect 8208 5720 8260 5772
rect 9496 5720 9548 5772
rect 8116 5652 8168 5704
rect 12164 5720 12216 5772
rect 9956 5652 10008 5704
rect 10968 5652 11020 5704
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 12900 5788 12952 5840
rect 12532 5720 12584 5772
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 12992 5720 13044 5772
rect 13360 5652 13412 5704
rect 6920 5516 6972 5568
rect 8208 5584 8260 5636
rect 10876 5584 10928 5636
rect 11704 5584 11756 5636
rect 10416 5516 10468 5568
rect 11244 5516 11296 5568
rect 12348 5516 12400 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 3332 5312 3384 5364
rect 4436 5355 4488 5364
rect 4436 5321 4445 5355
rect 4445 5321 4479 5355
rect 4479 5321 4488 5355
rect 4436 5312 4488 5321
rect 2596 5244 2648 5296
rect 8024 5244 8076 5296
rect 9772 5312 9824 5364
rect 8392 5244 8444 5296
rect 9680 5244 9732 5296
rect 10140 5312 10192 5364
rect 10876 5312 10928 5364
rect 12348 5312 12400 5364
rect 13176 5312 13228 5364
rect 9956 5244 10008 5296
rect 2780 5108 2832 5160
rect 3608 5108 3660 5160
rect 4804 5108 4856 5160
rect 3792 5040 3844 5092
rect 4436 5040 4488 5092
rect 6460 5108 6512 5160
rect 5172 5083 5224 5092
rect 5172 5049 5206 5083
rect 5206 5049 5224 5083
rect 5172 5040 5224 5049
rect 5540 5040 5592 5092
rect 6644 5040 6696 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 5724 4972 5776 5024
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 8392 5108 8444 5160
rect 6920 5040 6972 5092
rect 10140 5176 10192 5228
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 7196 4972 7248 5024
rect 7748 4972 7800 5024
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 12624 5244 12676 5296
rect 13820 5244 13872 5296
rect 11428 5176 11480 5228
rect 10968 5108 11020 5117
rect 11612 5108 11664 5160
rect 10232 5040 10284 5092
rect 11336 5040 11388 5092
rect 12440 5040 12492 5092
rect 12992 5040 13044 5092
rect 13176 5176 13228 5228
rect 14096 5108 14148 5160
rect 13544 5040 13596 5092
rect 14556 5040 14608 5092
rect 10508 5015 10560 5024
rect 10508 4981 10517 5015
rect 10517 4981 10551 5015
rect 10551 4981 10560 5015
rect 10508 4972 10560 4981
rect 11152 4972 11204 5024
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 6644 4768 6696 4820
rect 6920 4768 6972 4820
rect 9680 4768 9732 4820
rect 11428 4768 11480 4820
rect 12808 4768 12860 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14188 4768 14240 4820
rect 2044 4632 2096 4684
rect 3056 4632 3108 4684
rect 4620 4675 4672 4684
rect 4620 4641 4629 4675
rect 4629 4641 4663 4675
rect 4663 4641 4672 4675
rect 4620 4632 4672 4641
rect 3240 4496 3292 4548
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 3700 4564 3752 4616
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 5264 4632 5316 4684
rect 5540 4632 5592 4684
rect 8300 4632 8352 4684
rect 9312 4675 9364 4684
rect 4896 4564 4948 4573
rect 2780 4428 2832 4437
rect 4160 4428 4212 4480
rect 4620 4428 4672 4480
rect 7196 4564 7248 4616
rect 5264 4496 5316 4548
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 9772 4632 9824 4684
rect 10692 4632 10744 4684
rect 8760 4564 8812 4616
rect 9588 4564 9640 4616
rect 5632 4428 5684 4480
rect 6092 4428 6144 4480
rect 6828 4471 6880 4480
rect 6828 4437 6837 4471
rect 6837 4437 6871 4471
rect 6871 4437 6880 4471
rect 6828 4428 6880 4437
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 9680 4539 9732 4548
rect 9680 4505 9689 4539
rect 9689 4505 9723 4539
rect 9723 4505 9732 4539
rect 9680 4496 9732 4505
rect 12348 4700 12400 4752
rect 13544 4700 13596 4752
rect 13728 4743 13780 4752
rect 13728 4709 13737 4743
rect 13737 4709 13771 4743
rect 13771 4709 13780 4743
rect 13728 4700 13780 4709
rect 10968 4632 11020 4684
rect 11060 4564 11112 4616
rect 12164 4632 12216 4684
rect 12624 4607 12676 4616
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 12992 4564 13044 4616
rect 14740 4564 14792 4616
rect 14648 4539 14700 4548
rect 14648 4505 14657 4539
rect 14657 4505 14691 4539
rect 14691 4505 14700 4539
rect 14648 4496 14700 4505
rect 11336 4428 11388 4480
rect 12624 4428 12676 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 3240 4224 3292 4276
rect 4068 4224 4120 4276
rect 8208 4267 8260 4276
rect 1860 4156 1912 4208
rect 2872 4156 2924 4208
rect 2136 4088 2188 4140
rect 2320 4088 2372 4140
rect 4252 4088 4304 4140
rect 4896 4156 4948 4208
rect 6184 4156 6236 4208
rect 8208 4233 8217 4267
rect 8217 4233 8251 4267
rect 8251 4233 8260 4267
rect 8208 4224 8260 4233
rect 9680 4224 9732 4276
rect 9864 4224 9916 4276
rect 10416 4224 10468 4276
rect 10692 4224 10744 4276
rect 13176 4224 13228 4276
rect 4436 4088 4488 4140
rect 2412 4020 2464 4072
rect 4896 4063 4948 4072
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 4896 4020 4948 4029
rect 6092 4020 6144 4072
rect 9680 4088 9732 4140
rect 10232 4088 10284 4140
rect 11060 4131 11112 4140
rect 11060 4097 11069 4131
rect 11069 4097 11103 4131
rect 11103 4097 11112 4131
rect 11060 4088 11112 4097
rect 1400 3952 1452 4004
rect 4528 3952 4580 4004
rect 5264 3952 5316 4004
rect 6276 3952 6328 4004
rect 8208 4020 8260 4072
rect 12164 4088 12216 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 14740 4131 14792 4140
rect 12992 4088 13044 4097
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 14924 4088 14976 4140
rect 16764 4088 16816 4140
rect 7196 3952 7248 4004
rect 7288 3952 7340 4004
rect 3056 3884 3108 3936
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 7564 3884 7616 3936
rect 7932 3884 7984 3936
rect 9036 3952 9088 4004
rect 9496 3952 9548 4004
rect 13268 4020 13320 4072
rect 14004 4020 14056 4072
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 13544 3952 13596 4004
rect 13912 3995 13964 4004
rect 13912 3961 13921 3995
rect 13921 3961 13955 3995
rect 13955 3961 13964 3995
rect 13912 3952 13964 3961
rect 10048 3884 10100 3936
rect 10140 3884 10192 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12072 3884 12124 3936
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 12992 3884 13044 3936
rect 14096 3884 14148 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 2044 3723 2096 3732
rect 2044 3689 2053 3723
rect 2053 3689 2087 3723
rect 2087 3689 2096 3723
rect 2044 3680 2096 3689
rect 2780 3680 2832 3732
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 3700 3680 3752 3732
rect 5172 3680 5224 3732
rect 9220 3680 9272 3732
rect 9864 3680 9916 3732
rect 9956 3680 10008 3732
rect 11244 3723 11296 3732
rect 3424 3612 3476 3664
rect 5264 3612 5316 3664
rect 6092 3612 6144 3664
rect 6368 3612 6420 3664
rect 6828 3612 6880 3664
rect 4068 3544 4120 3596
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 4896 3544 4948 3596
rect 5632 3587 5684 3596
rect 5632 3553 5666 3587
rect 5666 3553 5684 3587
rect 5632 3544 5684 3553
rect 6736 3544 6788 3596
rect 6920 3544 6972 3596
rect 9312 3544 9364 3596
rect 9404 3544 9456 3596
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 2412 3408 2464 3460
rect 3424 3408 3476 3460
rect 4712 3476 4764 3528
rect 4252 3408 4304 3460
rect 4988 3408 5040 3460
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 4436 3340 4488 3392
rect 5080 3340 5132 3392
rect 6368 3476 6420 3528
rect 6644 3476 6696 3528
rect 7196 3519 7248 3528
rect 7196 3485 7205 3519
rect 7205 3485 7239 3519
rect 7239 3485 7248 3519
rect 7196 3476 7248 3485
rect 9128 3476 9180 3528
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 12992 3680 13044 3732
rect 10600 3612 10652 3664
rect 12716 3612 12768 3664
rect 10784 3544 10836 3596
rect 11336 3476 11388 3528
rect 12808 3544 12860 3596
rect 14464 3680 14516 3732
rect 13544 3655 13596 3664
rect 13544 3621 13553 3655
rect 13553 3621 13587 3655
rect 13587 3621 13596 3655
rect 13544 3612 13596 3621
rect 13268 3587 13320 3596
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 14556 3544 14608 3596
rect 14740 3544 14792 3596
rect 5540 3340 5592 3392
rect 6644 3340 6696 3392
rect 6828 3340 6880 3392
rect 10048 3408 10100 3460
rect 16396 3476 16448 3528
rect 10876 3383 10928 3392
rect 10876 3349 10885 3383
rect 10885 3349 10919 3383
rect 10919 3349 10928 3383
rect 10876 3340 10928 3349
rect 12072 3383 12124 3392
rect 12072 3349 12081 3383
rect 12081 3349 12115 3383
rect 12115 3349 12124 3383
rect 12072 3340 12124 3349
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 1768 3136 1820 3188
rect 2228 3068 2280 3120
rect 4436 3136 4488 3188
rect 4528 3136 4580 3188
rect 5172 3136 5224 3188
rect 5540 3136 5592 3188
rect 6092 3136 6144 3188
rect 6460 3136 6512 3188
rect 4896 3068 4948 3120
rect 8116 3136 8168 3188
rect 9404 3136 9456 3188
rect 10048 3136 10100 3188
rect 10784 3136 10836 3188
rect 12440 3136 12492 3188
rect 10140 3068 10192 3120
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 3976 3000 4028 3052
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4620 3000 4672 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 10232 3000 10284 3052
rect 11612 3043 11664 3052
rect 11612 3009 11621 3043
rect 11621 3009 11655 3043
rect 11655 3009 11664 3043
rect 11612 3000 11664 3009
rect 4436 2932 4488 2984
rect 4988 2932 5040 2984
rect 5448 2932 5500 2984
rect 8208 2932 8260 2984
rect 8944 2932 8996 2984
rect 13544 3000 13596 3052
rect 16028 3000 16080 3052
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 12532 2932 12584 2984
rect 14372 2932 14424 2984
rect 1860 2907 1912 2916
rect 1860 2873 1869 2907
rect 1869 2873 1903 2907
rect 1903 2873 1912 2907
rect 1860 2864 1912 2873
rect 2872 2907 2924 2916
rect 2872 2873 2881 2907
rect 2881 2873 2915 2907
rect 2915 2873 2924 2907
rect 2872 2864 2924 2873
rect 7748 2864 7800 2916
rect 11704 2864 11756 2916
rect 15752 2864 15804 2916
rect 5632 2796 5684 2848
rect 7012 2796 7064 2848
rect 7840 2796 7892 2848
rect 10048 2796 10100 2848
rect 11152 2796 11204 2848
rect 11336 2796 11388 2848
rect 11980 2796 12032 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 4896 2635 4948 2644
rect 4896 2601 4905 2635
rect 4905 2601 4939 2635
rect 4939 2601 4948 2635
rect 4896 2592 4948 2601
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 9128 2592 9180 2644
rect 10140 2635 10192 2644
rect 10140 2601 10149 2635
rect 10149 2601 10183 2635
rect 10183 2601 10192 2635
rect 10140 2592 10192 2601
rect 6828 2524 6880 2576
rect 1952 2456 2004 2508
rect 2872 2456 2924 2508
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 112 2252 164 2304
rect 5724 2388 5776 2440
rect 6644 2456 6696 2508
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 7840 2456 7892 2508
rect 8668 2456 8720 2508
rect 6736 2388 6788 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9404 2524 9456 2576
rect 10416 2592 10468 2644
rect 10508 2592 10560 2644
rect 12072 2592 12124 2644
rect 12440 2592 12492 2644
rect 14372 2592 14424 2644
rect 10784 2524 10836 2576
rect 12164 2524 12216 2576
rect 9312 2456 9364 2508
rect 11336 2499 11388 2508
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 9220 2388 9272 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10692 2388 10744 2440
rect 9956 2320 10008 2372
rect 12532 2456 12584 2508
rect 14004 2456 14056 2508
rect 12716 2388 12768 2440
rect 15384 2388 15436 2440
rect 4988 2252 5040 2304
rect 10784 2252 10836 2304
rect 12164 2295 12216 2304
rect 12164 2261 12173 2295
rect 12173 2261 12207 2295
rect 12207 2261 12216 2295
rect 12164 2252 12216 2261
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 6000 2048 6052 2100
rect 10324 2048 10376 2100
rect 10876 2048 10928 2100
rect 10968 2048 11020 2100
rect 11888 2048 11940 2100
rect 3056 1980 3108 2032
rect 7932 1980 7984 2032
rect 8208 1980 8260 2032
rect 12164 1980 12216 2032
rect 13360 1980 13412 2032
rect 14188 1980 14240 2032
rect 3792 1912 3844 1964
rect 7472 1912 7524 1964
rect 8668 1912 8720 1964
rect 5816 1844 5868 1896
rect 6368 1844 6420 1896
rect 11980 1844 12032 1896
rect 12256 1844 12308 1896
rect 12716 1844 12768 1896
rect 2504 1776 2556 1828
rect 12532 1776 12584 1828
rect 7840 1708 7892 1760
rect 8208 1708 8260 1760
rect 11612 1708 11664 1760
rect 12348 1708 12400 1760
rect 7288 1640 7340 1692
rect 12808 1640 12860 1692
rect 7196 1572 7248 1624
rect 8760 1572 8812 1624
rect 9588 1572 9640 1624
rect 11336 1572 11388 1624
rect 1308 1436 1360 1488
rect 8576 1232 8628 1284
rect 9036 1232 9088 1284
<< metal2 >>
rect 110 19200 166 20000
rect 386 19200 442 20000
rect 754 19200 810 20000
rect 1122 19200 1178 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2410 19200 2466 20000
rect 2778 19200 2834 20000
rect 2962 19408 3018 19417
rect 2962 19343 3018 19352
rect 1412 15910 1440 19200
rect 1780 16130 1808 19200
rect 2148 17270 2176 19200
rect 2136 17264 2188 17270
rect 2136 17206 2188 17212
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1504 16102 1808 16130
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1400 12708 1452 12714
rect 1400 12650 1452 12656
rect 1412 11393 1440 12650
rect 1398 11384 1454 11393
rect 1398 11319 1454 11328
rect 1400 9444 1452 9450
rect 1400 9386 1452 9392
rect 1306 6488 1362 6497
rect 1306 6423 1362 6432
rect 1122 6216 1178 6225
rect 1122 6151 1178 6160
rect 754 5128 810 5137
rect 754 5063 810 5072
rect 386 4720 442 4729
rect 386 4655 442 4664
rect 112 2304 164 2310
rect 112 2246 164 2252
rect 124 800 152 2246
rect 400 800 428 4655
rect 768 800 796 5063
rect 1136 800 1164 6151
rect 1320 1494 1348 6423
rect 1412 4457 1440 9386
rect 1398 4448 1454 4457
rect 1398 4383 1454 4392
rect 1400 4004 1452 4010
rect 1400 3946 1452 3952
rect 1412 2417 1440 3946
rect 1504 2825 1532 16102
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1596 14074 1624 14894
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10266 1624 10406
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 5914 1624 9454
rect 1688 7449 1716 15642
rect 1780 11354 1808 15982
rect 1860 14884 1912 14890
rect 1860 14826 1912 14832
rect 1872 14385 1900 14826
rect 1858 14376 1914 14385
rect 1858 14311 1914 14320
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1872 11898 1900 12378
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1964 11370 1992 16594
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 2056 13870 2084 15914
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2042 13560 2098 13569
rect 2042 13495 2044 13504
rect 2096 13495 2098 13504
rect 2044 13466 2096 13472
rect 2042 12336 2098 12345
rect 2042 12271 2044 12280
rect 2096 12271 2098 12280
rect 2044 12242 2096 12248
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1872 11342 1992 11370
rect 1872 10441 1900 11342
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1964 10810 1992 11154
rect 2148 11098 2176 16594
rect 2424 15994 2452 19200
rect 2792 18601 2820 19200
rect 2778 18592 2834 18601
rect 2778 18527 2834 18536
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 17202 2820 18391
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2976 17134 3004 19343
rect 3146 19200 3202 20000
rect 3514 19200 3570 20000
rect 3790 19200 3846 20000
rect 4158 19200 4214 20000
rect 4526 19200 4582 20000
rect 4802 19200 4858 20000
rect 5170 19200 5226 20000
rect 5538 19200 5594 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7194 19200 7250 20000
rect 7562 19200 7618 20000
rect 7930 19200 7986 20000
rect 8206 19200 8262 20000
rect 8574 19200 8630 20000
rect 8942 19200 8998 20000
rect 9218 19200 9274 20000
rect 9586 19200 9642 20000
rect 9954 19200 10010 20000
rect 10322 19200 10378 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11610 19200 11666 20000
rect 11978 19200 12034 20000
rect 12346 19200 12402 20000
rect 12622 19200 12678 20000
rect 12990 19200 13046 20000
rect 13358 19200 13414 20000
rect 13726 19200 13782 20000
rect 14002 19200 14058 20000
rect 14370 19200 14426 20000
rect 14738 19200 14794 20000
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15750 19200 15806 20000
rect 16026 19200 16082 20000
rect 16394 19200 16450 20000
rect 16762 19200 16818 20000
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2056 11070 2176 11098
rect 2240 15966 2452 15994
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1858 10432 1914 10441
rect 1858 10367 1914 10376
rect 2056 9466 2084 11070
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2148 10198 2176 10950
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 1872 9438 2084 9466
rect 1872 9178 1900 9438
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9178 2084 9318
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1674 7440 1730 7449
rect 1674 7375 1730 7384
rect 1674 6352 1730 6361
rect 1674 6287 1730 6296
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1490 2816 1546 2825
rect 1490 2751 1546 2760
rect 1398 2408 1454 2417
rect 1398 2343 1454 2352
rect 1308 1488 1360 1494
rect 1308 1430 1360 1436
rect 1596 1306 1624 5607
rect 1688 3074 1716 6287
rect 1780 3194 1808 8366
rect 2240 8242 2268 15966
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 12628 2360 15846
rect 2700 15162 2728 15982
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2872 15496 2924 15502
rect 2976 15473 3004 15914
rect 2872 15438 2924 15444
rect 2962 15464 3018 15473
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2410 14376 2466 14385
rect 2410 14311 2466 14320
rect 2504 14340 2556 14346
rect 2424 13326 2452 14311
rect 2504 14282 2556 14288
rect 2516 13938 2544 14282
rect 2608 14074 2636 14962
rect 2792 14362 2820 15302
rect 2884 14498 2912 15438
rect 2962 15399 3018 15408
rect 3068 14890 3096 17274
rect 3160 17218 3188 19200
rect 3528 17882 3556 19200
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3804 17762 3832 19200
rect 4172 17864 4200 19200
rect 4172 17836 4292 17864
rect 3804 17734 4200 17762
rect 4172 17610 4200 17734
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3160 17202 3280 17218
rect 3160 17196 3292 17202
rect 3160 17190 3240 17196
rect 3240 17138 3292 17144
rect 3976 17128 4028 17134
rect 3882 17096 3938 17105
rect 4028 17076 4108 17082
rect 3976 17070 4108 17076
rect 3988 17054 4108 17070
rect 3882 17031 3884 17040
rect 3936 17031 3938 17040
rect 3884 17002 3936 17008
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 2884 14470 3004 14498
rect 2700 14334 2820 14362
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2700 13682 2728 14334
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13802 2820 14214
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2700 13654 2820 13682
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12986 2544 13262
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2686 12744 2742 12753
rect 2332 12600 2452 12628
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2332 11558 2360 12174
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2318 10568 2374 10577
rect 2318 10503 2320 10512
rect 2372 10503 2374 10512
rect 2320 10474 2372 10480
rect 2148 8214 2268 8242
rect 1950 7984 2006 7993
rect 1950 7919 2006 7928
rect 1858 7032 1914 7041
rect 1964 7002 1992 7919
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7002 2084 7822
rect 1858 6967 1914 6976
rect 1952 6996 2004 7002
rect 1872 6458 1900 6967
rect 1952 6938 2004 6944
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2148 6882 2176 8214
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2240 7342 2268 7958
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 1964 6854 2176 6882
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1964 5642 1992 6854
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 5914 2084 6598
rect 2240 6458 2268 6734
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2148 5794 2176 6054
rect 2056 5766 2176 5794
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 2056 5522 2084 5766
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 1964 5494 2084 5522
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1872 4214 1900 4966
rect 1964 4865 1992 5494
rect 1950 4856 2006 4865
rect 1950 4791 2006 4800
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1688 3046 1808 3074
rect 1412 1278 1624 1306
rect 1412 800 1440 1278
rect 1780 800 1808 3046
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1872 1465 1900 2858
rect 1964 2514 1992 4791
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 2056 3777 2084 4626
rect 2148 4321 2176 5578
rect 2134 4312 2190 4321
rect 2134 4247 2190 4256
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2042 3768 2098 3777
rect 2042 3703 2044 3712
rect 2096 3703 2098 3712
rect 2044 3674 2096 3680
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1858 1456 1914 1465
rect 1858 1391 1914 1400
rect 2148 800 2176 4082
rect 2240 3534 2268 6258
rect 2332 4146 2360 7414
rect 2424 6934 2452 12600
rect 2608 9654 2636 12718
rect 2686 12679 2742 12688
rect 2700 11694 2728 12679
rect 2792 11694 2820 13654
rect 2884 12481 2912 14350
rect 2976 13433 3004 14470
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3068 13530 3096 14418
rect 3160 13920 3188 16526
rect 3252 16425 3280 16526
rect 3238 16416 3294 16425
rect 3238 16351 3294 16360
rect 3344 16250 3372 16662
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3252 15094 3280 15370
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3804 15162 3832 15438
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3436 14328 3464 15030
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3344 14300 3464 14328
rect 3160 13892 3280 13920
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2962 13424 3018 13433
rect 2962 13359 3018 13368
rect 3160 12832 3188 13738
rect 3068 12804 3188 12832
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2870 12472 2926 12481
rect 2976 12442 3004 12582
rect 2870 12407 2926 12416
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 10606 2820 11630
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2976 10538 3004 11698
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2792 9110 2820 9862
rect 2976 9586 3004 9998
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 8566 2636 8978
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2596 8560 2648 8566
rect 2884 8514 2912 8910
rect 2596 8502 2648 8508
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 3126 2268 3470
rect 2424 3466 2452 4014
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2228 3120 2280 3126
rect 2228 3062 2280 3068
rect 2410 2952 2466 2961
rect 2410 2887 2466 2896
rect 2424 800 2452 2887
rect 2516 1834 2544 8230
rect 2608 7886 2636 8502
rect 2700 8486 2912 8514
rect 2976 8514 3004 9522
rect 3068 9489 3096 12804
rect 3146 11656 3202 11665
rect 3146 11591 3148 11600
rect 3200 11591 3202 11600
rect 3148 11562 3200 11568
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10713 3188 11086
rect 3146 10704 3202 10713
rect 3146 10639 3202 10648
rect 3146 10160 3202 10169
rect 3146 10095 3148 10104
rect 3200 10095 3202 10104
rect 3148 10066 3200 10072
rect 3054 9480 3110 9489
rect 3054 9415 3110 9424
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9178 3188 9318
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8634 3188 8774
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2976 8486 3188 8514
rect 2700 8090 2728 8486
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 7970 2820 8366
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2700 7942 2820 7970
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2700 7154 2728 7942
rect 2884 7546 2912 8298
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 8090 3004 8230
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2976 7478 3004 7754
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2700 7126 2912 7154
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2608 5001 2636 5238
rect 2594 4992 2650 5001
rect 2594 4927 2650 4936
rect 2700 3641 2728 6870
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2792 5166 2820 6802
rect 2884 5658 2912 7126
rect 2976 6254 3004 7278
rect 3068 6662 3096 8298
rect 3160 8242 3188 8486
rect 3252 8401 3280 13892
rect 3344 8906 3372 14300
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 10266 3464 10474
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3514 9480 3570 9489
rect 3514 9415 3516 9424
rect 3568 9415 3570 9424
rect 3516 9386 3568 9392
rect 3620 9042 3648 9522
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3804 8906 3832 14962
rect 3896 12374 3924 15914
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 3988 11801 4016 16594
rect 4080 15026 4108 17054
rect 4264 16182 4292 17836
rect 4540 17746 4568 19200
rect 4816 18086 4844 19200
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 5184 18018 5212 19200
rect 5172 18012 5224 18018
rect 5172 17954 5224 17960
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 5552 17542 5580 19200
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4344 16040 4396 16046
rect 4342 16008 4344 16017
rect 4396 16008 4398 16017
rect 4342 15943 4398 15952
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4066 14512 4122 14521
rect 4066 14447 4122 14456
rect 4080 13802 4108 14447
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4172 13190 4200 15846
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 13841 4292 14758
rect 4250 13832 4306 13841
rect 4250 13767 4306 13776
rect 4356 13734 4384 15302
rect 4448 14958 4476 16730
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14482 4476 14758
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4250 13016 4306 13025
rect 4250 12951 4252 12960
rect 4304 12951 4306 12960
rect 4252 12922 4304 12928
rect 4068 12912 4120 12918
rect 4120 12860 4292 12866
rect 4068 12854 4292 12860
rect 4080 12838 4292 12854
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3896 11354 3924 11562
rect 3974 11520 4030 11529
rect 3974 11455 4030 11464
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3988 11218 4016 11455
rect 4080 11354 4108 12174
rect 4172 11762 4200 12378
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3882 10024 3938 10033
rect 3882 9959 3938 9968
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3896 8401 3924 9959
rect 3238 8392 3294 8401
rect 3238 8327 3294 8336
rect 3882 8392 3938 8401
rect 3882 8327 3938 8336
rect 3884 8288 3936 8294
rect 3330 8256 3386 8265
rect 3160 8214 3330 8242
rect 3884 8230 3936 8236
rect 3330 8191 3386 8200
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7546 3280 7822
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3238 7304 3294 7313
rect 3344 7274 3372 8191
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3804 7342 3832 7822
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3238 7239 3294 7248
rect 3332 7268 3384 7274
rect 3252 6934 3280 7239
rect 3332 7210 3384 7216
rect 3804 7206 3832 7278
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3528 6798 3556 7142
rect 3790 6896 3846 6905
rect 3790 6831 3846 6840
rect 3240 6792 3292 6798
rect 3238 6760 3240 6769
rect 3516 6792 3568 6798
rect 3292 6760 3294 6769
rect 3238 6695 3294 6704
rect 3344 6740 3516 6746
rect 3344 6734 3568 6740
rect 3344 6718 3556 6734
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 3160 5914 3188 6598
rect 3344 6186 3372 6718
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3804 6254 3832 6831
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3436 5710 3464 5850
rect 3240 5704 3292 5710
rect 2884 5630 3188 5658
rect 3424 5704 3476 5710
rect 3240 5646 3292 5652
rect 3344 5664 3424 5692
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 3738 2820 4422
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2686 3632 2742 3641
rect 2686 3567 2742 3576
rect 2778 3088 2834 3097
rect 2778 3023 2834 3032
rect 2504 1828 2556 1834
rect 2504 1770 2556 1776
rect 2792 800 2820 3023
rect 2884 2922 2912 4150
rect 2976 3058 3004 5510
rect 3054 4720 3110 4729
rect 3054 4655 3056 4664
rect 3108 4655 3110 4664
rect 3056 4626 3108 4632
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 2884 513 2912 2450
rect 3068 2038 3096 3878
rect 3160 3505 3188 5630
rect 3252 4554 3280 5646
rect 3344 5370 3372 5664
rect 3424 5646 3476 5652
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3332 5364 3384 5370
rect 3804 5352 3832 6190
rect 3332 5306 3384 5312
rect 3712 5324 3832 5352
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3620 5001 3648 5102
rect 3606 4992 3662 5001
rect 3606 4927 3662 4936
rect 3712 4622 3740 5324
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3424 4616 3476 4622
rect 3344 4576 3424 4604
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3252 3738 3280 4218
rect 3344 3913 3372 4576
rect 3424 4558 3476 4564
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3700 3936 3752 3942
rect 3330 3904 3386 3913
rect 3700 3878 3752 3884
rect 3330 3839 3386 3848
rect 3712 3738 3740 3878
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3146 3496 3202 3505
rect 3330 3496 3386 3505
rect 3146 3431 3202 3440
rect 3252 3454 3330 3482
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 3252 1816 3280 3454
rect 3436 3466 3464 3606
rect 3330 3431 3386 3440
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3804 3346 3832 5034
rect 3896 4321 3924 8230
rect 3988 6304 4016 11154
rect 4172 10742 4200 11494
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 4080 9450 4108 9551
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 4172 9217 4200 9930
rect 4264 9450 4292 12838
rect 4356 12442 4384 13262
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4342 11928 4398 11937
rect 4342 11863 4398 11872
rect 4356 11354 4384 11863
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10606 4384 11086
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4158 9208 4214 9217
rect 4356 9178 4384 10542
rect 4448 9586 4476 13126
rect 4540 12374 4568 14350
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4540 11132 4568 12310
rect 4632 11558 4660 16050
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15638 5212 15846
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5368 15570 5396 16594
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 15570 5488 16390
rect 5552 15706 5580 16730
rect 5828 16572 5856 19200
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 6012 17066 6040 17750
rect 6196 17338 6224 19200
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 5908 16584 5960 16590
rect 5828 16544 5908 16572
rect 5908 16526 5960 16532
rect 6288 16522 6316 17138
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4816 14929 4844 14962
rect 4896 14952 4948 14958
rect 4802 14920 4858 14929
rect 4896 14894 4948 14900
rect 4802 14855 4858 14864
rect 4908 14226 4936 14894
rect 5000 14890 5028 15438
rect 5368 15366 5396 15506
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5460 14958 5488 15506
rect 5630 15056 5686 15065
rect 5630 14991 5686 15000
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5000 14346 5028 14826
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5092 14226 5120 14282
rect 4908 14198 5120 14226
rect 4908 13938 4936 14198
rect 5276 13977 5304 14418
rect 5460 14346 5488 14418
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5262 13968 5318 13977
rect 4896 13932 4948 13938
rect 5262 13903 5318 13912
rect 4896 13874 4948 13880
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13462 4844 13670
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4724 13297 4752 13330
rect 4710 13288 4766 13297
rect 4710 13223 4766 13232
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4724 12714 4752 12922
rect 4908 12918 4936 13874
rect 5460 13326 5488 14282
rect 5552 13802 5580 14418
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 4804 12912 4856 12918
rect 4802 12880 4804 12889
rect 4896 12912 4948 12918
rect 4856 12880 4858 12889
rect 5092 12889 5120 13262
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4896 12854 4948 12860
rect 5078 12880 5134 12889
rect 4802 12815 4858 12824
rect 5078 12815 5134 12824
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 5092 12442 5120 12815
rect 5184 12782 5212 13126
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5000 12322 5028 12378
rect 5460 12322 5488 12718
rect 5644 12356 5672 14991
rect 5736 13870 5764 16050
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5828 14822 5856 15506
rect 5816 14816 5868 14822
rect 6288 14793 6316 16458
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 16046 6500 16390
rect 6564 16153 6592 19200
rect 6932 17762 6960 19200
rect 7208 17950 7236 19200
rect 7196 17944 7248 17950
rect 7196 17886 7248 17892
rect 6932 17734 7052 17762
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6932 17338 6960 17614
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6550 16144 6606 16153
rect 6550 16079 6606 16088
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 5816 14758 5868 14764
rect 6274 14784 6330 14793
rect 5886 14716 6182 14736
rect 6274 14719 6330 14728
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6012 14385 6040 14418
rect 5998 14376 6054 14385
rect 5998 14311 6054 14320
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5920 13025 5948 13330
rect 5906 13016 5962 13025
rect 5906 12951 5962 12960
rect 6288 12918 6316 13738
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 5644 12328 5856 12356
rect 5000 12294 5488 12322
rect 5540 12232 5592 12238
rect 5170 12200 5226 12209
rect 5540 12174 5592 12180
rect 5170 12135 5226 12144
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4620 11280 4672 11286
rect 4618 11248 4620 11257
rect 4672 11248 4674 11257
rect 4618 11183 4674 11192
rect 4540 11104 4752 11132
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4158 9143 4214 9152
rect 4344 9172 4396 9178
rect 4172 9042 4200 9143
rect 4344 9114 4396 9120
rect 4540 9081 4568 10134
rect 4724 9738 4752 11104
rect 4816 10674 4844 11630
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11286 4936 11494
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 5184 10742 5212 12135
rect 5354 11928 5410 11937
rect 5552 11898 5580 12174
rect 5354 11863 5410 11872
rect 5540 11892 5592 11898
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5276 10674 5304 11086
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 4816 9926 4844 10610
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 4804 9920 4856 9926
rect 4856 9868 4936 9874
rect 4804 9862 4936 9868
rect 4816 9846 4936 9862
rect 4724 9710 4844 9738
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4526 9072 4582 9081
rect 4160 9036 4212 9042
rect 4526 9007 4582 9016
rect 4620 9036 4672 9042
rect 4160 8978 4212 8984
rect 4620 8978 4672 8984
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4080 6497 4108 8842
rect 4342 8800 4398 8809
rect 4342 8735 4398 8744
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 4264 6390 4292 8434
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 3988 6276 4108 6304
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3882 4312 3938 4321
rect 3882 4247 3938 4256
rect 3882 3360 3938 3369
rect 3804 3318 3882 3346
rect 3421 3292 3717 3312
rect 3882 3295 3938 3304
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3988 3058 4016 6122
rect 4080 6100 4108 6276
rect 4080 6072 4292 6100
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 4282 4108 5510
rect 4264 5409 4292 6072
rect 4250 5400 4306 5409
rect 4250 5335 4306 5344
rect 4158 4992 4214 5001
rect 4158 4927 4214 4936
rect 4172 4486 4200 4927
rect 4264 4865 4292 5335
rect 4250 4856 4306 4865
rect 4250 4791 4306 4800
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 4250 4176 4306 4185
rect 4250 4111 4252 4120
rect 4080 3942 4108 4111
rect 4304 4111 4306 4120
rect 4252 4082 4304 4088
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4080 3602 4108 3878
rect 4172 3777 4200 3878
rect 4158 3768 4214 3777
rect 4158 3703 4214 3712
rect 4356 3618 4384 8735
rect 4632 8634 4660 8978
rect 4724 8634 4752 9318
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4448 7857 4476 7890
rect 4434 7848 4490 7857
rect 4434 7783 4490 7792
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 6730 4476 7686
rect 4540 7206 4568 8434
rect 4632 7478 4660 8570
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4448 5370 4476 5578
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4448 4729 4476 5034
rect 4434 4720 4490 4729
rect 4434 4655 4490 4664
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4448 3754 4476 4082
rect 4540 4010 4568 5646
rect 4618 4856 4674 4865
rect 4618 4791 4674 4800
rect 4632 4690 4660 4791
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4448 3726 4568 3754
rect 4068 3596 4120 3602
rect 4356 3590 4476 3618
rect 4068 3538 4120 3544
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3058 4200 3334
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4264 2938 4292 3402
rect 4448 3398 4476 3590
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4540 3346 4568 3726
rect 4632 3602 4660 4422
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4724 3534 4752 7754
rect 4816 7449 4844 9710
rect 4908 9518 4936 9846
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 9110 4936 9454
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5184 9178 5212 9386
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 5078 8528 5134 8537
rect 5078 8463 5134 8472
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4802 7440 4858 7449
rect 4802 7375 4858 7384
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4816 6730 4844 7278
rect 4908 7041 4936 7822
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 4894 7032 4950 7041
rect 4894 6967 4950 6976
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 6254 4844 6666
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 6118 4844 6190
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5778 4844 6054
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4816 4729 4844 5102
rect 4802 4720 4858 4729
rect 4802 4655 4858 4664
rect 4816 4060 4844 4655
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4908 4214 4936 4558
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4896 4072 4948 4078
rect 4816 4032 4896 4060
rect 4896 4014 4948 4020
rect 4908 3602 4936 4014
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4908 3346 4936 3538
rect 5000 3466 5028 7754
rect 5092 7750 5120 8463
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5184 7750 5212 8298
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6633 5120 6734
rect 5078 6624 5134 6633
rect 5078 6559 5134 6568
rect 5184 6458 5212 7210
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5184 5914 5212 6122
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5078 5808 5134 5817
rect 5276 5794 5304 10474
rect 5368 6905 5396 11863
rect 5540 11834 5592 11840
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11286 5764 11494
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5446 10704 5502 10713
rect 5446 10639 5502 10648
rect 5460 10538 5488 10639
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 5644 9722 5672 10474
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 7818 5488 9454
rect 5552 8945 5580 9658
rect 5630 9208 5686 9217
rect 5630 9143 5686 9152
rect 5538 8936 5594 8945
rect 5538 8871 5594 8880
rect 5644 8838 5672 9143
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5632 8424 5684 8430
rect 5736 8412 5764 9998
rect 5684 8384 5764 8412
rect 5632 8366 5684 8372
rect 5540 8288 5592 8294
rect 5538 8256 5540 8265
rect 5592 8256 5594 8265
rect 5538 8191 5594 8200
rect 5644 7954 5672 8366
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5354 6896 5410 6905
rect 5354 6831 5410 6840
rect 5276 5766 5396 5794
rect 5078 5743 5134 5752
rect 5092 3482 5120 5743
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5184 5098 5212 5646
rect 5276 5545 5304 5646
rect 5262 5536 5318 5545
rect 5262 5471 5318 5480
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5184 3913 5212 5034
rect 5262 4720 5318 4729
rect 5262 4655 5264 4664
rect 5316 4655 5318 4664
rect 5264 4626 5316 4632
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5276 4457 5304 4490
rect 5262 4448 5318 4457
rect 5262 4383 5318 4392
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5170 3904 5226 3913
rect 5170 3839 5226 3848
rect 5184 3738 5212 3839
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3670 5304 3946
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 4988 3460 5040 3466
rect 5092 3454 5212 3482
rect 4988 3402 5040 3408
rect 5080 3392 5132 3398
rect 4540 3318 4660 3346
rect 4908 3318 5028 3346
rect 5080 3334 5132 3340
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4448 3097 4476 3130
rect 4434 3088 4490 3097
rect 4434 3023 4490 3032
rect 4172 2910 4292 2938
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3514 2000 3570 2009
rect 3514 1935 3570 1944
rect 3792 1964 3844 1970
rect 3160 1788 3280 1816
rect 3160 800 3188 1788
rect 3528 800 3556 1935
rect 3792 1906 3844 1912
rect 3804 800 3832 1906
rect 4172 800 4200 2910
rect 4448 2650 4476 2926
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4540 800 4568 3130
rect 4632 3058 4660 3318
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4908 2650 4936 3062
rect 5000 2990 5028 3318
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5000 2310 5028 2926
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5092 1442 5120 3334
rect 5184 3194 5212 3454
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5368 3074 5396 5766
rect 4816 1414 5120 1442
rect 5184 3046 5396 3074
rect 4816 800 4844 1414
rect 5184 800 5212 3046
rect 5460 2990 5488 7142
rect 5540 6928 5592 6934
rect 5538 6896 5540 6905
rect 5592 6896 5594 6905
rect 5538 6831 5594 6840
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5552 5098 5580 6734
rect 5644 6730 5672 7890
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5552 5001 5580 5034
rect 5724 5024 5776 5030
rect 5538 4992 5594 5001
rect 5724 4966 5776 4972
rect 5538 4927 5594 4936
rect 5736 4729 5764 4966
rect 5722 4720 5778 4729
rect 5540 4684 5592 4690
rect 5722 4655 5778 4664
rect 5540 4626 5592 4632
rect 5552 3398 5580 4626
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5722 4448 5778 4457
rect 5644 3602 5672 4422
rect 5722 4383 5778 4392
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5552 800 5580 3130
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2650 5672 2790
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5736 2446 5764 4383
rect 5828 2632 5856 12328
rect 6288 11642 6316 12378
rect 6380 11898 6408 15846
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6458 14648 6514 14657
rect 6458 14583 6514 14592
rect 6472 12152 6500 14583
rect 6564 12889 6592 15302
rect 6656 14521 6684 16594
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6748 16454 6776 16526
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6840 16250 6868 16594
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6932 15450 6960 16050
rect 7024 15609 7052 17734
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7010 15600 7066 15609
rect 7010 15535 7066 15544
rect 6932 15422 7052 15450
rect 6920 14952 6972 14958
rect 6826 14920 6882 14929
rect 6920 14894 6972 14900
rect 6826 14855 6882 14864
rect 6642 14512 6698 14521
rect 6840 14482 6868 14855
rect 6642 14447 6698 14456
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6932 14414 6960 14894
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 7024 14362 7052 15422
rect 7116 14464 7144 17070
rect 7208 16561 7236 17070
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7194 16552 7250 16561
rect 7194 16487 7250 16496
rect 7208 15910 7236 16487
rect 7392 15910 7420 17002
rect 7196 15904 7248 15910
rect 7380 15904 7432 15910
rect 7196 15846 7248 15852
rect 7378 15872 7380 15881
rect 7432 15872 7434 15881
rect 7208 15473 7236 15846
rect 7378 15807 7434 15816
rect 7484 15706 7512 17138
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7194 15464 7250 15473
rect 7194 15399 7250 15408
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7116 14436 7236 14464
rect 7102 14376 7158 14385
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13870 6776 14214
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6736 13864 6788 13870
rect 6642 13832 6698 13841
rect 6736 13806 6788 13812
rect 6642 13767 6698 13776
rect 6656 13433 6684 13767
rect 6642 13424 6698 13433
rect 6642 13359 6698 13368
rect 6550 12880 6606 12889
rect 6550 12815 6606 12824
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6748 12617 6776 12718
rect 6840 12628 6868 13942
rect 6932 13870 6960 14350
rect 7024 14334 7102 14362
rect 7102 14311 7158 14320
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 12782 6960 13806
rect 7116 13802 7144 14311
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6920 12776 6972 12782
rect 6972 12736 7052 12764
rect 6920 12718 6972 12724
rect 6734 12608 6790 12617
rect 6840 12600 6960 12628
rect 6734 12543 6790 12552
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 12232 6696 12238
rect 6642 12200 6644 12209
rect 6696 12200 6698 12209
rect 6472 12124 6592 12152
rect 6642 12135 6698 12144
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6196 11626 6316 11642
rect 6184 11620 6316 11626
rect 6236 11614 6316 11620
rect 6184 11562 6236 11568
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6196 9364 6224 10066
rect 6288 9518 6316 11494
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6368 9376 6420 9382
rect 6196 9336 6316 9364
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 6288 8906 6316 9336
rect 6368 9318 6420 9324
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6288 8634 6316 8842
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6274 8256 6330 8265
rect 5886 8188 6182 8208
rect 6274 8191 6330 8200
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 6288 7954 6316 8191
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6104 6186 6132 6870
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 5030 6316 5714
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6182 4448 6238 4457
rect 6104 4078 6132 4422
rect 6182 4383 6238 4392
rect 6196 4214 6224 4383
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6288 4010 6316 4966
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 6380 3670 6408 9318
rect 6472 9178 6500 10406
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6104 3194 6132 3606
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 5828 2604 6224 2632
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6012 2106 6040 2450
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 5828 800 5856 1838
rect 6196 800 6224 2604
rect 6380 1902 6408 3470
rect 6472 3194 6500 5102
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6368 1896 6420 1902
rect 6368 1838 6420 1844
rect 6564 800 6592 12124
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6656 11558 6684 11630
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6748 11354 6776 12242
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6840 11218 6868 11698
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 10674 6868 11154
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6656 10198 6684 10406
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6840 10044 6868 10610
rect 6932 10538 6960 12600
rect 7024 12306 7052 12736
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7116 12442 7144 12650
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7208 11626 7236 14436
rect 7392 13530 7420 15302
rect 7484 14958 7512 15642
rect 7576 15366 7604 19200
rect 7944 17241 7972 19200
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7930 17232 7986 17241
rect 7930 17167 7986 17176
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7484 13394 7512 13806
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7564 13388 7616 13394
rect 7668 13376 7696 16458
rect 7760 14249 7788 16594
rect 7852 16114 7880 16662
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7944 15586 7972 16934
rect 8036 16794 8064 17274
rect 8220 17218 8248 19200
rect 8588 17649 8616 19200
rect 8574 17640 8630 17649
rect 8574 17575 8630 17584
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8220 17202 8432 17218
rect 8220 17196 8444 17202
rect 8220 17190 8392 17196
rect 8392 17138 8444 17144
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8668 16992 8720 16998
rect 8390 16960 8446 16969
rect 8668 16934 8720 16940
rect 8390 16895 8446 16904
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8404 16658 8432 16895
rect 8574 16688 8630 16697
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8392 16652 8444 16658
rect 8574 16623 8630 16632
rect 8392 16594 8444 16600
rect 8024 16584 8076 16590
rect 8312 16561 8340 16594
rect 8588 16590 8616 16623
rect 8576 16584 8628 16590
rect 8024 16526 8076 16532
rect 8298 16552 8354 16561
rect 8036 15745 8064 16526
rect 8576 16526 8628 16532
rect 8298 16487 8354 16496
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8022 15736 8078 15745
rect 8022 15671 8078 15680
rect 8116 15700 8168 15706
rect 7852 15558 7972 15586
rect 7852 14482 7880 15558
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7746 14240 7802 14249
rect 7746 14175 7802 14184
rect 7760 13802 7788 14175
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7852 13462 7880 13942
rect 7944 13530 7972 15438
rect 8036 14929 8064 15671
rect 8116 15642 8168 15648
rect 8022 14920 8078 14929
rect 8022 14855 8078 14864
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8036 13569 8064 14418
rect 8128 13938 8156 15642
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8022 13560 8078 13569
rect 7932 13524 7984 13530
rect 8022 13495 8078 13504
rect 7932 13466 7984 13472
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7616 13348 7696 13376
rect 7564 13330 7616 13336
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12646 7880 13126
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 8036 12753 8064 12854
rect 8128 12850 8156 13874
rect 8220 13462 8248 15506
rect 8312 15502 8340 15982
rect 8496 15881 8524 15982
rect 8482 15872 8538 15881
rect 8482 15807 8538 15816
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8300 15496 8352 15502
rect 8588 15473 8616 15506
rect 8300 15438 8352 15444
rect 8574 15464 8630 15473
rect 8574 15399 8630 15408
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8298 14784 8354 14793
rect 8298 14719 8354 14728
rect 8312 14414 8340 14719
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8496 14346 8524 14826
rect 8588 14550 8616 14962
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8312 13870 8340 13942
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8588 13258 8616 13738
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8300 12776 8352 12782
rect 8022 12744 8078 12753
rect 8022 12679 8078 12688
rect 8220 12736 8300 12764
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 8036 12374 8064 12679
rect 8220 12442 8248 12736
rect 8300 12718 8352 12724
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 7378 12200 7434 12209
rect 7378 12135 7434 12144
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7208 10266 7236 10474
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 6920 10056 6972 10062
rect 6840 10016 6920 10044
rect 6840 9586 6868 10016
rect 6920 9998 6972 10004
rect 7392 9738 7420 12135
rect 8220 11898 8248 12378
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7930 11656 7986 11665
rect 7930 11591 7986 11600
rect 7470 11112 7526 11121
rect 7470 11047 7526 11056
rect 7300 9710 7420 9738
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 7194 9480 7250 9489
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6656 7993 6684 8502
rect 6642 7984 6698 7993
rect 6642 7919 6698 7928
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5098 6684 5646
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6642 4856 6698 4865
rect 6642 4791 6644 4800
rect 6696 4791 6698 4800
rect 6644 4762 6696 4768
rect 6748 3720 6776 9454
rect 7104 9444 7156 9450
rect 7194 9415 7250 9424
rect 7104 9386 7156 9392
rect 7116 9110 7144 9386
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 7410 6868 8366
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 6254 6868 7346
rect 6932 7206 6960 7686
rect 7208 7313 7236 9415
rect 7194 7304 7250 7313
rect 7012 7268 7064 7274
rect 7194 7239 7250 7248
rect 7012 7210 7064 7216
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 7024 7041 7052 7210
rect 7010 7032 7066 7041
rect 7010 6967 7066 6976
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5098 6960 5510
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6656 3692 6776 3720
rect 6656 3534 6684 3692
rect 6840 3670 6868 4422
rect 6932 4185 6960 4762
rect 6918 4176 6974 4185
rect 6918 4111 6974 4120
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6932 3602 6960 4111
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6656 2514 6684 3334
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6748 2446 6776 3538
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 2582 6868 3334
rect 7024 2854 7052 6967
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6458 7236 6598
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7208 6202 7236 6394
rect 7116 6186 7236 6202
rect 7104 6180 7236 6186
rect 7156 6174 7236 6180
rect 7104 6122 7156 6128
rect 7300 5817 7328 9710
rect 7286 5808 7342 5817
rect 7104 5772 7156 5778
rect 7156 5732 7236 5760
rect 7286 5743 7342 5752
rect 7380 5772 7432 5778
rect 7104 5714 7156 5720
rect 7208 5030 7236 5732
rect 7380 5714 7432 5720
rect 7286 5264 7342 5273
rect 7392 5250 7420 5714
rect 7484 5352 7512 11047
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7852 9382 7880 10678
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7746 9208 7802 9217
rect 7746 9143 7802 9152
rect 7760 8974 7788 9143
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7748 8968 7800 8974
rect 7576 8928 7748 8956
rect 7576 7954 7604 8928
rect 7748 8910 7800 8916
rect 7852 8401 7880 9046
rect 7838 8392 7894 8401
rect 7838 8327 7894 8336
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7576 7392 7604 7890
rect 7840 7404 7892 7410
rect 7576 7364 7840 7392
rect 7760 6866 7788 7364
rect 7840 7346 7892 7352
rect 7564 6860 7616 6866
rect 7748 6860 7800 6866
rect 7616 6820 7696 6848
rect 7564 6802 7616 6808
rect 7668 5778 7696 6820
rect 7748 6802 7800 6808
rect 7838 6624 7894 6633
rect 7838 6559 7894 6568
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7484 5324 7604 5352
rect 7470 5264 7526 5273
rect 7392 5222 7470 5250
rect 7286 5199 7342 5208
rect 7470 5199 7526 5208
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4622 7236 4966
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7208 4010 7236 4558
rect 7300 4010 7328 5199
rect 7576 4298 7604 5324
rect 7760 5030 7788 6054
rect 7852 5681 7880 6559
rect 7838 5672 7894 5681
rect 7838 5607 7894 5616
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7484 4270 7604 4298
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7102 3904 7158 3913
rect 7102 3839 7158 3848
rect 7116 3233 7144 3839
rect 7208 3534 7236 3946
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7102 3224 7158 3233
rect 7102 3159 7158 3168
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6918 2408 6974 2417
rect 6918 2343 6974 2352
rect 6932 800 6960 2343
rect 7300 1698 7328 2450
rect 7484 1970 7512 4270
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7288 1692 7340 1698
rect 7288 1634 7340 1640
rect 7196 1624 7248 1630
rect 7196 1566 7248 1572
rect 7208 800 7236 1566
rect 7576 800 7604 3878
rect 7760 2922 7788 4966
rect 7944 4128 7972 11591
rect 8036 8809 8064 11766
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8588 11082 8616 11222
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8680 10742 8708 16934
rect 8772 16425 8800 17002
rect 8956 16810 8984 19200
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9048 16998 9076 17818
rect 9232 17066 9260 19200
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8956 16782 9168 16810
rect 9140 16590 9168 16782
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9324 16697 9352 16730
rect 9310 16688 9366 16697
rect 9310 16623 9366 16632
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9416 16522 9444 18022
rect 9496 18012 9548 18018
rect 9496 17954 9548 17960
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 8758 16416 8814 16425
rect 8758 16351 8814 16360
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8772 15162 8800 15574
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8772 13802 8800 14826
rect 8864 14249 8892 16050
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 8850 14240 8906 14249
rect 8850 14175 8906 14184
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8772 12442 8800 13466
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8864 13025 8892 13330
rect 8850 13016 8906 13025
rect 8850 12951 8906 12960
rect 8850 12880 8906 12889
rect 8850 12815 8906 12824
rect 8864 12442 8892 12815
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8956 12288 8984 15370
rect 8772 12260 8984 12288
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8116 10464 8168 10470
rect 8114 10432 8116 10441
rect 8772 10452 8800 12260
rect 8942 12200 8998 12209
rect 8942 12135 8998 12144
rect 8850 11248 8906 11257
rect 8850 11183 8906 11192
rect 8168 10432 8170 10441
rect 8114 10367 8170 10376
rect 8680 10424 8800 10452
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8576 9648 8628 9654
rect 8482 9616 8538 9625
rect 8680 9636 8708 10424
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8628 9608 8708 9636
rect 8576 9590 8628 9596
rect 8482 9551 8538 9560
rect 8496 9518 8524 9551
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9110 8248 9318
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8022 8800 8078 8809
rect 8022 8735 8078 8744
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8680 8634 8708 9046
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8220 7954 8248 8502
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8680 7818 8708 8230
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8772 7721 8800 10202
rect 8864 8974 8892 11183
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8864 8362 8892 8570
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8758 7712 8814 7721
rect 8352 7644 8648 7664
rect 8758 7647 8814 7656
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 7002 8156 7142
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8220 6934 8248 7414
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 6934 8708 7346
rect 8772 7342 8800 7647
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8668 6928 8720 6934
rect 8864 6905 8892 7890
rect 8668 6870 8720 6876
rect 8850 6896 8906 6905
rect 8022 6488 8078 6497
rect 8220 6458 8248 6870
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8022 6423 8078 6432
rect 8208 6452 8260 6458
rect 8036 6202 8064 6423
rect 8208 6394 8260 6400
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8036 6174 8248 6202
rect 8220 5778 8248 6174
rect 8496 6089 8524 6326
rect 8576 6248 8628 6254
rect 8680 6236 8708 6870
rect 8850 6831 8906 6840
rect 8628 6208 8708 6236
rect 8760 6248 8812 6254
rect 8576 6190 8628 6196
rect 8760 6190 8812 6196
rect 8668 6112 8720 6118
rect 8482 6080 8538 6089
rect 8772 6089 8800 6190
rect 8668 6054 8720 6060
rect 8758 6080 8814 6089
rect 8482 6015 8538 6024
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8024 5296 8076 5302
rect 8022 5264 8024 5273
rect 8076 5264 8078 5273
rect 8022 5199 8078 5208
rect 8022 4992 8078 5001
rect 8022 4927 8078 4936
rect 7852 4100 7972 4128
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7852 2854 7880 4100
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7944 3097 7972 3878
rect 7930 3088 7986 3097
rect 7930 3023 7986 3032
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7852 2514 7880 2790
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 7852 1766 7880 2450
rect 7932 2032 7984 2038
rect 8036 2020 8064 4927
rect 8128 3194 8156 5646
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8220 5545 8248 5578
rect 8206 5536 8262 5545
rect 8206 5471 8262 5480
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8404 5166 8432 5238
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4570 8340 4626
rect 8220 4542 8340 4570
rect 8220 4282 8248 4542
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8220 2990 8248 4014
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8680 3176 8708 6054
rect 8758 6015 8814 6024
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8588 3148 8708 3176
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8220 2038 8248 2926
rect 8588 2446 8616 3148
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 7984 1992 8064 2020
rect 8208 2032 8260 2038
rect 7932 1974 7984 1980
rect 8208 1974 8260 1980
rect 7840 1760 7892 1766
rect 7840 1702 7892 1708
rect 7944 800 7972 1974
rect 8680 1970 8708 2450
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8208 1760 8260 1766
rect 8208 1702 8260 1708
rect 8220 800 8248 1702
rect 8772 1630 8800 4558
rect 8864 2836 8892 6831
rect 8956 2990 8984 12135
rect 9048 10713 9076 16458
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 9140 15026 9168 15370
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9232 14890 9260 15982
rect 9324 15337 9352 15982
rect 9508 15910 9536 17954
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9310 15328 9366 15337
rect 9310 15263 9366 15272
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9324 14929 9352 14962
rect 9310 14920 9366 14929
rect 9220 14884 9272 14890
rect 9310 14855 9366 14864
rect 9220 14826 9272 14832
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9034 10704 9090 10713
rect 9034 10639 9090 10648
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 8498 9076 10474
rect 9140 9217 9168 14554
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9232 9500 9260 14418
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9324 12714 9352 14010
rect 9416 13802 9444 15846
rect 9600 15638 9628 19200
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16522 9720 16934
rect 9784 16561 9812 17070
rect 9770 16552 9826 16561
rect 9680 16516 9732 16522
rect 9770 16487 9826 16496
rect 9680 16458 9732 16464
rect 9876 16454 9904 17546
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9968 16250 9996 19200
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9864 16040 9916 16046
rect 9784 16000 9864 16028
rect 9680 15904 9732 15910
rect 9678 15872 9680 15881
rect 9732 15872 9734 15881
rect 9678 15807 9734 15816
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9508 13530 9536 15506
rect 9678 15192 9734 15201
rect 9784 15178 9812 16000
rect 9864 15982 9916 15988
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9876 15201 9904 15846
rect 9954 15736 10010 15745
rect 9954 15671 10010 15680
rect 9968 15502 9996 15671
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9734 15150 9812 15178
rect 9862 15192 9918 15201
rect 9678 15127 9734 15136
rect 9862 15127 9918 15136
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9586 14920 9642 14929
rect 9586 14855 9642 14864
rect 9600 14822 9628 14855
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9784 14550 9812 14962
rect 10060 14770 10088 16662
rect 9968 14742 10088 14770
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9600 14074 9628 14418
rect 9692 14113 9720 14418
rect 9772 14408 9824 14414
rect 9864 14408 9916 14414
rect 9772 14350 9824 14356
rect 9862 14376 9864 14385
rect 9916 14376 9918 14385
rect 9678 14104 9734 14113
rect 9588 14068 9640 14074
rect 9784 14074 9812 14350
rect 9862 14311 9918 14320
rect 9862 14240 9918 14249
rect 9862 14175 9918 14184
rect 9678 14039 9734 14048
rect 9772 14068 9824 14074
rect 9588 14010 9640 14016
rect 9772 14010 9824 14016
rect 9770 13968 9826 13977
rect 9770 13903 9826 13912
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9416 12306 9444 13330
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9312 12232 9364 12238
rect 9310 12200 9312 12209
rect 9364 12200 9366 12209
rect 9310 12135 9366 12144
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9324 10470 9352 11562
rect 9416 10810 9444 12242
rect 9508 11558 9536 13126
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9600 11937 9628 12650
rect 9692 12442 9720 13670
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9586 11928 9642 11937
rect 9586 11863 9642 11872
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 9738 9352 10406
rect 9416 10266 9444 10474
rect 9494 10296 9550 10305
rect 9404 10260 9456 10266
rect 9494 10231 9550 10240
rect 9404 10202 9456 10208
rect 9508 10198 9536 10231
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9494 9752 9550 9761
rect 9324 9710 9494 9738
rect 9494 9687 9550 9696
rect 9508 9586 9536 9687
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9600 9518 9628 11562
rect 9588 9512 9640 9518
rect 9232 9472 9444 9500
rect 9312 9376 9364 9382
rect 9310 9344 9312 9353
rect 9364 9344 9366 9353
rect 9310 9279 9366 9288
rect 9126 9208 9182 9217
rect 9126 9143 9182 9152
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9126 8256 9182 8265
rect 9126 8191 9182 8200
rect 9140 7886 9168 8191
rect 9232 7954 9260 9114
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9128 7880 9180 7886
rect 9416 7834 9444 9472
rect 9588 9454 9640 9460
rect 9600 9217 9628 9454
rect 9586 9208 9642 9217
rect 9692 9178 9720 12242
rect 9784 11665 9812 13903
rect 9876 13870 9904 14175
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9968 13530 9996 14742
rect 10046 14648 10102 14657
rect 10046 14583 10102 14592
rect 10060 14385 10088 14583
rect 10152 14550 10180 17070
rect 10244 16454 10272 17682
rect 10336 16969 10364 19200
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10520 17338 10548 17546
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10508 16992 10560 16998
rect 10322 16960 10378 16969
rect 10508 16934 10560 16940
rect 10322 16895 10378 16904
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10336 14958 10364 16594
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10336 14657 10364 14894
rect 10322 14648 10378 14657
rect 10322 14583 10378 14592
rect 10140 14544 10192 14550
rect 10428 14532 10456 16594
rect 10520 16590 10548 16934
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10520 15881 10548 15982
rect 10506 15872 10562 15881
rect 10506 15807 10562 15816
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10140 14486 10192 14492
rect 10244 14504 10456 14532
rect 10046 14376 10102 14385
rect 10046 14311 10102 14320
rect 10046 13696 10102 13705
rect 10046 13631 10102 13640
rect 9956 13524 10008 13530
rect 9876 13484 9956 13512
rect 9876 12481 9904 13484
rect 9956 13466 10008 13472
rect 10060 13326 10088 13631
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9968 13025 9996 13126
rect 9954 13016 10010 13025
rect 9954 12951 10010 12960
rect 10060 12889 10088 13262
rect 10046 12880 10102 12889
rect 10046 12815 10102 12824
rect 9862 12472 9918 12481
rect 9862 12407 9918 12416
rect 9956 12436 10008 12442
rect 9876 11762 9904 12407
rect 9956 12378 10008 12384
rect 9968 11898 9996 12378
rect 10048 12300 10100 12306
rect 10152 12288 10180 14486
rect 10244 13705 10272 14504
rect 10520 14482 10548 15438
rect 10612 14822 10640 19200
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17338 10732 17478
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10980 16980 11008 19200
rect 11152 17808 11204 17814
rect 11348 17762 11376 19200
rect 11152 17750 11204 17756
rect 10704 16952 11008 16980
rect 10704 16776 10732 16952
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 10704 16748 10916 16776
rect 10782 16552 10838 16561
rect 10782 16487 10838 16496
rect 10690 16280 10746 16289
rect 10690 16215 10746 16224
rect 10704 15570 10732 16215
rect 10796 16182 10824 16487
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10888 16114 10916 16748
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 11164 15688 11192 17750
rect 11256 17734 11376 17762
rect 11256 16726 11284 17734
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11072 15660 11192 15688
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10508 14476 10560 14482
rect 10336 14436 10508 14464
rect 10230 13696 10286 13705
rect 10230 13631 10286 13640
rect 10336 13240 10364 14436
rect 10508 14418 10560 14424
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10414 14104 10470 14113
rect 10414 14039 10416 14048
rect 10468 14039 10470 14048
rect 10416 14010 10468 14016
rect 10414 13968 10470 13977
rect 10414 13903 10470 13912
rect 10244 13212 10364 13240
rect 10244 12918 10272 13212
rect 10428 13138 10456 13903
rect 10520 13734 10548 14214
rect 10612 14113 10640 14758
rect 10704 14249 10732 15506
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 15065 11008 15438
rect 11072 15162 11100 15660
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10966 15056 11022 15065
rect 10966 14991 11022 15000
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 10968 14272 11020 14278
rect 10690 14240 10746 14249
rect 10968 14214 11020 14220
rect 10690 14175 10746 14184
rect 10598 14104 10654 14113
rect 10598 14039 10654 14048
rect 10980 14006 11008 14214
rect 11072 14074 11100 14447
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10336 13110 10456 13138
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10100 12260 10180 12288
rect 10048 12242 10100 12248
rect 10138 12200 10194 12209
rect 10048 12164 10100 12170
rect 10138 12135 10194 12144
rect 10048 12106 10100 12112
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10060 11762 10088 12106
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9770 11656 9826 11665
rect 9770 11591 9826 11600
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 10606 9812 11494
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9784 10130 9812 10542
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9784 9586 9812 10066
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9586 9143 9642 9152
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9494 8392 9550 8401
rect 9494 8327 9550 8336
rect 9588 8356 9640 8362
rect 9508 7954 9536 8327
rect 9588 8298 9640 8304
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9128 7822 9180 7828
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9048 6089 9076 7482
rect 9034 6080 9090 6089
rect 9034 6015 9090 6024
rect 9140 5681 9168 7822
rect 9232 7806 9444 7834
rect 9126 5672 9182 5681
rect 9126 5607 9182 5616
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8864 2808 8984 2836
rect 8760 1624 8812 1630
rect 8760 1566 8812 1572
rect 8576 1284 8628 1290
rect 8576 1226 8628 1232
rect 8588 800 8616 1226
rect 8956 800 8984 2808
rect 9048 1290 9076 3946
rect 9140 3618 9168 4422
rect 9232 3738 9260 7806
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 4690 9352 7686
rect 9600 7324 9628 8298
rect 9692 8090 9720 8774
rect 9784 8673 9812 8842
rect 9770 8664 9826 8673
rect 9770 8599 9826 8608
rect 9876 8378 9904 11562
rect 9968 9178 9996 11698
rect 10060 11218 10088 11698
rect 10152 11694 10180 12135
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10244 11014 10272 12582
rect 10336 11558 10364 13110
rect 10416 12980 10468 12986
rect 10468 12940 10548 12968
rect 10416 12922 10468 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10428 12753 10456 12786
rect 10414 12744 10470 12753
rect 10414 12679 10470 12688
rect 10520 11898 10548 12940
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 11393 10364 11494
rect 10322 11384 10378 11393
rect 10322 11319 10378 11328
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10232 11008 10284 11014
rect 10046 10976 10102 10985
rect 10232 10950 10284 10956
rect 10046 10911 10102 10920
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9784 8362 9904 8378
rect 9772 8356 9904 8362
rect 9824 8350 9904 8356
rect 9772 8298 9824 8304
rect 9864 8288 9916 8294
rect 9770 8256 9826 8265
rect 9864 8230 9916 8236
rect 9770 8191 9826 8200
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9784 8022 9812 8191
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9680 7336 9732 7342
rect 9600 7296 9680 7324
rect 9680 7278 9732 7284
rect 9876 7206 9904 8230
rect 9864 7200 9916 7206
rect 9586 7168 9642 7177
rect 9864 7142 9916 7148
rect 9586 7103 9642 7112
rect 9402 7032 9458 7041
rect 9402 6967 9458 6976
rect 9416 6798 9444 6967
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9140 3590 9260 3618
rect 9324 3602 9352 4626
rect 9508 4457 9536 5714
rect 9600 5545 9628 7103
rect 9862 6488 9918 6497
rect 9862 6423 9918 6432
rect 9876 6118 9904 6423
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9586 5536 9642 5545
rect 9586 5471 9642 5480
rect 9586 5400 9642 5409
rect 9586 5335 9642 5344
rect 9772 5364 9824 5370
rect 9600 4622 9628 5335
rect 9772 5306 9824 5312
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9692 4826 9720 5238
rect 9784 4842 9812 5306
rect 9876 5001 9904 6054
rect 9968 5710 9996 8978
rect 10060 8906 10088 10911
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 10266 10180 10610
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10152 9625 10180 10202
rect 10244 10130 10272 10474
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10138 9616 10194 9625
rect 10138 9551 10194 9560
rect 10138 9480 10194 9489
rect 10138 9415 10194 9424
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10152 8634 10180 9415
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10060 7177 10088 8570
rect 10138 8392 10194 8401
rect 10138 8327 10194 8336
rect 10244 8344 10272 10066
rect 10336 10062 10364 11086
rect 10612 11064 10640 13942
rect 10690 13832 10746 13841
rect 10690 13767 10746 13776
rect 10428 11036 10640 11064
rect 10428 10441 10456 11036
rect 10506 10976 10562 10985
rect 10704 10962 10732 13767
rect 11164 13734 11192 15438
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 11152 13524 11204 13530
rect 10796 13484 11152 13512
rect 10796 13190 10824 13484
rect 11152 13466 11204 13472
rect 10888 13348 11100 13376
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10888 12850 10916 13348
rect 10966 13288 11022 13297
rect 11072 13258 11100 13348
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10966 13223 11022 13232
rect 11060 13252 11112 13258
rect 10980 12986 11008 13223
rect 11060 13194 11112 13200
rect 11058 13152 11114 13161
rect 11058 13087 11114 13096
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 11072 12753 11100 13087
rect 11164 12782 11192 13262
rect 11152 12776 11204 12782
rect 11058 12744 11114 12753
rect 11152 12718 11204 12724
rect 11058 12679 11114 12688
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 11164 12374 11192 12718
rect 11256 12714 11284 15982
rect 11348 15502 11376 17614
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11440 16794 11468 17478
rect 11518 17232 11574 17241
rect 11518 17167 11574 17176
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11440 16289 11468 16730
rect 11426 16280 11482 16289
rect 11426 16215 11482 16224
rect 11532 15910 11560 17167
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11440 15042 11468 15506
rect 11518 15056 11574 15065
rect 11348 14414 11376 15030
rect 11440 15014 11518 15042
rect 11518 14991 11520 15000
rect 11572 14991 11574 15000
rect 11520 14962 11572 14968
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11334 14104 11390 14113
rect 11334 14039 11390 14048
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11152 12368 11204 12374
rect 11348 12322 11376 14039
rect 11440 13569 11468 14894
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11532 13938 11560 14826
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11426 13560 11482 13569
rect 11426 13495 11482 13504
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11152 12310 11204 12316
rect 11256 12306 11376 12322
rect 11244 12300 11376 12306
rect 11296 12294 11376 12300
rect 11244 12242 11296 12248
rect 11256 11778 11284 12242
rect 11336 12232 11388 12238
rect 11334 12200 11336 12209
rect 11388 12200 11390 12209
rect 11334 12135 11390 12144
rect 11164 11750 11284 11778
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 11164 11218 11192 11750
rect 11242 11656 11298 11665
rect 11242 11591 11298 11600
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10506 10911 10562 10920
rect 10612 10934 10732 10962
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10520 10810 10548 10911
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10612 10674 10640 10934
rect 10690 10840 10746 10849
rect 10690 10775 10746 10784
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10508 10464 10560 10470
rect 10414 10432 10470 10441
rect 10508 10406 10560 10412
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10414 10367 10470 10376
rect 10414 10296 10470 10305
rect 10414 10231 10416 10240
rect 10468 10231 10470 10240
rect 10416 10202 10468 10208
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9761 10364 9998
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10322 9616 10378 9625
rect 10322 9551 10378 9560
rect 10336 9382 10364 9551
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8498 10456 8910
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10324 8356 10376 8362
rect 10152 8242 10180 8327
rect 10244 8316 10324 8344
rect 10324 8298 10376 8304
rect 10152 8214 10364 8242
rect 10230 8120 10286 8129
rect 10336 8090 10364 8214
rect 10230 8055 10286 8064
rect 10324 8084 10376 8090
rect 10244 7324 10272 8055
rect 10324 8026 10376 8032
rect 10152 7296 10272 7324
rect 10152 7206 10180 7296
rect 10140 7200 10192 7206
rect 10046 7168 10102 7177
rect 10140 7142 10192 7148
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10046 7103 10102 7112
rect 10060 6458 10088 7103
rect 10152 6934 10180 7142
rect 10244 7002 10272 7142
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10230 6488 10286 6497
rect 10048 6452 10100 6458
rect 10230 6423 10286 6432
rect 10048 6394 10100 6400
rect 10244 5914 10272 6423
rect 10428 6390 10456 8434
rect 10520 8430 10548 10406
rect 10612 9722 10640 10406
rect 10704 10266 10732 10775
rect 10888 10674 10916 10950
rect 11164 10810 11192 11154
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10704 9654 10732 9998
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10874 9752 10930 9761
rect 11072 9722 11100 9862
rect 10874 9687 10930 9696
rect 11060 9716 11112 9722
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10888 9364 10916 9687
rect 11060 9658 11112 9664
rect 10598 9344 10654 9353
rect 10704 9336 10916 9364
rect 10704 9330 10732 9336
rect 10654 9302 10732 9330
rect 10598 9279 10654 9288
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10520 7585 10548 8026
rect 10506 7576 10562 7585
rect 10506 7511 10562 7520
rect 10612 7410 10640 8910
rect 10704 8022 10732 9114
rect 11058 9072 11114 9081
rect 11058 9007 11114 9016
rect 11164 9024 11192 10746
rect 11256 9092 11284 11591
rect 11348 11218 11376 12135
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10305 11376 10406
rect 11334 10296 11390 10305
rect 11334 10231 11390 10240
rect 11440 9625 11468 13398
rect 11518 13288 11574 13297
rect 11518 13223 11574 13232
rect 11532 12646 11560 13223
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11624 12209 11652 19200
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 15337 11744 15506
rect 11702 15328 11758 15337
rect 11702 15263 11758 15272
rect 11702 15192 11758 15201
rect 11702 15127 11758 15136
rect 11716 13802 11744 15127
rect 11808 15026 11836 16594
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 12850 11744 13330
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11610 12200 11666 12209
rect 11610 12135 11666 12144
rect 11518 12064 11574 12073
rect 11518 11999 11574 12008
rect 11532 11898 11560 11999
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11532 11529 11560 11562
rect 11518 11520 11574 11529
rect 11518 11455 11574 11464
rect 11624 11354 11652 11766
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11716 10520 11744 11562
rect 11624 10492 11744 10520
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9761 11560 10066
rect 11624 10062 11652 10492
rect 11702 10432 11758 10441
rect 11702 10367 11758 10376
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11518 9752 11574 9761
rect 11518 9687 11574 9696
rect 11520 9648 11572 9654
rect 11426 9616 11482 9625
rect 11520 9590 11572 9596
rect 11426 9551 11482 9560
rect 11428 9512 11480 9518
rect 11334 9480 11390 9489
rect 11532 9500 11560 9590
rect 11480 9472 11560 9500
rect 11428 9454 11480 9460
rect 11334 9415 11390 9424
rect 11348 9382 11376 9415
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11624 9217 11652 9998
rect 11610 9208 11666 9217
rect 11610 9143 11666 9152
rect 11256 9064 11652 9092
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10796 8430 10824 8842
rect 11072 8498 11100 9007
rect 11164 8996 11284 9024
rect 11150 8936 11206 8945
rect 11150 8871 11206 8880
rect 11164 8634 11192 8871
rect 11256 8809 11284 8996
rect 11336 8968 11388 8974
rect 11334 8936 11336 8945
rect 11520 8968 11572 8974
rect 11388 8936 11390 8945
rect 11334 8871 11390 8880
rect 11440 8928 11520 8956
rect 11242 8800 11298 8809
rect 11242 8735 11298 8744
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11440 8514 11468 8928
rect 11520 8910 11572 8916
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11348 8486 11468 8514
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11256 8265 11284 8298
rect 11242 8256 11298 8265
rect 10817 8188 11113 8208
rect 11242 8191 11298 8200
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 11242 8120 11298 8129
rect 11242 8055 11244 8064
rect 11296 8055 11298 8064
rect 11244 8026 11296 8032
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10704 7290 10732 7822
rect 10888 7546 10916 7890
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10980 7410 11008 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10520 7262 10732 7290
rect 10520 7177 10548 7262
rect 10796 7188 10824 7346
rect 11164 7274 11192 7346
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 10506 7168 10562 7177
rect 10506 7103 10562 7112
rect 10612 7160 10824 7188
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10140 5364 10192 5370
rect 10060 5324 10140 5352
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9862 4992 9918 5001
rect 9862 4927 9918 4936
rect 9680 4820 9732 4826
rect 9784 4814 9904 4842
rect 9680 4762 9732 4768
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9494 4448 9550 4457
rect 9494 4383 9550 4392
rect 9494 4312 9550 4321
rect 9692 4282 9720 4490
rect 9494 4247 9550 4256
rect 9680 4276 9732 4282
rect 9508 4010 9536 4247
rect 9680 4218 9732 4224
rect 9678 4176 9734 4185
rect 9678 4111 9680 4120
rect 9732 4111 9734 4120
rect 9680 4082 9732 4088
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 2650 9168 3470
rect 9232 3233 9260 3590
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9218 3224 9274 3233
rect 9274 3182 9352 3210
rect 9416 3194 9444 3538
rect 9218 3159 9274 3168
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9232 2446 9260 2994
rect 9324 2514 9352 3182
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9678 2952 9734 2961
rect 9678 2887 9734 2896
rect 9404 2576 9456 2582
rect 9692 2553 9720 2887
rect 9404 2518 9456 2524
rect 9678 2544 9734 2553
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9416 2292 9444 2518
rect 9678 2479 9734 2488
rect 9784 2417 9812 4626
rect 9876 4570 9904 4814
rect 9968 4672 9996 5238
rect 10060 4842 10088 5324
rect 10140 5306 10192 5312
rect 10230 5264 10286 5273
rect 10140 5228 10192 5234
rect 10230 5199 10286 5208
rect 10140 5170 10192 5176
rect 10152 5001 10180 5170
rect 10244 5098 10272 5199
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10138 4992 10194 5001
rect 10138 4927 10194 4936
rect 10060 4814 10272 4842
rect 9968 4644 10088 4672
rect 9876 4542 9996 4570
rect 9862 4312 9918 4321
rect 9862 4247 9864 4256
rect 9916 4247 9918 4256
rect 9864 4218 9916 4224
rect 9968 3738 9996 4542
rect 10060 3942 10088 4644
rect 10138 4176 10194 4185
rect 10244 4146 10272 4814
rect 10138 4111 10194 4120
rect 10232 4140 10284 4146
rect 10152 3942 10180 4111
rect 10232 4082 10284 4088
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9876 2496 9904 3674
rect 10060 3466 10088 3878
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10060 2854 10088 3130
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10048 2848 10100 2854
rect 10152 2825 10180 3062
rect 10244 3058 10272 4082
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10048 2790 10100 2796
rect 10138 2816 10194 2825
rect 10138 2751 10194 2760
rect 10138 2680 10194 2689
rect 10138 2615 10140 2624
rect 10192 2615 10194 2624
rect 10140 2586 10192 2592
rect 9876 2468 9996 2496
rect 9770 2408 9826 2417
rect 9968 2378 9996 2468
rect 10336 2446 10364 6190
rect 10520 6089 10548 6938
rect 10506 6080 10562 6089
rect 10506 6015 10562 6024
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10428 4282 10456 5510
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4865 10548 4966
rect 10506 4856 10562 4865
rect 10506 4791 10562 4800
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10506 4176 10562 4185
rect 10506 4111 10562 4120
rect 10520 3913 10548 4111
rect 10506 3904 10562 3913
rect 10506 3839 10562 3848
rect 10612 3754 10640 7160
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 11256 6984 11284 7890
rect 11348 7721 11376 8486
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11334 7712 11390 7721
rect 11334 7647 11390 7656
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11072 6956 11284 6984
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 11072 6882 11100 6956
rect 10796 6186 10824 6870
rect 11072 6854 11192 6882
rect 10874 6624 10930 6633
rect 10874 6559 10930 6568
rect 11058 6624 11114 6633
rect 11058 6559 11114 6568
rect 10888 6254 10916 6559
rect 10968 6452 11020 6458
rect 11072 6440 11100 6559
rect 11020 6412 11100 6440
rect 10968 6394 11020 6400
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 11164 5896 11192 6854
rect 11348 6662 11376 7482
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11440 6497 11468 8298
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11624 7970 11652 9064
rect 11716 8072 11744 10367
rect 11808 9761 11836 14554
rect 11900 11626 11928 17070
rect 11992 13297 12020 19200
rect 12072 17944 12124 17950
rect 12072 17886 12124 17892
rect 12084 16794 12112 17886
rect 12360 17377 12388 19200
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12346 17368 12402 17377
rect 12346 17303 12402 17312
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12084 15745 12112 16594
rect 12070 15736 12126 15745
rect 12070 15671 12126 15680
rect 12070 15600 12126 15609
rect 12070 15535 12126 15544
rect 12164 15564 12216 15570
rect 12084 15434 12112 15535
rect 12164 15506 12216 15512
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11978 13288 12034 13297
rect 11978 13223 12034 13232
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11992 12730 12020 13126
rect 12084 12850 12112 14962
rect 12176 13569 12204 15506
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12268 14482 12296 15370
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12162 13560 12218 13569
rect 12268 13530 12296 14418
rect 12360 13977 12388 16594
rect 12452 16046 12480 17546
rect 12532 17128 12584 17134
rect 12530 17096 12532 17105
rect 12584 17096 12586 17105
rect 12530 17031 12586 17040
rect 12636 16266 12664 19200
rect 12898 17640 12954 17649
rect 12898 17575 12954 17584
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16794 12848 17138
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12544 16238 12664 16266
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12346 13968 12402 13977
rect 12346 13903 12402 13912
rect 12452 13841 12480 15982
rect 12438 13832 12494 13841
rect 12438 13767 12494 13776
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12438 13696 12494 13705
rect 12162 13495 12218 13504
rect 12256 13524 12308 13530
rect 12176 12850 12204 13495
rect 12256 13466 12308 13472
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 11992 12702 12112 12730
rect 11978 12472 12034 12481
rect 12084 12442 12112 12702
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 11978 12407 12034 12416
rect 12072 12436 12124 12442
rect 11992 12306 12020 12407
rect 12072 12378 12124 12384
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11794 9752 11850 9761
rect 11900 9738 11928 11290
rect 11992 11257 12020 12242
rect 12176 11937 12204 12650
rect 12162 11928 12218 11937
rect 12162 11863 12218 11872
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12084 11665 12112 11766
rect 12070 11656 12126 11665
rect 12070 11591 12126 11600
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12176 11370 12204 11562
rect 12084 11342 12204 11370
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 12084 11098 12112 11342
rect 12164 11280 12216 11286
rect 12162 11248 12164 11257
rect 12216 11248 12218 11257
rect 12162 11183 12218 11192
rect 11980 11076 12032 11082
rect 12084 11070 12204 11098
rect 11980 11018 12032 11024
rect 11992 9926 12020 11018
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10266 12112 10950
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11900 9710 12020 9738
rect 12176 9722 12204 11070
rect 11794 9687 11850 9696
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11808 8566 11836 9522
rect 11900 9178 11928 9522
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11992 9092 12020 9710
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12176 9625 12204 9658
rect 12162 9616 12218 9625
rect 12162 9551 12218 9560
rect 12162 9208 12218 9217
rect 12162 9143 12218 9152
rect 11886 9072 11942 9081
rect 11992 9064 12112 9092
rect 11886 9007 11942 9016
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11808 8401 11836 8502
rect 11900 8498 11928 9007
rect 12084 8956 12112 9064
rect 12176 9042 12204 9143
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 11992 8928 12112 8956
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11794 8392 11850 8401
rect 11794 8327 11850 8336
rect 11716 8044 11928 8072
rect 11532 6780 11560 7958
rect 11624 7942 11836 7970
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11624 7721 11652 7822
rect 11610 7712 11666 7721
rect 11610 7647 11666 7656
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 6934 11744 7142
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11612 6792 11664 6798
rect 11532 6752 11612 6780
rect 11612 6734 11664 6740
rect 11426 6488 11482 6497
rect 11426 6423 11482 6432
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11334 6080 11390 6089
rect 11072 5868 11192 5896
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10888 5370 10916 5578
rect 10980 5409 11008 5646
rect 10966 5400 11022 5409
rect 10876 5364 10928 5370
rect 10966 5335 11022 5344
rect 10876 5306 10928 5312
rect 10968 5160 11020 5166
rect 11072 5148 11100 5868
rect 11256 5658 11284 6054
rect 11334 6015 11390 6024
rect 11348 5846 11376 6015
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11624 5710 11652 6734
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11164 5630 11284 5658
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11716 5642 11744 6258
rect 11704 5636 11756 5642
rect 11164 5352 11192 5630
rect 11704 5578 11756 5584
rect 11244 5568 11296 5574
rect 11296 5528 11468 5556
rect 11244 5510 11296 5516
rect 11164 5324 11284 5352
rect 11150 5264 11206 5273
rect 11150 5199 11152 5208
rect 11204 5199 11206 5208
rect 11152 5170 11204 5176
rect 11020 5120 11100 5148
rect 10968 5102 11020 5108
rect 10980 5012 11008 5102
rect 10704 4984 11008 5012
rect 11152 5024 11204 5030
rect 10704 4690 10732 4984
rect 11152 4966 11204 4972
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10980 4321 11008 4626
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10690 4312 10746 4321
rect 10690 4247 10692 4256
rect 10744 4247 10746 4256
rect 10966 4312 11022 4321
rect 10966 4247 11022 4256
rect 10692 4218 10744 4224
rect 10428 3726 10640 3754
rect 10428 2650 10456 3726
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10506 3360 10562 3369
rect 10506 3295 10562 3304
rect 10520 2650 10548 3295
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 9770 2343 9826 2352
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9232 2264 9444 2292
rect 9954 2272 10010 2281
rect 9036 1284 9088 1290
rect 9036 1226 9088 1232
rect 9232 800 9260 2264
rect 9954 2207 10010 2216
rect 9588 1624 9640 1630
rect 9588 1566 9640 1572
rect 9600 800 9628 1566
rect 9968 800 9996 2207
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 10336 800 10364 2042
rect 10612 800 10640 3606
rect 10704 2446 10732 4218
rect 11072 4146 11100 4558
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 3194 10824 3538
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10888 3097 10916 3334
rect 10874 3088 10930 3097
rect 10874 3023 10930 3032
rect 11164 2854 11192 4966
rect 11256 3738 11284 5324
rect 11334 5264 11390 5273
rect 11440 5234 11468 5528
rect 11334 5199 11390 5208
rect 11428 5228 11480 5234
rect 11348 5098 11376 5199
rect 11428 5170 11480 5176
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11440 4729 11468 4762
rect 11426 4720 11482 4729
rect 11426 4655 11482 4664
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11348 3534 11376 4422
rect 11426 4312 11482 4321
rect 11426 4247 11482 4256
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11334 2952 11390 2961
rect 11334 2887 11390 2896
rect 11348 2854 11376 2887
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10796 2310 10824 2518
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 10874 2408 10930 2417
rect 10874 2343 10930 2352
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10888 2106 10916 2343
rect 11348 2281 11376 2450
rect 11334 2272 11390 2281
rect 11334 2207 11390 2216
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 10980 800 11008 2042
rect 11348 1630 11376 2207
rect 11336 1624 11388 1630
rect 11336 1566 11388 1572
rect 11440 1442 11468 4247
rect 11624 3058 11652 5102
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11716 2922 11744 3878
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11612 1760 11664 1766
rect 11808 1748 11836 7942
rect 11900 2106 11928 8044
rect 11992 2854 12020 8928
rect 12164 8900 12216 8906
rect 12084 8860 12164 8888
rect 12084 8401 12112 8860
rect 12164 8842 12216 8848
rect 12162 8800 12218 8809
rect 12162 8735 12218 8744
rect 12070 8392 12126 8401
rect 12070 8327 12126 8336
rect 12176 7954 12204 8735
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12070 7440 12126 7449
rect 12070 7375 12126 7384
rect 12084 3942 12112 7375
rect 12176 6934 12204 7890
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12176 5778 12204 6870
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12176 4690 12204 5714
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11978 2680 12034 2689
rect 12084 2650 12112 3334
rect 11978 2615 12034 2624
rect 12072 2644 12124 2650
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 11992 1902 12020 2615
rect 12072 2586 12124 2592
rect 12176 2582 12204 4082
rect 12268 2961 12296 13330
rect 12360 13161 12388 13670
rect 12438 13631 12494 13640
rect 12452 13394 12480 13631
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12360 12442 12388 12854
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12452 12220 12480 13194
rect 12544 13025 12572 16238
rect 12624 16176 12676 16182
rect 12622 16144 12624 16153
rect 12676 16144 12678 16153
rect 12622 16079 12678 16088
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 14958 12664 15302
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12530 13016 12586 13025
rect 12530 12951 12586 12960
rect 12530 12472 12586 12481
rect 12530 12407 12586 12416
rect 12636 12424 12664 14758
rect 12728 14618 12756 16594
rect 12912 16130 12940 17575
rect 12820 16102 12940 16130
rect 12820 15094 12848 16102
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12820 14521 12848 14894
rect 12806 14512 12862 14521
rect 12806 14447 12808 14456
rect 12860 14447 12862 14456
rect 12808 14418 12860 14424
rect 12820 14387 12848 14418
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13326 12756 13806
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12728 12850 12756 13262
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12820 12617 12848 14282
rect 12806 12608 12862 12617
rect 12806 12543 12862 12552
rect 12544 12322 12572 12407
rect 12636 12396 12848 12424
rect 12544 12294 12756 12322
rect 12532 12232 12584 12238
rect 12452 12192 12532 12220
rect 12532 12174 12584 12180
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12438 12064 12494 12073
rect 12360 11354 12388 12038
rect 12438 11999 12494 12008
rect 12452 11694 12480 11999
rect 12728 11914 12756 12294
rect 12544 11886 12756 11914
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12544 11354 12572 11886
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12360 11218 12388 11290
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12636 11150 12664 11698
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12728 11354 12756 11494
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12440 11144 12492 11150
rect 12346 11112 12402 11121
rect 12440 11086 12492 11092
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12346 11047 12348 11056
rect 12400 11047 12402 11056
rect 12348 11018 12400 11024
rect 12452 10810 12480 11086
rect 12440 10804 12492 10810
rect 12360 10764 12440 10792
rect 12360 9761 12388 10764
rect 12440 10746 12492 10752
rect 12636 10538 12664 11086
rect 12728 10674 12756 11154
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 12452 10266 12480 10367
rect 12440 10260 12492 10266
rect 12820 10248 12848 12396
rect 12912 11506 12940 15982
rect 13004 14482 13032 19200
rect 13372 17524 13400 19200
rect 13188 17496 13400 17524
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12990 14376 13046 14385
rect 12990 14311 12992 14320
rect 13044 14311 13046 14320
rect 12992 14282 13044 14288
rect 13096 13462 13124 15506
rect 13188 15026 13216 17496
rect 13282 17436 13578 17456
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13556 16794 13584 17002
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13082 13152 13138 13161
rect 13082 13087 13138 13096
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 13004 11626 13032 12922
rect 13096 12628 13124 13087
rect 13188 12782 13216 14214
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13648 13802 13676 15574
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13740 13530 13768 19200
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13280 13433 13308 13466
rect 13266 13424 13322 13433
rect 13266 13359 13322 13368
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13096 12600 13216 12628
rect 13082 12472 13138 12481
rect 13082 12407 13138 12416
rect 13096 12102 13124 12407
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13084 11824 13136 11830
rect 13082 11792 13084 11801
rect 13136 11792 13138 11801
rect 13082 11727 13138 11736
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12912 11478 13032 11506
rect 13004 10810 13032 11478
rect 13096 10849 13124 11562
rect 13082 10840 13138 10849
rect 12992 10804 13044 10810
rect 13082 10775 13138 10784
rect 12992 10746 13044 10752
rect 12440 10202 12492 10208
rect 12636 10220 12848 10248
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12346 9752 12402 9761
rect 12346 9687 12402 9696
rect 12452 9586 12480 9998
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12544 9382 12572 9998
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12636 9194 12664 10220
rect 13004 10169 13032 10746
rect 13082 10568 13138 10577
rect 13082 10503 13138 10512
rect 12714 10160 12770 10169
rect 12714 10095 12770 10104
rect 12990 10160 13046 10169
rect 12990 10095 13046 10104
rect 12452 9166 12664 9194
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12360 8945 12388 8978
rect 12346 8936 12402 8945
rect 12346 8871 12402 8880
rect 12348 8832 12400 8838
rect 12346 8800 12348 8809
rect 12400 8800 12402 8809
rect 12346 8735 12402 8744
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12360 7274 12388 8434
rect 12452 8265 12480 9166
rect 12622 9072 12678 9081
rect 12622 9007 12678 9016
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12438 8256 12494 8265
rect 12438 8191 12494 8200
rect 12544 8090 12572 8910
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12636 8022 12664 9007
rect 12728 8786 12756 10095
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12820 9092 12848 9998
rect 12992 9920 13044 9926
rect 12990 9888 12992 9897
rect 13044 9888 13046 9897
rect 12990 9823 13046 9832
rect 12898 9752 12954 9761
rect 12898 9687 12954 9696
rect 12912 9217 12940 9687
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12898 9208 12954 9217
rect 12898 9143 12954 9152
rect 12820 9081 12940 9092
rect 12820 9072 12954 9081
rect 12820 9064 12898 9072
rect 12898 9007 12954 9016
rect 12728 8758 12848 8786
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12624 8016 12676 8022
rect 12438 7984 12494 7993
rect 12624 7958 12676 7964
rect 12438 7919 12494 7928
rect 12452 7546 12480 7919
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12728 7478 12756 8230
rect 12820 8090 12848 8758
rect 12912 8673 12940 9007
rect 13004 8974 13032 9522
rect 13096 9382 13124 10503
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12898 8664 12954 8673
rect 13004 8634 13032 8910
rect 13084 8832 13136 8838
rect 13082 8800 13084 8809
rect 13136 8800 13138 8809
rect 13082 8735 13138 8744
rect 12898 8599 12954 8608
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12912 8401 12940 8434
rect 13188 8430 13216 12600
rect 13266 12608 13322 12617
rect 13266 12543 13322 12552
rect 13280 12442 13308 12543
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13740 12322 13768 13330
rect 13832 13326 13860 13874
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13924 12986 13952 15982
rect 14016 14929 14044 19200
rect 14384 15473 14412 19200
rect 14370 15464 14426 15473
rect 14370 15399 14426 15408
rect 14002 14920 14058 14929
rect 14002 14855 14058 14864
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12753 13860 12786
rect 13912 12776 13964 12782
rect 13818 12744 13874 12753
rect 13912 12718 13964 12724
rect 13818 12679 13874 12688
rect 13636 12300 13688 12306
rect 13740 12294 13860 12322
rect 13636 12242 13688 12248
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13280 11121 13308 11698
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13266 11112 13322 11121
rect 13464 11098 13492 11630
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 11234 13584 11494
rect 13648 11354 13676 12242
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13556 11206 13676 11234
rect 13544 11144 13596 11150
rect 13542 11112 13544 11121
rect 13596 11112 13598 11121
rect 13464 11070 13542 11098
rect 13266 11047 13322 11056
rect 13542 11047 13598 11056
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13544 10736 13596 10742
rect 13450 10704 13506 10713
rect 13268 10668 13320 10674
rect 13544 10678 13596 10684
rect 13450 10639 13452 10648
rect 13268 10610 13320 10616
rect 13504 10639 13506 10648
rect 13452 10610 13504 10616
rect 13280 10198 13308 10610
rect 13556 10470 13584 10678
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13464 10266 13492 10406
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13648 9994 13676 11206
rect 13740 10810 13768 12174
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 10062 13768 10542
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13740 9081 13768 9522
rect 13832 9382 13860 12294
rect 13924 11642 13952 12718
rect 14016 11830 14044 14855
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 13924 11614 14044 11642
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13726 9072 13782 9081
rect 13636 9036 13688 9042
rect 13726 9007 13782 9016
rect 13636 8978 13688 8984
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13648 8634 13676 8978
rect 13740 8974 13768 9007
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13832 8514 13860 9318
rect 13924 9110 13952 11494
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13648 8486 13860 8514
rect 13176 8424 13228 8430
rect 12898 8392 12954 8401
rect 12898 8327 12954 8336
rect 13096 8384 13176 8412
rect 12990 8120 13046 8129
rect 12808 8084 12860 8090
rect 12990 8055 13046 8064
rect 12808 8026 12860 8032
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12452 6866 12480 7278
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 12346 6624 12402 6633
rect 12346 6559 12402 6568
rect 12360 6168 12388 6559
rect 12452 6338 12480 6695
rect 12544 6458 12572 6938
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12452 6310 12572 6338
rect 12360 6140 12480 6168
rect 12346 6080 12402 6089
rect 12346 6015 12402 6024
rect 12360 5914 12388 6015
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 5370 12388 5510
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5098 12480 6140
rect 12544 6066 12572 6310
rect 12636 6186 12664 6802
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12544 6038 12664 6066
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12346 4992 12402 5001
rect 12346 4927 12402 4936
rect 12360 4758 12388 4927
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12254 2952 12310 2961
rect 12254 2887 12310 2896
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12176 2038 12204 2246
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 11980 1896 12032 1902
rect 11980 1838 12032 1844
rect 12256 1896 12308 1902
rect 12256 1838 12308 1844
rect 11808 1720 12020 1748
rect 11612 1702 11664 1708
rect 11348 1414 11468 1442
rect 11348 800 11376 1414
rect 11624 800 11652 1702
rect 11992 800 12020 1720
rect 12268 1442 12296 1838
rect 12360 1766 12388 4694
rect 12544 4570 12572 5714
rect 12636 5302 12664 6038
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12452 4542 12572 4570
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12452 3194 12480 4542
rect 12636 4486 12664 4558
rect 12624 4480 12676 4486
rect 12530 4448 12586 4457
rect 12624 4422 12676 4428
rect 12530 4383 12586 4392
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 2990 12572 4383
rect 12728 3670 12756 7210
rect 12820 7002 12848 7754
rect 12912 7410 12940 7890
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13004 7206 13032 8055
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 13096 6934 13124 8384
rect 13176 8366 13228 8372
rect 13280 7886 13308 8434
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7410 13216 7686
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13648 7528 13676 8486
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13740 8090 13768 8298
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13556 7500 13676 7528
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13084 6928 13136 6934
rect 12806 6896 12862 6905
rect 13084 6870 13136 6876
rect 12806 6831 12862 6840
rect 12820 5914 12848 6831
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 6186 12940 6598
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 13004 6118 13032 6734
rect 13188 6610 13216 7210
rect 13280 6730 13308 7414
rect 13556 7274 13584 7500
rect 13634 7304 13690 7313
rect 13544 7268 13596 7274
rect 13634 7239 13690 7248
rect 13544 7210 13596 7216
rect 13648 7206 13676 7239
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13634 7032 13690 7041
rect 13634 6967 13690 6976
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13096 6582 13216 6610
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12820 4826 12848 5714
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12806 4312 12862 4321
rect 12806 4247 12862 4256
rect 12820 3942 12848 4247
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12452 2650 12480 2926
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12544 1834 12572 2450
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12622 2136 12678 2145
rect 12622 2071 12678 2080
rect 12532 1828 12584 1834
rect 12532 1770 12584 1776
rect 12348 1760 12400 1766
rect 12348 1702 12400 1708
rect 12268 1414 12388 1442
rect 12360 800 12388 1414
rect 12636 800 12664 2071
rect 12728 1902 12756 2382
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 12820 1698 12848 3538
rect 12912 3233 12940 5782
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 5409 13032 5714
rect 12990 5400 13046 5409
rect 12990 5335 13046 5344
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 13004 4622 13032 5034
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13004 4146 13032 4558
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3738 13032 3878
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13096 3618 13124 6582
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5370 13216 6054
rect 13280 5953 13308 6122
rect 13266 5944 13322 5953
rect 13266 5879 13322 5888
rect 13372 5710 13400 6258
rect 13452 6112 13504 6118
rect 13450 6080 13452 6089
rect 13504 6080 13506 6089
rect 13450 6015 13506 6024
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13188 4282 13216 5170
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13556 4758 13584 5034
rect 13648 4826 13676 6967
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 6390 13768 6666
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13740 5914 13768 6190
rect 13832 6118 13860 8230
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13832 5681 13860 6054
rect 13818 5672 13874 5681
rect 13818 5607 13874 5616
rect 13832 5302 13860 5607
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13726 4856 13782 4865
rect 13636 4820 13688 4826
rect 13726 4791 13782 4800
rect 13636 4762 13688 4768
rect 13740 4758 13768 4791
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13004 3590 13124 3618
rect 13280 3602 13308 4014
rect 13544 4004 13596 4010
rect 13740 3992 13768 4694
rect 13924 4162 13952 8774
rect 14016 7546 14044 11614
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 7002 14044 7142
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14016 5914 14044 6802
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14002 5536 14058 5545
rect 14002 5471 14058 5480
rect 14016 4978 14044 5471
rect 14108 5166 14136 14350
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14200 12782 14228 13806
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14200 11257 14228 12242
rect 14186 11248 14242 11257
rect 14186 11183 14242 11192
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14200 10674 14228 11086
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10033 14228 10406
rect 14186 10024 14242 10033
rect 14186 9959 14242 9968
rect 14292 9466 14320 14418
rect 14384 13258 14412 15399
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14476 13530 14504 14826
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14568 12968 14596 14962
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14384 12940 14596 12968
rect 14384 10305 14412 12940
rect 14554 12880 14610 12889
rect 14554 12815 14610 12824
rect 14568 12782 14596 12815
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14476 11218 14504 11766
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14370 10296 14426 10305
rect 14370 10231 14426 10240
rect 14384 10130 14412 10231
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14200 9450 14320 9466
rect 14188 9444 14320 9450
rect 14240 9438 14320 9444
rect 14188 9386 14240 9392
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14200 7410 14228 7822
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14200 5817 14228 7142
rect 14186 5808 14242 5817
rect 14186 5743 14242 5752
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14096 5024 14148 5030
rect 14016 4972 14096 4978
rect 14016 4966 14148 4972
rect 14016 4950 14136 4966
rect 13544 3946 13596 3952
rect 13648 3964 13768 3992
rect 13832 4134 13952 4162
rect 13556 3670 13584 3946
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13268 3596 13320 3602
rect 12898 3224 12954 3233
rect 12898 3159 12954 3168
rect 12808 1692 12860 1698
rect 12808 1634 12860 1640
rect 13004 800 13032 3590
rect 13268 3538 13320 3544
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13544 3052 13596 3058
rect 13648 3040 13676 3964
rect 13726 3904 13782 3913
rect 13726 3839 13782 3848
rect 13596 3012 13676 3040
rect 13544 2994 13596 3000
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13360 2032 13412 2038
rect 13360 1974 13412 1980
rect 13372 800 13400 1974
rect 13740 800 13768 3839
rect 13832 2825 13860 4134
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13924 3641 13952 3946
rect 13910 3632 13966 3641
rect 13910 3567 13966 3576
rect 13818 2816 13874 2825
rect 13818 2751 13874 2760
rect 14016 2514 14044 4014
rect 14108 3942 14136 4950
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14016 800 14044 2450
rect 14200 2038 14228 4762
rect 14292 4185 14320 9318
rect 14278 4176 14334 4185
rect 14278 4111 14334 4120
rect 14384 3505 14412 9862
rect 14476 9722 14504 11154
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14462 9208 14518 9217
rect 14462 9143 14518 9152
rect 14476 9042 14504 9143
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14464 8560 14516 8566
rect 14462 8528 14464 8537
rect 14516 8528 14518 8537
rect 14462 8463 14518 8472
rect 14568 8430 14596 11222
rect 14660 9518 14688 13194
rect 14752 11694 14780 19200
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14476 6798 14504 7754
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14476 3738 14504 6258
rect 14568 5098 14596 8366
rect 14752 7954 14780 10678
rect 14844 10033 14872 12650
rect 14830 10024 14886 10033
rect 14830 9959 14886 9968
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 6361 14688 7686
rect 14646 6352 14702 6361
rect 14646 6287 14702 6296
rect 14556 5092 14608 5098
rect 14556 5034 14608 5040
rect 14752 4622 14780 7890
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 4616 14792 4622
rect 14646 4584 14702 4593
rect 14740 4558 14792 4564
rect 14646 4519 14648 4528
rect 14700 4519 14702 4528
rect 14648 4490 14700 4496
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14556 4072 14608 4078
rect 14752 4049 14780 4082
rect 14556 4014 14608 4020
rect 14738 4040 14794 4049
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14568 3602 14596 4014
rect 14844 4026 14872 7482
rect 14936 4146 14964 13806
rect 15028 12306 15056 19200
rect 15396 15434 15424 19200
rect 15764 16561 15792 19200
rect 16040 17542 16068 19200
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15750 16552 15806 16561
rect 15750 16487 15806 16496
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 16408 15065 16436 19200
rect 16776 15366 16804 19200
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16394 15056 16450 15065
rect 16394 14991 16450 15000
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15014 12200 15070 12209
rect 15014 12135 15070 12144
rect 15028 7342 15056 12135
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15028 6322 15056 7278
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15014 6216 15070 6225
rect 15014 6151 15070 6160
rect 15028 6118 15056 6151
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15014 5128 15070 5137
rect 15014 5063 15070 5072
rect 15028 5030 15056 5063
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14844 3998 15056 4026
rect 14738 3975 14794 3984
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14370 3496 14426 3505
rect 14370 3431 14426 3440
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14384 2650 14412 2926
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14188 2032 14240 2038
rect 14188 1974 14240 1980
rect 14384 800 14412 2586
rect 14752 800 14780 3538
rect 15028 800 15056 3998
rect 15120 3369 15148 11698
rect 15304 10606 15332 13398
rect 15292 10600 15344 10606
rect 15212 10560 15292 10588
rect 15212 8265 15240 10560
rect 15292 10542 15344 10548
rect 15198 8256 15254 8265
rect 15198 8191 15254 8200
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 15106 3360 15162 3369
rect 15106 3295 15162 3304
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15396 800 15424 2382
rect 15764 800 15792 2858
rect 16040 800 16068 2994
rect 16408 800 16436 3470
rect 16776 800 16804 4082
rect 2870 504 2926 513
rect 2870 439 2926 448
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
<< via2 >>
rect 2962 19352 3018 19408
rect 1398 11328 1454 11384
rect 1306 6432 1362 6488
rect 1122 6160 1178 6216
rect 754 5072 810 5128
rect 386 4664 442 4720
rect 1398 4392 1454 4448
rect 1858 14320 1914 14376
rect 2042 13524 2098 13560
rect 2042 13504 2044 13524
rect 2044 13504 2096 13524
rect 2096 13504 2098 13524
rect 2042 12300 2098 12336
rect 2042 12280 2044 12300
rect 2044 12280 2096 12300
rect 2096 12280 2098 12300
rect 2778 18536 2834 18592
rect 2778 18400 2834 18456
rect 1858 10376 1914 10432
rect 1674 7384 1730 7440
rect 1674 6296 1730 6352
rect 1582 5616 1638 5672
rect 1490 2760 1546 2816
rect 1398 2352 1454 2408
rect 2410 14320 2466 14376
rect 2962 15408 3018 15464
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 3882 17060 3938 17096
rect 3882 17040 3884 17060
rect 3884 17040 3936 17060
rect 3936 17040 3938 17060
rect 2318 10532 2374 10568
rect 2318 10512 2320 10532
rect 2320 10512 2372 10532
rect 2372 10512 2374 10532
rect 1950 7928 2006 7984
rect 1858 6976 1914 7032
rect 1950 4800 2006 4856
rect 2134 4256 2190 4312
rect 2042 3732 2098 3768
rect 2042 3712 2044 3732
rect 2044 3712 2096 3732
rect 2096 3712 2098 3732
rect 1858 1400 1914 1456
rect 2686 12688 2742 12744
rect 3238 16360 3294 16416
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 2962 13368 3018 13424
rect 2870 12416 2926 12472
rect 2410 2896 2466 2952
rect 3146 11620 3202 11656
rect 3146 11600 3148 11620
rect 3148 11600 3200 11620
rect 3200 11600 3202 11620
rect 3146 10648 3202 10704
rect 3146 10124 3202 10160
rect 3146 10104 3148 10124
rect 3148 10104 3200 10124
rect 3200 10104 3202 10124
rect 3054 9424 3110 9480
rect 2594 4936 2650 4992
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3514 9444 3570 9480
rect 3514 9424 3516 9444
rect 3516 9424 3568 9444
rect 3568 9424 3570 9444
rect 4342 15988 4344 16008
rect 4344 15988 4396 16008
rect 4396 15988 4398 16008
rect 4342 15952 4398 15988
rect 4066 14456 4122 14512
rect 4250 13776 4306 13832
rect 4250 12980 4306 13016
rect 4250 12960 4252 12980
rect 4252 12960 4304 12980
rect 4304 12960 4306 12980
rect 3974 11736 4030 11792
rect 3974 11464 4030 11520
rect 3882 9968 3938 10024
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3238 8336 3294 8392
rect 3882 8336 3938 8392
rect 3330 8200 3386 8256
rect 3238 7248 3294 7304
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3790 6840 3846 6896
rect 3238 6740 3240 6760
rect 3240 6740 3292 6760
rect 3292 6740 3294 6760
rect 3238 6704 3294 6740
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 2686 3576 2742 3632
rect 2778 3032 2834 3088
rect 3054 4684 3110 4720
rect 3054 4664 3056 4684
rect 3056 4664 3108 4684
rect 3108 4664 3110 4684
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3606 4936 3662 4992
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3330 3848 3386 3904
rect 3146 3440 3202 3496
rect 3330 3440 3386 3496
rect 4066 9560 4122 9616
rect 4342 11872 4398 11928
rect 4158 9152 4214 9208
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 4802 14864 4858 14920
rect 5630 15000 5686 15056
rect 5262 13912 5318 13968
rect 4710 13232 4766 13288
rect 4802 12860 4804 12880
rect 4804 12860 4856 12880
rect 4856 12860 4858 12880
rect 4802 12824 4858 12860
rect 5078 12824 5134 12880
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 6550 16088 6606 16144
rect 6274 14728 6330 14784
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5998 14320 6054 14376
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5906 12960 5962 13016
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5170 12144 5226 12200
rect 4618 11228 4620 11248
rect 4620 11228 4672 11248
rect 4672 11228 4674 11248
rect 4618 11192 4674 11228
rect 5354 11872 5410 11928
rect 4526 9016 4582 9072
rect 4342 8744 4398 8800
rect 4066 6432 4122 6488
rect 3882 4256 3938 4312
rect 3882 3304 3938 3360
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 4250 5344 4306 5400
rect 4158 4936 4214 4992
rect 4250 4800 4306 4856
rect 4066 4120 4122 4176
rect 4250 4140 4306 4176
rect 4250 4120 4252 4140
rect 4252 4120 4304 4140
rect 4304 4120 4306 4140
rect 4158 3712 4214 3768
rect 4434 7792 4490 7848
rect 4434 4664 4490 4720
rect 4618 4800 4674 4856
rect 5078 8472 5134 8528
rect 4802 7384 4858 7440
rect 4894 6976 4950 7032
rect 4802 4664 4858 4720
rect 5078 6568 5134 6624
rect 5078 5752 5134 5808
rect 5446 10648 5502 10704
rect 5630 9152 5686 9208
rect 5538 8880 5594 8936
rect 5538 8236 5540 8256
rect 5540 8236 5592 8256
rect 5592 8236 5594 8256
rect 5538 8200 5594 8236
rect 5354 6840 5410 6896
rect 5262 5480 5318 5536
rect 5262 4684 5318 4720
rect 5262 4664 5264 4684
rect 5264 4664 5316 4684
rect 5316 4664 5318 4684
rect 5262 4392 5318 4448
rect 5170 3848 5226 3904
rect 4434 3032 4490 3088
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 3514 1944 3570 2000
rect 5538 6876 5540 6896
rect 5540 6876 5592 6896
rect 5592 6876 5594 6896
rect 5538 6840 5594 6876
rect 5538 4936 5594 4992
rect 5722 4664 5778 4720
rect 5722 4392 5778 4448
rect 6458 14592 6514 14648
rect 7010 15544 7066 15600
rect 6826 14864 6882 14920
rect 6642 14456 6698 14512
rect 7194 16496 7250 16552
rect 7378 15852 7380 15872
rect 7380 15852 7432 15872
rect 7432 15852 7434 15872
rect 7378 15816 7434 15852
rect 7194 15408 7250 15464
rect 6642 13776 6698 13832
rect 6642 13368 6698 13424
rect 6550 12824 6606 12880
rect 7102 14320 7158 14376
rect 6734 12552 6790 12608
rect 6642 12180 6644 12200
rect 6644 12180 6696 12200
rect 6696 12180 6698 12200
rect 6642 12144 6698 12180
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 6274 8200 6330 8256
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 6182 4392 6238 4448
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 7930 17176 7986 17232
rect 8574 17584 8630 17640
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 8390 16904 8446 16960
rect 8574 16632 8630 16688
rect 8298 16496 8354 16552
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8022 15680 8078 15736
rect 7746 14184 7802 14240
rect 8022 14864 8078 14920
rect 8022 13504 8078 13560
rect 8482 15816 8538 15872
rect 8574 15408 8630 15464
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8298 14728 8354 14784
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8022 12688 8078 12744
rect 7378 12144 7434 12200
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 7930 11600 7986 11656
rect 7470 11056 7526 11112
rect 6642 7928 6698 7984
rect 6642 4820 6698 4856
rect 6642 4800 6644 4820
rect 6644 4800 6696 4820
rect 6696 4800 6698 4820
rect 7194 9424 7250 9480
rect 7194 7248 7250 7304
rect 7010 6976 7066 7032
rect 6918 4120 6974 4176
rect 7286 5752 7342 5808
rect 7286 5208 7342 5264
rect 7746 9152 7802 9208
rect 7838 8336 7894 8392
rect 7838 6568 7894 6624
rect 7470 5208 7526 5264
rect 7838 5616 7894 5672
rect 7102 3848 7158 3904
rect 7102 3168 7158 3224
rect 6918 2352 6974 2408
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 9310 16632 9366 16688
rect 8758 16360 8814 16416
rect 8850 14184 8906 14240
rect 8850 12960 8906 13016
rect 8850 12824 8906 12880
rect 8942 12144 8998 12200
rect 8850 11192 8906 11248
rect 8114 10412 8116 10432
rect 8116 10412 8168 10432
rect 8168 10412 8170 10432
rect 8114 10376 8170 10412
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8482 9560 8538 9616
rect 8022 8744 8078 8800
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8758 7656 8814 7712
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8022 6432 8078 6488
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8850 6840 8906 6896
rect 8482 6024 8538 6080
rect 8022 5244 8024 5264
rect 8024 5244 8076 5264
rect 8076 5244 8078 5264
rect 8022 5208 8078 5244
rect 8022 4936 8078 4992
rect 7930 3032 7986 3088
rect 8206 5480 8262 5536
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8758 6024 8814 6080
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 9310 15272 9366 15328
rect 9310 14864 9366 14920
rect 9034 10648 9090 10704
rect 9770 16496 9826 16552
rect 9678 15852 9680 15872
rect 9680 15852 9732 15872
rect 9732 15852 9734 15872
rect 9678 15816 9734 15852
rect 9678 15136 9734 15192
rect 9954 15680 10010 15736
rect 9862 15136 9918 15192
rect 9586 14864 9642 14920
rect 9862 14356 9864 14376
rect 9864 14356 9916 14376
rect 9916 14356 9918 14376
rect 9678 14048 9734 14104
rect 9862 14320 9918 14356
rect 9862 14184 9918 14240
rect 9770 13912 9826 13968
rect 9310 12180 9312 12200
rect 9312 12180 9364 12200
rect 9364 12180 9366 12200
rect 9310 12144 9366 12180
rect 9586 11872 9642 11928
rect 9494 10240 9550 10296
rect 9494 9696 9550 9752
rect 9310 9324 9312 9344
rect 9312 9324 9364 9344
rect 9364 9324 9366 9344
rect 9310 9288 9366 9324
rect 9126 9152 9182 9208
rect 9126 8200 9182 8256
rect 9586 9152 9642 9208
rect 10046 14592 10102 14648
rect 10322 16904 10378 16960
rect 10322 14592 10378 14648
rect 10506 15816 10562 15872
rect 10046 14320 10102 14376
rect 10046 13640 10102 13696
rect 9954 12960 10010 13016
rect 10046 12824 10102 12880
rect 9862 12416 9918 12472
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 10782 16496 10838 16552
rect 10690 16224 10746 16280
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10230 13640 10286 13696
rect 10414 14068 10470 14104
rect 10414 14048 10416 14068
rect 10416 14048 10468 14068
rect 10468 14048 10470 14068
rect 10414 13912 10470 13968
rect 10966 15000 11022 15056
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 11058 14456 11114 14512
rect 10690 14184 10746 14240
rect 10598 14048 10654 14104
rect 10138 12144 10194 12200
rect 9770 11600 9826 11656
rect 9494 8336 9550 8392
rect 9034 6024 9090 6080
rect 9126 5616 9182 5672
rect 9770 8608 9826 8664
rect 10414 12688 10470 12744
rect 10322 11328 10378 11384
rect 10046 10920 10102 10976
rect 9770 8200 9826 8256
rect 9586 7112 9642 7168
rect 9402 6976 9458 7032
rect 9862 6432 9918 6488
rect 9586 5480 9642 5536
rect 9586 5344 9642 5400
rect 10138 9560 10194 9616
rect 10138 9424 10194 9480
rect 10138 8336 10194 8392
rect 10690 13776 10746 13832
rect 10506 10920 10562 10976
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10966 13232 11022 13288
rect 11058 13096 11114 13152
rect 11058 12688 11114 12744
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 11518 17176 11574 17232
rect 11426 16224 11482 16280
rect 11518 15020 11574 15056
rect 11518 15000 11520 15020
rect 11520 15000 11572 15020
rect 11572 15000 11574 15020
rect 11334 14048 11390 14104
rect 11426 13504 11482 13560
rect 11334 12180 11336 12200
rect 11336 12180 11388 12200
rect 11388 12180 11390 12200
rect 11334 12144 11390 12180
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 11242 11600 11298 11656
rect 10690 10784 10746 10840
rect 10414 10376 10470 10432
rect 10414 10260 10470 10296
rect 10414 10240 10416 10260
rect 10416 10240 10468 10260
rect 10468 10240 10470 10260
rect 10322 9696 10378 9752
rect 10322 9560 10378 9616
rect 10230 8064 10286 8120
rect 10046 7112 10102 7168
rect 10230 6432 10286 6488
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10874 9696 10930 9752
rect 10598 9288 10654 9344
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10506 7520 10562 7576
rect 11058 9016 11114 9072
rect 11334 10240 11390 10296
rect 11518 13232 11574 13288
rect 11702 15272 11758 15328
rect 11702 15136 11758 15192
rect 11610 12144 11666 12200
rect 11518 12008 11574 12064
rect 11518 11464 11574 11520
rect 11702 10376 11758 10432
rect 11518 9696 11574 9752
rect 11426 9560 11482 9616
rect 11334 9424 11390 9480
rect 11610 9152 11666 9208
rect 11150 8880 11206 8936
rect 11334 8916 11336 8936
rect 11336 8916 11388 8936
rect 11388 8916 11390 8936
rect 11334 8880 11390 8916
rect 11242 8744 11298 8800
rect 11242 8200 11298 8256
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 11242 8084 11298 8120
rect 11242 8064 11244 8084
rect 11244 8064 11296 8084
rect 11296 8064 11298 8084
rect 10506 7112 10562 7168
rect 9862 4936 9918 4992
rect 9494 4392 9550 4448
rect 9494 4256 9550 4312
rect 9678 4140 9734 4176
rect 9678 4120 9680 4140
rect 9680 4120 9732 4140
rect 9732 4120 9734 4140
rect 9218 3168 9274 3224
rect 9678 2896 9734 2952
rect 9678 2488 9734 2544
rect 10230 5208 10286 5264
rect 10138 4936 10194 4992
rect 9862 4276 9918 4312
rect 9862 4256 9864 4276
rect 9864 4256 9916 4276
rect 9916 4256 9918 4276
rect 10138 4120 10194 4176
rect 10138 2760 10194 2816
rect 10138 2644 10194 2680
rect 10138 2624 10140 2644
rect 10140 2624 10192 2644
rect 10192 2624 10194 2644
rect 9770 2352 9826 2408
rect 10506 6024 10562 6080
rect 10506 4800 10562 4856
rect 10506 4120 10562 4176
rect 10506 3848 10562 3904
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 11334 7656 11390 7712
rect 10874 6568 10930 6624
rect 11058 6568 11114 6624
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 12346 17312 12402 17368
rect 12070 15680 12126 15736
rect 12070 15544 12126 15600
rect 11978 13232 12034 13288
rect 12162 13504 12218 13560
rect 12530 17076 12532 17096
rect 12532 17076 12584 17096
rect 12584 17076 12586 17096
rect 12530 17040 12586 17076
rect 12898 17584 12954 17640
rect 12346 13912 12402 13968
rect 12438 13776 12494 13832
rect 11978 12416 12034 12472
rect 11794 9696 11850 9752
rect 12162 11872 12218 11928
rect 12070 11600 12126 11656
rect 11978 11192 12034 11248
rect 12162 11228 12164 11248
rect 12164 11228 12216 11248
rect 12216 11228 12218 11248
rect 12162 11192 12218 11228
rect 12162 9560 12218 9616
rect 12162 9152 12218 9208
rect 11886 9016 11942 9072
rect 11794 8336 11850 8392
rect 11610 7656 11666 7712
rect 11426 6432 11482 6488
rect 10966 5344 11022 5400
rect 11334 6024 11390 6080
rect 11150 5228 11206 5264
rect 11150 5208 11152 5228
rect 11152 5208 11204 5228
rect 11204 5208 11206 5228
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10690 4276 10746 4312
rect 10690 4256 10692 4276
rect 10692 4256 10744 4276
rect 10744 4256 10746 4276
rect 10966 4256 11022 4312
rect 10506 3304 10562 3360
rect 9954 2216 10010 2272
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10874 3032 10930 3088
rect 11334 5208 11390 5264
rect 11426 4664 11482 4720
rect 11426 4256 11482 4312
rect 11334 2896 11390 2952
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 10874 2352 10930 2408
rect 11334 2216 11390 2272
rect 12162 8744 12218 8800
rect 12070 8336 12126 8392
rect 12070 7384 12126 7440
rect 11978 2624 12034 2680
rect 12438 13640 12494 13696
rect 12346 13096 12402 13152
rect 12622 16124 12624 16144
rect 12624 16124 12676 16144
rect 12676 16124 12678 16144
rect 12622 16088 12678 16124
rect 12530 12960 12586 13016
rect 12530 12416 12586 12472
rect 12806 14476 12862 14512
rect 12806 14456 12808 14476
rect 12808 14456 12860 14476
rect 12860 14456 12862 14476
rect 12806 12552 12862 12608
rect 12438 12008 12494 12064
rect 12346 11076 12402 11112
rect 12346 11056 12348 11076
rect 12348 11056 12400 11076
rect 12400 11056 12402 11076
rect 12438 10376 12494 10432
rect 12990 14340 13046 14376
rect 12990 14320 12992 14340
rect 12992 14320 13044 14340
rect 13044 14320 13046 14340
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13082 13096 13138 13152
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13266 13368 13322 13424
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13082 12416 13138 12472
rect 13082 11772 13084 11792
rect 13084 11772 13136 11792
rect 13136 11772 13138 11792
rect 13082 11736 13138 11772
rect 13082 10784 13138 10840
rect 12346 9696 12402 9752
rect 13082 10512 13138 10568
rect 12714 10104 12770 10160
rect 12990 10104 13046 10160
rect 12346 8880 12402 8936
rect 12346 8780 12348 8800
rect 12348 8780 12400 8800
rect 12400 8780 12402 8800
rect 12346 8744 12402 8780
rect 12622 9016 12678 9072
rect 12438 8200 12494 8256
rect 12990 9868 12992 9888
rect 12992 9868 13044 9888
rect 13044 9868 13046 9888
rect 12990 9832 13046 9868
rect 12898 9696 12954 9752
rect 12898 9152 12954 9208
rect 12898 9016 12954 9072
rect 12438 7928 12494 7984
rect 12898 8608 12954 8664
rect 13082 8780 13084 8800
rect 13084 8780 13136 8800
rect 13136 8780 13138 8800
rect 13082 8744 13138 8780
rect 13266 12552 13322 12608
rect 14370 15408 14426 15464
rect 14002 14864 14058 14920
rect 13818 12688 13874 12744
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13266 11056 13322 11112
rect 13542 11092 13544 11112
rect 13544 11092 13596 11112
rect 13596 11092 13598 11112
rect 13542 11056 13598 11092
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13450 10668 13506 10704
rect 13450 10648 13452 10668
rect 13452 10648 13504 10668
rect 13504 10648 13506 10668
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13726 9016 13782 9072
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 12898 8336 12954 8392
rect 12990 8064 13046 8120
rect 12438 6704 12494 6760
rect 12346 6568 12402 6624
rect 12346 6024 12402 6080
rect 12346 4936 12402 4992
rect 12254 2896 12310 2952
rect 12530 4392 12586 4448
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 12806 6840 12862 6896
rect 13634 7248 13690 7304
rect 13634 6976 13690 7032
rect 12806 4256 12862 4312
rect 12622 2080 12678 2136
rect 12990 5344 13046 5400
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13266 5888 13322 5944
rect 13450 6060 13452 6080
rect 13452 6060 13504 6080
rect 13504 6060 13506 6080
rect 13450 6024 13506 6060
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13818 5616 13874 5672
rect 13726 4800 13782 4856
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 14002 5480 14058 5536
rect 14186 11192 14242 11248
rect 14186 9968 14242 10024
rect 14554 12824 14610 12880
rect 14370 10240 14426 10296
rect 14186 5752 14242 5808
rect 12898 3168 12954 3224
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13726 3848 13782 3904
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 13910 3576 13966 3632
rect 13818 2760 13874 2816
rect 14278 4120 14334 4176
rect 14462 9152 14518 9208
rect 14462 8508 14464 8528
rect 14464 8508 14516 8528
rect 14516 8508 14518 8528
rect 14462 8472 14518 8508
rect 14830 9968 14886 10024
rect 14646 6296 14702 6352
rect 14646 4548 14702 4584
rect 14646 4528 14648 4548
rect 14648 4528 14700 4548
rect 14700 4528 14702 4548
rect 14738 3984 14794 4040
rect 15750 16496 15806 16552
rect 16394 15000 16450 15056
rect 15014 12144 15070 12200
rect 15014 6160 15070 6216
rect 15014 5072 15070 5128
rect 14370 3440 14426 3496
rect 15198 8200 15254 8256
rect 15106 3304 15162 3360
rect 2870 448 2926 504
<< metal3 >>
rect 0 19410 800 19440
rect 2957 19410 3023 19413
rect 0 19408 3023 19410
rect 0 19352 2962 19408
rect 3018 19352 3023 19408
rect 0 19350 3023 19352
rect 0 19320 800 19350
rect 2957 19347 3023 19350
rect 2773 18594 2839 18597
rect 9070 18594 9076 18596
rect 2773 18592 9076 18594
rect 2773 18536 2778 18592
rect 2834 18536 9076 18592
rect 2773 18534 9076 18536
rect 2773 18531 2839 18534
rect 9070 18532 9076 18534
rect 9140 18532 9146 18596
rect 0 18458 800 18488
rect 2773 18458 2839 18461
rect 0 18456 2839 18458
rect 0 18400 2778 18456
rect 2834 18400 2839 18456
rect 0 18398 2839 18400
rect 0 18368 800 18398
rect 2773 18395 2839 18398
rect 8569 17642 8635 17645
rect 12893 17642 12959 17645
rect 8569 17640 12959 17642
rect 8569 17584 8574 17640
rect 8630 17584 12898 17640
rect 12954 17584 12959 17640
rect 8569 17582 12959 17584
rect 8569 17579 8635 17582
rect 12893 17579 12959 17582
rect 3409 17440 3729 17441
rect 0 17280 800 17400
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 17375 13590 17376
rect 9990 17308 9996 17372
rect 10060 17370 10066 17372
rect 12341 17370 12407 17373
rect 10060 17368 12407 17370
rect 10060 17312 12346 17368
rect 12402 17312 12407 17368
rect 10060 17310 12407 17312
rect 10060 17308 10066 17310
rect 12341 17307 12407 17310
rect 7925 17234 7991 17237
rect 11513 17234 11579 17237
rect 7925 17232 11579 17234
rect 7925 17176 7930 17232
rect 7986 17176 11518 17232
rect 11574 17176 11579 17232
rect 7925 17174 11579 17176
rect 7925 17171 7991 17174
rect 11513 17171 11579 17174
rect 3877 17098 3943 17101
rect 11278 17098 11284 17100
rect 3877 17096 11284 17098
rect 3877 17040 3882 17096
rect 3938 17040 11284 17096
rect 3877 17038 11284 17040
rect 3877 17035 3943 17038
rect 11278 17036 11284 17038
rect 11348 17036 11354 17100
rect 12382 17036 12388 17100
rect 12452 17098 12458 17100
rect 12525 17098 12591 17101
rect 12452 17096 12591 17098
rect 12452 17040 12530 17096
rect 12586 17040 12591 17096
rect 12452 17038 12591 17040
rect 12452 17036 12458 17038
rect 12525 17035 12591 17038
rect 8385 16962 8451 16965
rect 10317 16962 10383 16965
rect 8385 16960 10383 16962
rect 8385 16904 8390 16960
rect 8446 16904 10322 16960
rect 10378 16904 10383 16960
rect 8385 16902 10383 16904
rect 8385 16899 8451 16902
rect 10317 16899 10383 16902
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 8569 16690 8635 16693
rect 9305 16690 9371 16693
rect 8569 16688 9371 16690
rect 8569 16632 8574 16688
rect 8630 16632 9310 16688
rect 9366 16632 9371 16688
rect 8569 16630 9371 16632
rect 8569 16627 8635 16630
rect 9305 16627 9371 16630
rect 16200 16600 17000 16720
rect 7189 16554 7255 16557
rect 8293 16554 8359 16557
rect 7189 16552 8359 16554
rect 7189 16496 7194 16552
rect 7250 16496 8298 16552
rect 8354 16496 8359 16552
rect 7189 16494 8359 16496
rect 7189 16491 7255 16494
rect 8293 16491 8359 16494
rect 9765 16556 9831 16557
rect 9765 16552 9812 16556
rect 9876 16554 9882 16556
rect 9765 16496 9770 16552
rect 9765 16492 9812 16496
rect 9876 16494 9922 16554
rect 9876 16492 9882 16494
rect 10174 16492 10180 16556
rect 10244 16554 10250 16556
rect 10777 16554 10843 16557
rect 15745 16554 15811 16557
rect 10244 16552 10843 16554
rect 10244 16496 10782 16552
rect 10838 16496 10843 16552
rect 10244 16494 10843 16496
rect 10244 16492 10250 16494
rect 9765 16491 9831 16492
rect 10777 16491 10843 16494
rect 12712 16552 15811 16554
rect 12712 16496 15750 16552
rect 15806 16496 15811 16552
rect 12712 16494 15811 16496
rect 0 16418 800 16448
rect 3233 16418 3299 16421
rect 0 16416 3299 16418
rect 0 16360 3238 16416
rect 3294 16360 3299 16416
rect 0 16358 3299 16360
rect 0 16328 800 16358
rect 3233 16355 3299 16358
rect 8753 16418 8819 16421
rect 8886 16418 8892 16420
rect 8753 16416 8892 16418
rect 8753 16360 8758 16416
rect 8814 16360 8892 16416
rect 8753 16358 8892 16360
rect 8753 16355 8819 16358
rect 8886 16356 8892 16358
rect 8956 16418 8962 16420
rect 12712 16418 12772 16494
rect 15745 16491 15811 16494
rect 8956 16358 12772 16418
rect 8956 16356 8962 16358
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 10685 16282 10751 16285
rect 11421 16282 11487 16285
rect 10685 16280 11487 16282
rect 10685 16224 10690 16280
rect 10746 16224 11426 16280
rect 11482 16224 11487 16280
rect 10685 16222 11487 16224
rect 10685 16219 10751 16222
rect 11421 16219 11487 16222
rect 6545 16146 6611 16149
rect 12617 16146 12683 16149
rect 6545 16144 12683 16146
rect 6545 16088 6550 16144
rect 6606 16088 12622 16144
rect 12678 16088 12683 16144
rect 6545 16086 12683 16088
rect 6545 16083 6611 16086
rect 12617 16083 12683 16086
rect 4337 16010 4403 16013
rect 13118 16010 13124 16012
rect 4337 16008 13124 16010
rect 4337 15952 4342 16008
rect 4398 15952 13124 16008
rect 4337 15950 13124 15952
rect 4337 15947 4403 15950
rect 13118 15948 13124 15950
rect 13188 15948 13194 16012
rect 7230 15812 7236 15876
rect 7300 15874 7306 15876
rect 7373 15874 7439 15877
rect 7300 15872 7439 15874
rect 7300 15816 7378 15872
rect 7434 15816 7439 15872
rect 7300 15814 7439 15816
rect 7300 15812 7306 15814
rect 7373 15811 7439 15814
rect 8477 15874 8543 15877
rect 8886 15874 8892 15876
rect 8477 15872 8892 15874
rect 8477 15816 8482 15872
rect 8538 15816 8892 15872
rect 8477 15814 8892 15816
rect 8477 15811 8543 15814
rect 8886 15812 8892 15814
rect 8956 15812 8962 15876
rect 9673 15874 9739 15877
rect 10501 15876 10567 15877
rect 10174 15874 10180 15876
rect 9673 15872 10180 15874
rect 9673 15816 9678 15872
rect 9734 15816 10180 15872
rect 9673 15814 10180 15816
rect 9673 15811 9739 15814
rect 10174 15812 10180 15814
rect 10244 15812 10250 15876
rect 10501 15874 10548 15876
rect 10456 15872 10548 15874
rect 10456 15816 10506 15872
rect 10456 15814 10548 15816
rect 10501 15812 10548 15814
rect 10612 15812 10618 15876
rect 10501 15811 10567 15812
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 8017 15738 8083 15741
rect 9949 15738 10015 15741
rect 12065 15740 12131 15741
rect 12014 15738 12020 15740
rect 8017 15736 10015 15738
rect 8017 15680 8022 15736
rect 8078 15680 9954 15736
rect 10010 15680 10015 15736
rect 8017 15678 10015 15680
rect 11974 15678 12020 15738
rect 12084 15736 12131 15740
rect 12126 15680 12131 15736
rect 8017 15675 8083 15678
rect 9949 15675 10015 15678
rect 12014 15676 12020 15678
rect 12084 15676 12131 15680
rect 12065 15675 12131 15676
rect 7005 15602 7071 15605
rect 12065 15602 12131 15605
rect 7005 15600 12131 15602
rect 7005 15544 7010 15600
rect 7066 15544 12070 15600
rect 12126 15544 12131 15600
rect 7005 15542 12131 15544
rect 7005 15539 7071 15542
rect 12065 15539 12131 15542
rect 0 15466 800 15496
rect 2957 15466 3023 15469
rect 0 15464 3023 15466
rect 0 15408 2962 15464
rect 3018 15408 3023 15464
rect 0 15406 3023 15408
rect 0 15376 800 15406
rect 2957 15403 3023 15406
rect 5574 15404 5580 15468
rect 5644 15466 5650 15468
rect 7189 15466 7255 15469
rect 5644 15464 7255 15466
rect 5644 15408 7194 15464
rect 7250 15408 7255 15464
rect 5644 15406 7255 15408
rect 5644 15404 5650 15406
rect 7189 15403 7255 15406
rect 8569 15466 8635 15469
rect 14365 15466 14431 15469
rect 8569 15464 14431 15466
rect 8569 15408 8574 15464
rect 8630 15408 14370 15464
rect 14426 15408 14431 15464
rect 8569 15406 14431 15408
rect 8569 15403 8635 15406
rect 14365 15403 14431 15406
rect 9305 15330 9371 15333
rect 11697 15330 11763 15333
rect 11830 15330 11836 15332
rect 9305 15328 11836 15330
rect 9305 15272 9310 15328
rect 9366 15272 11702 15328
rect 11758 15272 11836 15328
rect 9305 15270 11836 15272
rect 9305 15267 9371 15270
rect 11697 15267 11763 15270
rect 11830 15268 11836 15270
rect 11900 15268 11906 15332
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 9673 15196 9739 15197
rect 9622 15132 9628 15196
rect 9692 15194 9739 15196
rect 9857 15194 9923 15197
rect 11697 15194 11763 15197
rect 9692 15192 9784 15194
rect 9734 15136 9784 15192
rect 9692 15134 9784 15136
rect 9857 15192 11763 15194
rect 9857 15136 9862 15192
rect 9918 15136 11702 15192
rect 11758 15136 11763 15192
rect 9857 15134 11763 15136
rect 9692 15132 9739 15134
rect 9673 15131 9739 15132
rect 9857 15131 9923 15134
rect 11697 15131 11763 15134
rect 5625 15058 5691 15061
rect 10961 15058 11027 15061
rect 11513 15060 11579 15061
rect 11462 15058 11468 15060
rect 5625 15056 11027 15058
rect 5625 15000 5630 15056
rect 5686 15000 10966 15056
rect 11022 15000 11027 15056
rect 5625 14998 11027 15000
rect 11386 14998 11468 15058
rect 11532 15058 11579 15060
rect 16389 15058 16455 15061
rect 11532 15056 16455 15058
rect 11574 15000 16394 15056
rect 16450 15000 16455 15056
rect 5625 14995 5691 14998
rect 10961 14995 11027 14998
rect 11462 14996 11468 14998
rect 11532 14998 16455 15000
rect 11532 14996 11579 14998
rect 11513 14995 11579 14996
rect 16389 14995 16455 14998
rect 4797 14922 4863 14925
rect 6821 14922 6887 14925
rect 8017 14922 8083 14925
rect 9305 14924 9371 14925
rect 4797 14920 8083 14922
rect 4797 14864 4802 14920
rect 4858 14864 6826 14920
rect 6882 14864 8022 14920
rect 8078 14864 8083 14920
rect 4797 14862 8083 14864
rect 4797 14859 4863 14862
rect 6821 14859 6887 14862
rect 8017 14859 8083 14862
rect 9254 14860 9260 14924
rect 9324 14922 9371 14924
rect 9581 14922 9647 14925
rect 13997 14922 14063 14925
rect 9324 14920 9416 14922
rect 9366 14864 9416 14920
rect 9324 14862 9416 14864
rect 9581 14920 14063 14922
rect 9581 14864 9586 14920
rect 9642 14864 14002 14920
rect 14058 14864 14063 14920
rect 9581 14862 14063 14864
rect 9324 14860 9371 14862
rect 9305 14859 9371 14860
rect 9581 14859 9647 14862
rect 13997 14859 14063 14862
rect 6269 14786 6335 14789
rect 8293 14786 8359 14789
rect 6269 14784 8359 14786
rect 6269 14728 6274 14784
rect 6330 14728 8298 14784
rect 8354 14728 8359 14784
rect 6269 14726 8359 14728
rect 6269 14723 6335 14726
rect 8293 14723 8359 14726
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 4061 14514 4127 14517
rect 6272 14514 6332 14723
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 6453 14650 6519 14653
rect 10041 14650 10107 14653
rect 6453 14648 10107 14650
rect 6453 14592 6458 14648
rect 6514 14592 10046 14648
rect 10102 14592 10107 14648
rect 6453 14590 10107 14592
rect 6453 14587 6519 14590
rect 10041 14587 10107 14590
rect 10317 14652 10383 14653
rect 10317 14648 10364 14652
rect 10428 14650 10434 14652
rect 10317 14592 10322 14648
rect 10317 14588 10364 14592
rect 10428 14590 10474 14650
rect 10428 14588 10434 14590
rect 10317 14587 10383 14588
rect 4061 14512 6332 14514
rect 4061 14456 4066 14512
rect 4122 14456 6332 14512
rect 4061 14454 6332 14456
rect 6637 14514 6703 14517
rect 11053 14514 11119 14517
rect 12801 14516 12867 14517
rect 12750 14514 12756 14516
rect 6637 14512 11119 14514
rect 6637 14456 6642 14512
rect 6698 14456 11058 14512
rect 11114 14456 11119 14512
rect 6637 14454 11119 14456
rect 12710 14454 12756 14514
rect 12820 14512 12867 14516
rect 12862 14456 12867 14512
rect 4061 14451 4127 14454
rect 6637 14451 6703 14454
rect 11053 14451 11119 14454
rect 12750 14452 12756 14454
rect 12820 14452 12867 14456
rect 12801 14451 12867 14452
rect 0 14378 800 14408
rect 1853 14378 1919 14381
rect 0 14376 1919 14378
rect 0 14320 1858 14376
rect 1914 14320 1919 14376
rect 0 14318 1919 14320
rect 0 14288 800 14318
rect 1853 14315 1919 14318
rect 2405 14378 2471 14381
rect 5993 14378 6059 14381
rect 7097 14378 7163 14381
rect 9857 14378 9923 14381
rect 2405 14376 6930 14378
rect 2405 14320 2410 14376
rect 2466 14320 5998 14376
rect 6054 14320 6930 14376
rect 2405 14318 6930 14320
rect 2405 14315 2471 14318
rect 5993 14315 6059 14318
rect 6870 14242 6930 14318
rect 7097 14376 9923 14378
rect 7097 14320 7102 14376
rect 7158 14320 9862 14376
rect 9918 14320 9923 14376
rect 7097 14318 9923 14320
rect 7097 14315 7163 14318
rect 9857 14315 9923 14318
rect 10041 14378 10107 14381
rect 12985 14378 13051 14381
rect 10041 14376 13051 14378
rect 10041 14320 10046 14376
rect 10102 14320 12990 14376
rect 13046 14320 13051 14376
rect 10041 14318 13051 14320
rect 10041 14315 10107 14318
rect 12985 14315 13051 14318
rect 7741 14242 7807 14245
rect 6870 14240 7807 14242
rect 6870 14184 7746 14240
rect 7802 14184 7807 14240
rect 6870 14182 7807 14184
rect 7741 14179 7807 14182
rect 8845 14242 8911 14245
rect 9857 14242 9923 14245
rect 8845 14240 9923 14242
rect 8845 14184 8850 14240
rect 8906 14184 9862 14240
rect 9918 14184 9923 14240
rect 8845 14182 9923 14184
rect 8845 14179 8911 14182
rect 9857 14179 9923 14182
rect 10174 14180 10180 14244
rect 10244 14242 10250 14244
rect 10685 14242 10751 14245
rect 10244 14240 10751 14242
rect 10244 14184 10690 14240
rect 10746 14184 10751 14240
rect 10244 14182 10751 14184
rect 10244 14180 10250 14182
rect 10685 14179 10751 14182
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 9673 14106 9739 14109
rect 9990 14106 9996 14108
rect 9673 14104 9996 14106
rect 9673 14048 9678 14104
rect 9734 14048 9996 14104
rect 9673 14046 9996 14048
rect 9673 14043 9739 14046
rect 9990 14044 9996 14046
rect 10060 14044 10066 14108
rect 10409 14106 10475 14109
rect 10136 14104 10475 14106
rect 10136 14048 10414 14104
rect 10470 14048 10475 14104
rect 10136 14046 10475 14048
rect 5257 13970 5323 13973
rect 9765 13972 9831 13973
rect 9622 13970 9628 13972
rect 5257 13968 9628 13970
rect 5257 13912 5262 13968
rect 5318 13912 9628 13968
rect 5257 13910 9628 13912
rect 5257 13907 5323 13910
rect 9622 13908 9628 13910
rect 9692 13908 9698 13972
rect 9765 13968 9812 13972
rect 9876 13970 9882 13972
rect 9765 13912 9770 13968
rect 9765 13908 9812 13912
rect 9876 13910 9922 13970
rect 9876 13908 9882 13910
rect 9765 13907 9831 13908
rect 4245 13834 4311 13837
rect 6637 13834 6703 13837
rect 10136 13834 10196 14046
rect 10409 14043 10475 14046
rect 10593 14106 10659 14109
rect 11329 14106 11395 14109
rect 10593 14104 11395 14106
rect 10593 14048 10598 14104
rect 10654 14048 11334 14104
rect 11390 14048 11395 14104
rect 10593 14046 11395 14048
rect 10593 14043 10659 14046
rect 11329 14043 11395 14046
rect 10409 13970 10475 13973
rect 12341 13970 12407 13973
rect 10409 13968 12407 13970
rect 10409 13912 10414 13968
rect 10470 13912 12346 13968
rect 12402 13912 12407 13968
rect 10409 13910 12407 13912
rect 10409 13907 10475 13910
rect 12341 13907 12407 13910
rect 4245 13832 6562 13834
rect 4245 13776 4250 13832
rect 4306 13776 6562 13832
rect 4245 13774 6562 13776
rect 4245 13771 4311 13774
rect 6502 13698 6562 13774
rect 6637 13832 10196 13834
rect 6637 13776 6642 13832
rect 6698 13776 10196 13832
rect 6637 13774 10196 13776
rect 10685 13834 10751 13837
rect 12433 13834 12499 13837
rect 10685 13832 12499 13834
rect 10685 13776 10690 13832
rect 10746 13776 12438 13832
rect 12494 13776 12499 13832
rect 10685 13774 12499 13776
rect 6637 13771 6703 13774
rect 10685 13771 10751 13774
rect 12433 13771 12499 13774
rect 10041 13698 10107 13701
rect 10225 13698 10291 13701
rect 12433 13700 12499 13701
rect 12382 13698 12388 13700
rect 6502 13696 10291 13698
rect 6502 13640 10046 13696
rect 10102 13640 10230 13696
rect 10286 13640 10291 13696
rect 6502 13638 10291 13640
rect 12342 13638 12388 13698
rect 12452 13696 12499 13700
rect 12494 13640 12499 13696
rect 10041 13635 10107 13638
rect 10225 13635 10291 13638
rect 12382 13636 12388 13638
rect 12452 13636 12499 13640
rect 12433 13635 12499 13636
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 2037 13562 2103 13565
rect 8017 13562 8083 13565
rect 11421 13562 11487 13565
rect 11646 13562 11652 13564
rect 2037 13560 3204 13562
rect 2037 13504 2042 13560
rect 2098 13504 3204 13560
rect 2037 13502 3204 13504
rect 2037 13499 2103 13502
rect 0 13426 800 13456
rect 2957 13426 3023 13429
rect 0 13424 3023 13426
rect 0 13368 2962 13424
rect 3018 13368 3023 13424
rect 0 13366 3023 13368
rect 3144 13426 3204 13502
rect 8017 13560 9552 13562
rect 8017 13504 8022 13560
rect 8078 13504 9552 13560
rect 8017 13502 9552 13504
rect 8017 13499 8083 13502
rect 6637 13426 6703 13429
rect 3144 13424 6703 13426
rect 3144 13368 6642 13424
rect 6698 13368 6703 13424
rect 3144 13366 6703 13368
rect 9492 13426 9552 13502
rect 11421 13560 11652 13562
rect 11421 13504 11426 13560
rect 11482 13504 11652 13560
rect 11421 13502 11652 13504
rect 11421 13499 11487 13502
rect 11646 13500 11652 13502
rect 11716 13500 11722 13564
rect 12157 13562 12223 13565
rect 12382 13562 12388 13564
rect 12157 13560 12388 13562
rect 12157 13504 12162 13560
rect 12218 13504 12388 13560
rect 12157 13502 12388 13504
rect 12157 13499 12223 13502
rect 12382 13500 12388 13502
rect 12452 13500 12458 13564
rect 13261 13426 13327 13429
rect 9492 13424 13327 13426
rect 9492 13368 13266 13424
rect 13322 13368 13327 13424
rect 9492 13366 13327 13368
rect 0 13336 800 13366
rect 2957 13363 3023 13366
rect 6637 13363 6703 13366
rect 13261 13363 13327 13366
rect 4705 13290 4771 13293
rect 10961 13290 11027 13293
rect 4705 13288 11027 13290
rect 4705 13232 4710 13288
rect 4766 13232 10966 13288
rect 11022 13232 11027 13288
rect 4705 13230 11027 13232
rect 4705 13227 4771 13230
rect 10961 13227 11027 13230
rect 11513 13290 11579 13293
rect 11973 13290 12039 13293
rect 12198 13290 12204 13292
rect 11513 13288 12204 13290
rect 11513 13232 11518 13288
rect 11574 13232 11978 13288
rect 12034 13232 12204 13288
rect 11513 13230 12204 13232
rect 11513 13227 11579 13230
rect 11973 13227 12039 13230
rect 12198 13228 12204 13230
rect 12268 13228 12274 13292
rect 9070 13092 9076 13156
rect 9140 13154 9146 13156
rect 11053 13154 11119 13157
rect 9140 13152 11119 13154
rect 9140 13096 11058 13152
rect 11114 13096 11119 13152
rect 9140 13094 11119 13096
rect 9140 13092 9146 13094
rect 11053 13091 11119 13094
rect 12341 13154 12407 13157
rect 13077 13154 13143 13157
rect 12341 13152 13143 13154
rect 12341 13096 12346 13152
rect 12402 13096 13082 13152
rect 13138 13096 13143 13152
rect 12341 13094 13143 13096
rect 12341 13091 12407 13094
rect 13077 13091 13143 13094
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 4245 13018 4311 13021
rect 5901 13018 5967 13021
rect 4245 13016 5967 13018
rect 4245 12960 4250 13016
rect 4306 12960 5906 13016
rect 5962 12960 5967 13016
rect 4245 12958 5967 12960
rect 4245 12955 4311 12958
rect 5901 12955 5967 12958
rect 8845 13018 8911 13021
rect 9949 13018 10015 13021
rect 10542 13018 10548 13020
rect 8845 13016 10015 13018
rect 8845 12960 8850 13016
rect 8906 12960 9954 13016
rect 10010 12960 10015 13016
rect 8845 12958 10015 12960
rect 10466 12958 10548 13018
rect 8845 12955 8911 12958
rect 9949 12955 10015 12958
rect 10542 12956 10548 12958
rect 10612 13018 10618 13020
rect 12344 13018 12404 13091
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 10612 12958 12404 13018
rect 12525 13020 12591 13021
rect 12525 13016 12572 13020
rect 12636 13018 12642 13020
rect 12525 12960 12530 13016
rect 10612 12956 10656 12958
rect 4797 12882 4863 12885
rect 5073 12882 5139 12885
rect 4797 12880 5139 12882
rect 4797 12824 4802 12880
rect 4858 12824 5078 12880
rect 5134 12824 5139 12880
rect 4797 12822 5139 12824
rect 4797 12819 4863 12822
rect 5073 12819 5139 12822
rect 6545 12882 6611 12885
rect 8845 12882 8911 12885
rect 6545 12880 8911 12882
rect 6545 12824 6550 12880
rect 6606 12824 8850 12880
rect 8906 12824 8911 12880
rect 6545 12822 8911 12824
rect 6545 12819 6611 12822
rect 8845 12819 8911 12822
rect 9438 12820 9444 12884
rect 9508 12882 9514 12884
rect 10041 12882 10107 12885
rect 9508 12880 10107 12882
rect 9508 12824 10046 12880
rect 10102 12824 10107 12880
rect 9508 12822 10107 12824
rect 9508 12820 9514 12822
rect 10041 12819 10107 12822
rect 2681 12746 2747 12749
rect 8017 12746 8083 12749
rect 9254 12746 9260 12748
rect 2681 12744 6332 12746
rect 2681 12688 2686 12744
rect 2742 12688 6332 12744
rect 2681 12686 6332 12688
rect 2681 12683 2747 12686
rect 5874 12544 6194 12545
rect 0 12474 800 12504
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 2865 12474 2931 12477
rect 0 12472 2931 12474
rect 0 12416 2870 12472
rect 2926 12416 2931 12472
rect 0 12414 2931 12416
rect 6272 12474 6332 12686
rect 8017 12744 9260 12746
rect 8017 12688 8022 12744
rect 8078 12688 9260 12744
rect 8017 12686 9260 12688
rect 8017 12683 8083 12686
rect 9254 12684 9260 12686
rect 9324 12746 9330 12748
rect 10409 12746 10475 12749
rect 9324 12744 10475 12746
rect 9324 12688 10414 12744
rect 10470 12688 10475 12744
rect 9324 12686 10475 12688
rect 9324 12684 9330 12686
rect 10409 12683 10475 12686
rect 6729 12610 6795 12613
rect 10596 12610 10656 12956
rect 12525 12956 12572 12960
rect 12636 12958 12682 13018
rect 12636 12956 12642 12958
rect 12525 12955 12591 12956
rect 11278 12820 11284 12884
rect 11348 12882 11354 12884
rect 12934 12882 12940 12884
rect 11348 12822 12940 12882
rect 11348 12820 11354 12822
rect 12934 12820 12940 12822
rect 13004 12882 13010 12884
rect 14549 12882 14615 12885
rect 13004 12880 14615 12882
rect 13004 12824 14554 12880
rect 14610 12824 14615 12880
rect 13004 12822 14615 12824
rect 13004 12820 13010 12822
rect 14549 12819 14615 12822
rect 11053 12746 11119 12749
rect 13813 12746 13879 12749
rect 11053 12744 13879 12746
rect 11053 12688 11058 12744
rect 11114 12688 13818 12744
rect 13874 12688 13879 12744
rect 11053 12686 13879 12688
rect 11053 12683 11119 12686
rect 13813 12683 13879 12686
rect 12801 12610 12867 12613
rect 6729 12608 10656 12610
rect 6729 12552 6734 12608
rect 6790 12552 10656 12608
rect 6729 12550 10656 12552
rect 12574 12608 12867 12610
rect 12574 12552 12806 12608
rect 12862 12552 12867 12608
rect 12574 12550 12867 12552
rect 6729 12547 6795 12550
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 12574 12477 12634 12550
rect 12801 12547 12867 12550
rect 13118 12548 13124 12612
rect 13188 12610 13194 12612
rect 13261 12610 13327 12613
rect 13188 12608 13327 12610
rect 13188 12552 13266 12608
rect 13322 12552 13327 12608
rect 13188 12550 13327 12552
rect 13188 12548 13194 12550
rect 13261 12547 13327 12550
rect 9857 12474 9923 12477
rect 11973 12476 12039 12477
rect 11973 12474 12020 12476
rect 6272 12472 9923 12474
rect 6272 12416 9862 12472
rect 9918 12416 9923 12472
rect 6272 12414 9923 12416
rect 11928 12472 12020 12474
rect 11928 12416 11978 12472
rect 11928 12414 12020 12416
rect 0 12384 800 12414
rect 2865 12411 2931 12414
rect 9857 12411 9923 12414
rect 11973 12412 12020 12414
rect 12084 12412 12090 12476
rect 12525 12472 12634 12477
rect 12525 12416 12530 12472
rect 12586 12416 12634 12472
rect 12525 12414 12634 12416
rect 11973 12411 12039 12412
rect 12525 12411 12591 12414
rect 12750 12412 12756 12476
rect 12820 12474 12826 12476
rect 13077 12474 13143 12477
rect 12820 12472 13143 12474
rect 12820 12416 13082 12472
rect 13138 12416 13143 12472
rect 12820 12414 13143 12416
rect 12820 12412 12826 12414
rect 13077 12411 13143 12414
rect 2037 12338 2103 12341
rect 12750 12338 12756 12340
rect 2037 12336 12756 12338
rect 2037 12280 2042 12336
rect 2098 12280 12756 12336
rect 2037 12278 12756 12280
rect 2037 12275 2103 12278
rect 12750 12276 12756 12278
rect 12820 12276 12826 12340
rect 5165 12202 5231 12205
rect 6637 12202 6703 12205
rect 5165 12200 6703 12202
rect 5165 12144 5170 12200
rect 5226 12144 6642 12200
rect 6698 12144 6703 12200
rect 5165 12142 6703 12144
rect 5165 12139 5231 12142
rect 6637 12139 6703 12142
rect 7373 12202 7439 12205
rect 8937 12204 9003 12205
rect 7373 12200 8816 12202
rect 7373 12144 7378 12200
rect 7434 12144 8816 12200
rect 7373 12142 8816 12144
rect 7373 12139 7439 12142
rect 8756 12066 8816 12142
rect 8886 12140 8892 12204
rect 8956 12202 9003 12204
rect 9305 12202 9371 12205
rect 9622 12202 9628 12204
rect 8956 12200 9048 12202
rect 8998 12144 9048 12200
rect 8956 12142 9048 12144
rect 9305 12200 9628 12202
rect 9305 12144 9310 12200
rect 9366 12144 9628 12200
rect 9305 12142 9628 12144
rect 8956 12140 9003 12142
rect 8937 12139 9003 12140
rect 9305 12139 9371 12142
rect 9622 12140 9628 12142
rect 9692 12140 9698 12204
rect 9990 12140 9996 12204
rect 10060 12202 10066 12204
rect 10133 12202 10199 12205
rect 10060 12200 10199 12202
rect 10060 12144 10138 12200
rect 10194 12144 10199 12200
rect 10060 12142 10199 12144
rect 10060 12140 10066 12142
rect 10133 12139 10199 12142
rect 10358 12140 10364 12204
rect 10428 12202 10434 12204
rect 11329 12202 11395 12205
rect 10428 12200 11395 12202
rect 10428 12144 11334 12200
rect 11390 12144 11395 12200
rect 10428 12142 11395 12144
rect 10428 12140 10434 12142
rect 11329 12139 11395 12142
rect 11605 12202 11671 12205
rect 15009 12202 15075 12205
rect 11605 12200 15075 12202
rect 11605 12144 11610 12200
rect 11666 12144 15014 12200
rect 15070 12144 15075 12200
rect 11605 12142 15075 12144
rect 11605 12139 11671 12142
rect 15009 12139 15075 12142
rect 11513 12066 11579 12069
rect 8756 12064 11579 12066
rect 8756 12008 11518 12064
rect 11574 12008 11579 12064
rect 8756 12006 11579 12008
rect 11513 12003 11579 12006
rect 11646 12004 11652 12068
rect 11716 12066 11722 12068
rect 12433 12066 12499 12069
rect 11716 12064 12499 12066
rect 11716 12008 12438 12064
rect 12494 12008 12499 12064
rect 11716 12006 12499 12008
rect 11716 12004 11722 12006
rect 12433 12003 12499 12006
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 4337 11930 4403 11933
rect 5349 11930 5415 11933
rect 7230 11930 7236 11932
rect 4337 11928 7236 11930
rect 4337 11872 4342 11928
rect 4398 11872 5354 11928
rect 5410 11872 7236 11928
rect 4337 11870 7236 11872
rect 4337 11867 4403 11870
rect 5349 11867 5415 11870
rect 7230 11868 7236 11870
rect 7300 11868 7306 11932
rect 9254 11868 9260 11932
rect 9324 11930 9330 11932
rect 9581 11930 9647 11933
rect 9324 11928 9647 11930
rect 9324 11872 9586 11928
rect 9642 11872 9647 11928
rect 9324 11870 9647 11872
rect 9324 11868 9330 11870
rect 9581 11867 9647 11870
rect 12014 11868 12020 11932
rect 12084 11930 12090 11932
rect 12157 11930 12223 11933
rect 12084 11928 12223 11930
rect 12084 11872 12162 11928
rect 12218 11872 12223 11928
rect 12084 11870 12223 11872
rect 12084 11868 12090 11870
rect 12157 11867 12223 11870
rect 3969 11794 4035 11797
rect 13077 11794 13143 11797
rect 3969 11792 13143 11794
rect 3969 11736 3974 11792
rect 4030 11736 13082 11792
rect 13138 11736 13143 11792
rect 3969 11734 13143 11736
rect 3969 11731 4035 11734
rect 13077 11731 13143 11734
rect 3141 11658 3207 11661
rect 7925 11658 7991 11661
rect 9765 11658 9831 11661
rect 3141 11656 6332 11658
rect 3141 11600 3146 11656
rect 3202 11600 6332 11656
rect 3141 11598 6332 11600
rect 3141 11595 3207 11598
rect 3969 11522 4035 11525
rect 5574 11522 5580 11524
rect 3969 11520 5580 11522
rect 3969 11464 3974 11520
rect 4030 11464 5580 11520
rect 3969 11462 5580 11464
rect 3969 11459 4035 11462
rect 5574 11460 5580 11462
rect 5644 11460 5650 11524
rect 6272 11522 6332 11598
rect 7925 11656 9831 11658
rect 7925 11600 7930 11656
rect 7986 11600 9770 11656
rect 9826 11600 9831 11656
rect 7925 11598 9831 11600
rect 7925 11595 7991 11598
rect 9765 11595 9831 11598
rect 11237 11658 11303 11661
rect 11646 11658 11652 11660
rect 11237 11656 11652 11658
rect 11237 11600 11242 11656
rect 11298 11600 11652 11656
rect 11237 11598 11652 11600
rect 11237 11595 11303 11598
rect 11646 11596 11652 11598
rect 11716 11596 11722 11660
rect 12065 11656 12131 11661
rect 12065 11600 12070 11656
rect 12126 11600 12131 11656
rect 12065 11595 12131 11600
rect 9254 11522 9260 11524
rect 6272 11462 9260 11522
rect 9254 11460 9260 11462
rect 9324 11460 9330 11524
rect 11513 11522 11579 11525
rect 12068 11522 12128 11595
rect 11513 11520 12128 11522
rect 11513 11464 11518 11520
rect 11574 11464 12128 11520
rect 11513 11462 12128 11464
rect 11513 11459 11579 11462
rect 5874 11456 6194 11457
rect 0 11386 800 11416
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 1393 11386 1459 11389
rect 0 11384 1459 11386
rect 0 11328 1398 11384
rect 1454 11328 1459 11384
rect 0 11326 1459 11328
rect 0 11296 800 11326
rect 1393 11323 1459 11326
rect 10317 11388 10383 11389
rect 10317 11384 10364 11388
rect 10428 11386 10434 11388
rect 10317 11328 10322 11384
rect 10317 11324 10364 11328
rect 10428 11326 10474 11386
rect 10428 11324 10434 11326
rect 10317 11323 10383 11324
rect 4613 11250 4679 11253
rect 8845 11250 8911 11253
rect 4613 11248 8911 11250
rect 4613 11192 4618 11248
rect 4674 11192 8850 11248
rect 8906 11192 8911 11248
rect 4613 11190 8911 11192
rect 4613 11187 4679 11190
rect 8845 11187 8911 11190
rect 11646 11188 11652 11252
rect 11716 11250 11722 11252
rect 11973 11250 12039 11253
rect 11716 11248 12039 11250
rect 11716 11192 11978 11248
rect 12034 11192 12039 11248
rect 11716 11190 12039 11192
rect 11716 11188 11722 11190
rect 11973 11187 12039 11190
rect 12157 11250 12223 11253
rect 13854 11250 13860 11252
rect 12157 11248 13860 11250
rect 12157 11192 12162 11248
rect 12218 11192 13860 11248
rect 12157 11190 13860 11192
rect 12157 11187 12223 11190
rect 13854 11188 13860 11190
rect 13924 11250 13930 11252
rect 14181 11250 14247 11253
rect 13924 11248 14247 11250
rect 13924 11192 14186 11248
rect 14242 11192 14247 11248
rect 13924 11190 14247 11192
rect 13924 11188 13930 11190
rect 14181 11187 14247 11190
rect 7465 11114 7531 11117
rect 12341 11114 12407 11117
rect 13261 11114 13327 11117
rect 7465 11112 12407 11114
rect 7465 11056 7470 11112
rect 7526 11056 12346 11112
rect 12402 11056 12407 11112
rect 7465 11054 12407 11056
rect 7465 11051 7531 11054
rect 12341 11051 12407 11054
rect 13126 11112 13327 11114
rect 13126 11056 13266 11112
rect 13322 11056 13327 11112
rect 13126 11054 13327 11056
rect 10041 10978 10107 10981
rect 10174 10978 10180 10980
rect 10041 10976 10180 10978
rect 10041 10920 10046 10976
rect 10102 10920 10180 10976
rect 10041 10918 10180 10920
rect 10041 10915 10107 10918
rect 10174 10916 10180 10918
rect 10244 10916 10250 10980
rect 10501 10978 10567 10981
rect 13126 10978 13186 11054
rect 13261 11051 13327 11054
rect 13537 11114 13603 11117
rect 13670 11114 13676 11116
rect 13537 11112 13676 11114
rect 13537 11056 13542 11112
rect 13598 11056 13676 11112
rect 13537 11054 13676 11056
rect 13537 11051 13603 11054
rect 13670 11052 13676 11054
rect 13740 11052 13746 11116
rect 10501 10976 13186 10978
rect 10501 10920 10506 10976
rect 10562 10920 13186 10976
rect 10501 10918 13186 10920
rect 10501 10915 10567 10918
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 10685 10842 10751 10845
rect 13077 10842 13143 10845
rect 10685 10840 13143 10842
rect 10685 10784 10690 10840
rect 10746 10784 13082 10840
rect 13138 10784 13143 10840
rect 10685 10782 13143 10784
rect 10685 10779 10751 10782
rect 13077 10779 13143 10782
rect 3141 10706 3207 10709
rect 5441 10706 5507 10709
rect 3141 10704 5507 10706
rect 3141 10648 3146 10704
rect 3202 10648 5446 10704
rect 5502 10648 5507 10704
rect 3141 10646 5507 10648
rect 3141 10643 3207 10646
rect 5441 10643 5507 10646
rect 8886 10644 8892 10708
rect 8956 10706 8962 10708
rect 9029 10706 9095 10709
rect 8956 10704 9095 10706
rect 8956 10648 9034 10704
rect 9090 10648 9095 10704
rect 8956 10646 9095 10648
rect 8956 10644 8962 10646
rect 9029 10643 9095 10646
rect 12198 10644 12204 10708
rect 12268 10706 12274 10708
rect 13445 10706 13511 10709
rect 12268 10704 13511 10706
rect 12268 10648 13450 10704
rect 13506 10648 13511 10704
rect 12268 10646 13511 10648
rect 12268 10644 12274 10646
rect 13445 10643 13511 10646
rect 2313 10570 2379 10573
rect 13077 10570 13143 10573
rect 2313 10568 13143 10570
rect 2313 10512 2318 10568
rect 2374 10512 13082 10568
rect 13138 10512 13143 10568
rect 2313 10510 13143 10512
rect 2313 10507 2379 10510
rect 13077 10507 13143 10510
rect 0 10434 800 10464
rect 1853 10434 1919 10437
rect 0 10432 1919 10434
rect 0 10376 1858 10432
rect 1914 10376 1919 10432
rect 0 10374 1919 10376
rect 0 10344 800 10374
rect 1853 10371 1919 10374
rect 8109 10434 8175 10437
rect 10409 10434 10475 10437
rect 8109 10432 10475 10434
rect 8109 10376 8114 10432
rect 8170 10376 10414 10432
rect 10470 10376 10475 10432
rect 8109 10374 10475 10376
rect 8109 10371 8175 10374
rect 10409 10371 10475 10374
rect 11697 10434 11763 10437
rect 12433 10436 12499 10437
rect 12382 10434 12388 10436
rect 11697 10432 12388 10434
rect 12452 10434 12499 10436
rect 12452 10432 12544 10434
rect 11697 10376 11702 10432
rect 11758 10376 12388 10432
rect 12494 10376 12544 10432
rect 11697 10374 12388 10376
rect 11697 10371 11763 10374
rect 12382 10372 12388 10374
rect 12452 10374 12544 10376
rect 12452 10372 12499 10374
rect 12433 10371 12499 10372
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 9489 10298 9555 10301
rect 10409 10298 10475 10301
rect 9489 10296 10475 10298
rect 9489 10240 9494 10296
rect 9550 10240 10414 10296
rect 10470 10240 10475 10296
rect 9489 10238 10475 10240
rect 9489 10235 9555 10238
rect 10409 10235 10475 10238
rect 11329 10298 11395 10301
rect 14365 10298 14431 10301
rect 11329 10296 14431 10298
rect 11329 10240 11334 10296
rect 11390 10240 14370 10296
rect 14426 10240 14431 10296
rect 11329 10238 14431 10240
rect 11329 10235 11395 10238
rect 14365 10235 14431 10238
rect 3141 10162 3207 10165
rect 12709 10162 12775 10165
rect 3141 10160 12775 10162
rect 3141 10104 3146 10160
rect 3202 10104 12714 10160
rect 12770 10104 12775 10160
rect 3141 10102 12775 10104
rect 3141 10099 3207 10102
rect 12709 10099 12775 10102
rect 12985 10162 13051 10165
rect 13118 10162 13124 10164
rect 12985 10160 13124 10162
rect 12985 10104 12990 10160
rect 13046 10104 13124 10160
rect 12985 10102 13124 10104
rect 12985 10099 13051 10102
rect 13118 10100 13124 10102
rect 13188 10100 13194 10164
rect 3877 10026 3943 10029
rect 14181 10026 14247 10029
rect 3877 10024 14247 10026
rect 3877 9968 3882 10024
rect 3938 9968 14186 10024
rect 14242 9968 14247 10024
rect 3877 9966 14247 9968
rect 3877 9963 3943 9966
rect 14181 9963 14247 9966
rect 14825 10026 14891 10029
rect 16200 10026 17000 10056
rect 14825 10024 17000 10026
rect 14825 9968 14830 10024
rect 14886 9968 17000 10024
rect 14825 9966 17000 9968
rect 14825 9963 14891 9966
rect 16200 9936 17000 9966
rect 10542 9828 10548 9892
rect 10612 9890 10618 9892
rect 12566 9890 12572 9892
rect 10612 9830 12572 9890
rect 10612 9828 10618 9830
rect 12566 9828 12572 9830
rect 12636 9828 12642 9892
rect 12750 9828 12756 9892
rect 12820 9890 12826 9892
rect 12985 9890 13051 9893
rect 12820 9888 13051 9890
rect 12820 9832 12990 9888
rect 13046 9832 13051 9888
rect 12820 9830 13051 9832
rect 12820 9828 12826 9830
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 9489 9754 9555 9757
rect 10317 9754 10383 9757
rect 9489 9752 10383 9754
rect 9489 9696 9494 9752
rect 9550 9696 10322 9752
rect 10378 9696 10383 9752
rect 9489 9694 10383 9696
rect 9489 9691 9555 9694
rect 10317 9691 10383 9694
rect 10869 9754 10935 9757
rect 11513 9754 11579 9757
rect 10869 9752 11579 9754
rect 10869 9696 10874 9752
rect 10930 9696 11518 9752
rect 11574 9696 11579 9752
rect 10869 9694 11579 9696
rect 10869 9691 10935 9694
rect 11513 9691 11579 9694
rect 11789 9752 11855 9757
rect 12341 9754 12407 9757
rect 11789 9696 11794 9752
rect 11850 9696 11855 9752
rect 11789 9691 11855 9696
rect 12022 9752 12407 9754
rect 12022 9696 12346 9752
rect 12402 9696 12407 9752
rect 12022 9694 12407 9696
rect 12574 9754 12634 9828
rect 12985 9827 13051 9830
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 12893 9754 12959 9757
rect 12574 9752 12959 9754
rect 12574 9696 12898 9752
rect 12954 9696 12959 9752
rect 12574 9694 12959 9696
rect 4061 9618 4127 9621
rect 8477 9618 8543 9621
rect 10133 9620 10199 9621
rect 8886 9618 8892 9620
rect 4061 9616 8402 9618
rect 4061 9560 4066 9616
rect 4122 9560 8402 9616
rect 4061 9558 8402 9560
rect 4061 9555 4127 9558
rect 0 9482 800 9512
rect 3049 9482 3115 9485
rect 0 9480 3115 9482
rect 0 9424 3054 9480
rect 3110 9424 3115 9480
rect 0 9422 3115 9424
rect 0 9392 800 9422
rect 3049 9419 3115 9422
rect 3509 9482 3575 9485
rect 7189 9482 7255 9485
rect 3509 9480 7255 9482
rect 3509 9424 3514 9480
rect 3570 9424 7194 9480
rect 7250 9424 7255 9480
rect 3509 9422 7255 9424
rect 8342 9482 8402 9558
rect 8477 9616 8892 9618
rect 8477 9560 8482 9616
rect 8538 9560 8892 9616
rect 8477 9558 8892 9560
rect 8477 9555 8543 9558
rect 8886 9556 8892 9558
rect 8956 9556 8962 9620
rect 10133 9618 10180 9620
rect 10088 9616 10180 9618
rect 10088 9560 10138 9616
rect 10088 9558 10180 9560
rect 10133 9556 10180 9558
rect 10244 9556 10250 9620
rect 10317 9618 10383 9621
rect 11421 9618 11487 9621
rect 10317 9616 11487 9618
rect 10317 9560 10322 9616
rect 10378 9560 11426 9616
rect 11482 9560 11487 9616
rect 10317 9558 11487 9560
rect 10133 9555 10199 9556
rect 10317 9555 10383 9558
rect 11421 9555 11487 9558
rect 10133 9482 10199 9485
rect 11329 9484 11395 9485
rect 11278 9482 11284 9484
rect 8342 9480 10199 9482
rect 8342 9424 10138 9480
rect 10194 9424 10199 9480
rect 8342 9422 10199 9424
rect 11202 9422 11284 9482
rect 11348 9482 11395 9484
rect 11792 9482 11852 9691
rect 11348 9480 11852 9482
rect 11390 9424 11852 9480
rect 3509 9419 3575 9422
rect 7189 9419 7255 9422
rect 10133 9419 10199 9422
rect 11278 9420 11284 9422
rect 11348 9422 11852 9424
rect 11348 9420 11395 9422
rect 11329 9419 11395 9420
rect 9305 9346 9371 9349
rect 9438 9346 9444 9348
rect 9305 9344 9444 9346
rect 9305 9288 9310 9344
rect 9366 9288 9444 9344
rect 9305 9286 9444 9288
rect 9305 9283 9371 9286
rect 9438 9284 9444 9286
rect 9508 9346 9514 9348
rect 10593 9346 10659 9349
rect 9508 9344 10659 9346
rect 9508 9288 10598 9344
rect 10654 9288 10659 9344
rect 9508 9286 10659 9288
rect 9508 9284 9514 9286
rect 10593 9283 10659 9286
rect 11646 9284 11652 9348
rect 11716 9346 11722 9348
rect 11716 9286 11898 9346
rect 11716 9284 11722 9286
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 4153 9210 4219 9213
rect 5625 9210 5691 9213
rect 4153 9208 5691 9210
rect 4153 9152 4158 9208
rect 4214 9152 5630 9208
rect 5686 9152 5691 9208
rect 4153 9150 5691 9152
rect 4153 9147 4219 9150
rect 5625 9147 5691 9150
rect 7741 9210 7807 9213
rect 9121 9210 9187 9213
rect 7741 9208 9187 9210
rect 7741 9152 7746 9208
rect 7802 9152 9126 9208
rect 9182 9152 9187 9208
rect 7741 9150 9187 9152
rect 7741 9147 7807 9150
rect 9121 9147 9187 9150
rect 9581 9210 9647 9213
rect 11605 9212 11671 9213
rect 9990 9210 9996 9212
rect 9581 9208 9996 9210
rect 9581 9152 9586 9208
rect 9642 9152 9996 9208
rect 9581 9150 9996 9152
rect 9581 9147 9647 9150
rect 9990 9148 9996 9150
rect 10060 9148 10066 9212
rect 11605 9208 11652 9212
rect 11716 9210 11722 9212
rect 11605 9152 11610 9208
rect 11605 9148 11652 9152
rect 11716 9150 11762 9210
rect 11716 9148 11722 9150
rect 11605 9147 11671 9148
rect 11838 9077 11898 9286
rect 4521 9074 4587 9077
rect 11053 9074 11119 9077
rect 11462 9074 11468 9076
rect 4521 9072 11468 9074
rect 4521 9016 4526 9072
rect 4582 9016 11058 9072
rect 11114 9016 11468 9072
rect 4521 9014 11468 9016
rect 4521 9011 4587 9014
rect 11053 9011 11119 9014
rect 11462 9012 11468 9014
rect 11532 9012 11538 9076
rect 11838 9072 11947 9077
rect 11838 9016 11886 9072
rect 11942 9016 11947 9072
rect 11838 9014 11947 9016
rect 12022 9074 12082 9694
rect 12341 9691 12407 9694
rect 12893 9691 12959 9694
rect 12157 9618 12223 9621
rect 12566 9618 12572 9620
rect 12157 9616 12572 9618
rect 12157 9560 12162 9616
rect 12218 9560 12572 9616
rect 12157 9558 12572 9560
rect 12157 9555 12223 9558
rect 12566 9556 12572 9558
rect 12636 9556 12642 9620
rect 12157 9210 12223 9213
rect 12893 9210 12959 9213
rect 14457 9210 14523 9213
rect 12157 9208 14523 9210
rect 12157 9152 12162 9208
rect 12218 9152 12898 9208
rect 12954 9152 14462 9208
rect 14518 9152 14523 9208
rect 12157 9150 14523 9152
rect 12157 9147 12223 9150
rect 12893 9147 12959 9150
rect 14457 9147 14523 9150
rect 12617 9074 12683 9077
rect 12022 9072 12683 9074
rect 12022 9016 12622 9072
rect 12678 9016 12683 9072
rect 12022 9014 12683 9016
rect 11881 9011 11947 9014
rect 12617 9011 12683 9014
rect 12893 9074 12959 9077
rect 13721 9074 13787 9077
rect 12893 9072 13787 9074
rect 12893 9016 12898 9072
rect 12954 9016 13726 9072
rect 13782 9016 13787 9072
rect 12893 9014 13787 9016
rect 12893 9011 12959 9014
rect 13721 9011 13787 9014
rect 5533 8938 5599 8941
rect 11145 8938 11211 8941
rect 5533 8936 11211 8938
rect 5533 8880 5538 8936
rect 5594 8880 11150 8936
rect 11206 8880 11211 8936
rect 5533 8878 11211 8880
rect 5533 8875 5599 8878
rect 11145 8875 11211 8878
rect 11329 8938 11395 8941
rect 12341 8940 12407 8941
rect 12014 8938 12020 8940
rect 11329 8936 12020 8938
rect 11329 8880 11334 8936
rect 11390 8880 12020 8936
rect 11329 8878 12020 8880
rect 11329 8875 11395 8878
rect 12014 8876 12020 8878
rect 12084 8876 12090 8940
rect 12341 8938 12388 8940
rect 12296 8936 12388 8938
rect 12296 8880 12346 8936
rect 12296 8878 12388 8880
rect 12341 8876 12388 8878
rect 12452 8876 12458 8940
rect 12341 8875 12407 8876
rect 4337 8802 4403 8805
rect 8017 8802 8083 8805
rect 4337 8800 8083 8802
rect 4337 8744 4342 8800
rect 4398 8744 8022 8800
rect 8078 8744 8083 8800
rect 4337 8742 8083 8744
rect 4337 8739 4403 8742
rect 8017 8739 8083 8742
rect 11237 8802 11303 8805
rect 12157 8802 12223 8805
rect 11237 8800 12223 8802
rect 11237 8744 11242 8800
rect 11298 8744 12162 8800
rect 12218 8744 12223 8800
rect 11237 8742 12223 8744
rect 11237 8739 11303 8742
rect 12157 8739 12223 8742
rect 12341 8802 12407 8805
rect 13077 8802 13143 8805
rect 12341 8800 13143 8802
rect 12341 8744 12346 8800
rect 12402 8744 13082 8800
rect 13138 8744 13143 8800
rect 12341 8742 13143 8744
rect 12341 8739 12407 8742
rect 13077 8739 13143 8742
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 9765 8666 9831 8669
rect 12893 8666 12959 8669
rect 9765 8664 12959 8666
rect 9765 8608 9770 8664
rect 9826 8608 12898 8664
rect 12954 8608 12959 8664
rect 9765 8606 12959 8608
rect 9765 8603 9831 8606
rect 12893 8603 12959 8606
rect 5073 8530 5139 8533
rect 14457 8530 14523 8533
rect 5073 8528 14523 8530
rect 5073 8472 5078 8528
rect 5134 8472 14462 8528
rect 14518 8472 14523 8528
rect 5073 8470 14523 8472
rect 5073 8467 5139 8470
rect 14457 8467 14523 8470
rect 0 8394 800 8424
rect 3233 8394 3299 8397
rect 0 8392 3299 8394
rect 0 8336 3238 8392
rect 3294 8336 3299 8392
rect 0 8334 3299 8336
rect 0 8304 800 8334
rect 3233 8331 3299 8334
rect 3877 8396 3943 8397
rect 3877 8392 3924 8396
rect 3988 8394 3994 8396
rect 7833 8394 7899 8397
rect 9489 8394 9555 8397
rect 3877 8336 3882 8392
rect 3877 8332 3924 8336
rect 3988 8334 4034 8394
rect 7833 8392 9555 8394
rect 7833 8336 7838 8392
rect 7894 8336 9494 8392
rect 9550 8336 9555 8392
rect 7833 8334 9555 8336
rect 3988 8332 3994 8334
rect 3877 8331 3943 8332
rect 7833 8331 7899 8334
rect 9489 8331 9555 8334
rect 10133 8394 10199 8397
rect 10358 8394 10364 8396
rect 10133 8392 10364 8394
rect 10133 8336 10138 8392
rect 10194 8336 10364 8392
rect 10133 8334 10364 8336
rect 10133 8331 10199 8334
rect 10358 8332 10364 8334
rect 10428 8332 10434 8396
rect 11789 8394 11855 8397
rect 10550 8392 11855 8394
rect 10550 8336 11794 8392
rect 11850 8336 11855 8392
rect 10550 8334 11855 8336
rect 3325 8258 3391 8261
rect 5533 8258 5599 8261
rect 3325 8256 5599 8258
rect 3325 8200 3330 8256
rect 3386 8200 5538 8256
rect 5594 8200 5599 8256
rect 3325 8198 5599 8200
rect 3325 8195 3391 8198
rect 5533 8195 5599 8198
rect 6269 8258 6335 8261
rect 9121 8258 9187 8261
rect 6269 8256 9187 8258
rect 6269 8200 6274 8256
rect 6330 8200 9126 8256
rect 9182 8200 9187 8256
rect 6269 8198 9187 8200
rect 6269 8195 6335 8198
rect 9121 8195 9187 8198
rect 9765 8258 9831 8261
rect 10358 8258 10364 8260
rect 9765 8256 10364 8258
rect 9765 8200 9770 8256
rect 9826 8200 10364 8256
rect 9765 8198 10364 8200
rect 9765 8195 9831 8198
rect 10358 8196 10364 8198
rect 10428 8196 10434 8260
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 9806 8122 9812 8124
rect 6272 8062 9812 8122
rect 1945 7986 2011 7989
rect 6272 7986 6332 8062
rect 9806 8060 9812 8062
rect 9876 8060 9882 8124
rect 10225 8122 10291 8125
rect 10550 8122 10610 8334
rect 11789 8331 11855 8334
rect 12065 8394 12131 8397
rect 12893 8394 12959 8397
rect 12065 8392 12959 8394
rect 12065 8336 12070 8392
rect 12126 8336 12898 8392
rect 12954 8336 12959 8392
rect 12065 8334 12959 8336
rect 12065 8331 12131 8334
rect 12893 8331 12959 8334
rect 11237 8260 11303 8261
rect 11237 8258 11284 8260
rect 11192 8256 11284 8258
rect 11192 8200 11242 8256
rect 11192 8198 11284 8200
rect 11237 8196 11284 8198
rect 11348 8196 11354 8260
rect 12014 8196 12020 8260
rect 12084 8258 12090 8260
rect 12433 8258 12499 8261
rect 12084 8256 12499 8258
rect 12084 8200 12438 8256
rect 12494 8200 12499 8256
rect 12084 8198 12499 8200
rect 12084 8196 12090 8198
rect 11237 8195 11303 8196
rect 12433 8195 12499 8198
rect 15193 8258 15259 8261
rect 15193 8256 15394 8258
rect 15193 8200 15198 8256
rect 15254 8200 15394 8256
rect 15193 8198 15394 8200
rect 15193 8195 15259 8198
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 10225 8120 10610 8122
rect 10225 8064 10230 8120
rect 10286 8064 10610 8120
rect 10225 8062 10610 8064
rect 11237 8122 11303 8125
rect 12382 8122 12388 8124
rect 11237 8120 12388 8122
rect 11237 8064 11242 8120
rect 11298 8064 12388 8120
rect 11237 8062 12388 8064
rect 10225 8059 10291 8062
rect 11237 8059 11303 8062
rect 12382 8060 12388 8062
rect 12452 8060 12458 8124
rect 12985 8122 13051 8125
rect 15334 8122 15394 8198
rect 12985 8120 15394 8122
rect 12985 8064 12990 8120
rect 13046 8064 15394 8120
rect 12985 8062 15394 8064
rect 12985 8059 13051 8062
rect 1945 7984 6332 7986
rect 1945 7928 1950 7984
rect 2006 7928 6332 7984
rect 1945 7926 6332 7928
rect 6637 7986 6703 7989
rect 12433 7986 12499 7989
rect 6637 7984 12499 7986
rect 6637 7928 6642 7984
rect 6698 7928 12438 7984
rect 12494 7928 12499 7984
rect 6637 7926 12499 7928
rect 1945 7923 2011 7926
rect 6637 7923 6703 7926
rect 12433 7923 12499 7926
rect 4429 7850 4495 7853
rect 12750 7850 12756 7852
rect 4429 7848 12756 7850
rect 4429 7792 4434 7848
rect 4490 7792 12756 7848
rect 4429 7790 12756 7792
rect 4429 7787 4495 7790
rect 12750 7788 12756 7790
rect 12820 7788 12826 7852
rect 8753 7714 8819 7717
rect 11329 7714 11395 7717
rect 11605 7714 11671 7717
rect 8753 7712 11671 7714
rect 8753 7656 8758 7712
rect 8814 7656 11334 7712
rect 11390 7656 11610 7712
rect 11666 7656 11671 7712
rect 8753 7654 11671 7656
rect 8753 7651 8819 7654
rect 11329 7651 11395 7654
rect 11605 7651 11671 7654
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 10501 7578 10567 7581
rect 11462 7578 11468 7580
rect 10501 7576 11468 7578
rect 10501 7520 10506 7576
rect 10562 7520 11468 7576
rect 10501 7518 11468 7520
rect 10501 7515 10567 7518
rect 11462 7516 11468 7518
rect 11532 7516 11538 7580
rect 0 7442 800 7472
rect 1669 7442 1735 7445
rect 0 7440 1735 7442
rect 0 7384 1674 7440
rect 1730 7384 1735 7440
rect 0 7382 1735 7384
rect 0 7352 800 7382
rect 1669 7379 1735 7382
rect 4654 7380 4660 7444
rect 4724 7442 4730 7444
rect 4797 7442 4863 7445
rect 12065 7442 12131 7445
rect 4724 7440 4863 7442
rect 4724 7384 4802 7440
rect 4858 7384 4863 7440
rect 4724 7382 4863 7384
rect 4724 7380 4730 7382
rect 4797 7379 4863 7382
rect 7054 7440 12131 7442
rect 7054 7384 12070 7440
rect 12126 7384 12131 7440
rect 7054 7382 12131 7384
rect 3233 7306 3299 7309
rect 7054 7306 7114 7382
rect 12065 7379 12131 7382
rect 3233 7304 7114 7306
rect 3233 7248 3238 7304
rect 3294 7248 7114 7304
rect 3233 7246 7114 7248
rect 7189 7306 7255 7309
rect 13629 7306 13695 7309
rect 7189 7304 13695 7306
rect 7189 7248 7194 7304
rect 7250 7248 13634 7304
rect 13690 7248 13695 7304
rect 7189 7246 13695 7248
rect 3233 7243 3299 7246
rect 7189 7243 7255 7246
rect 13629 7243 13695 7246
rect 9581 7170 9647 7173
rect 10041 7170 10107 7173
rect 10501 7170 10567 7173
rect 9540 7168 9828 7170
rect 9540 7112 9586 7168
rect 9642 7112 9828 7168
rect 9540 7110 9828 7112
rect 9581 7107 9647 7110
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 1853 7034 1919 7037
rect 4889 7034 4955 7037
rect 1853 7032 4955 7034
rect 1853 6976 1858 7032
rect 1914 6976 4894 7032
rect 4950 6976 4955 7032
rect 1853 6974 4955 6976
rect 1853 6971 1919 6974
rect 4889 6971 4955 6974
rect 7005 7034 7071 7037
rect 9397 7034 9463 7037
rect 7005 7032 9463 7034
rect 7005 6976 7010 7032
rect 7066 6976 9402 7032
rect 9458 6976 9463 7032
rect 7005 6974 9463 6976
rect 7005 6971 7071 6974
rect 9397 6971 9463 6974
rect 3785 6898 3851 6901
rect 5349 6898 5415 6901
rect 3785 6896 5415 6898
rect 3785 6840 3790 6896
rect 3846 6840 5354 6896
rect 5410 6840 5415 6896
rect 3785 6838 5415 6840
rect 3785 6835 3851 6838
rect 5349 6835 5415 6838
rect 5533 6898 5599 6901
rect 8845 6898 8911 6901
rect 5533 6896 8911 6898
rect 5533 6840 5538 6896
rect 5594 6840 8850 6896
rect 8906 6840 8911 6896
rect 5533 6838 8911 6840
rect 5533 6835 5599 6838
rect 8845 6835 8911 6838
rect 9622 6836 9628 6900
rect 9692 6898 9698 6900
rect 9768 6898 9828 7110
rect 10041 7168 10567 7170
rect 10041 7112 10046 7168
rect 10102 7112 10506 7168
rect 10562 7112 10567 7168
rect 10041 7110 10567 7112
rect 10041 7107 10107 7110
rect 10501 7107 10567 7110
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 12566 6972 12572 7036
rect 12636 7034 12642 7036
rect 13629 7034 13695 7037
rect 12636 7032 13695 7034
rect 12636 6976 13634 7032
rect 13690 6976 13695 7032
rect 12636 6974 13695 6976
rect 12636 6972 12642 6974
rect 13629 6971 13695 6974
rect 9692 6838 9828 6898
rect 9692 6836 9698 6838
rect 10358 6836 10364 6900
rect 10428 6898 10434 6900
rect 12801 6898 12867 6901
rect 10428 6896 12867 6898
rect 10428 6840 12806 6896
rect 12862 6840 12867 6896
rect 10428 6838 12867 6840
rect 10428 6836 10434 6838
rect 12801 6835 12867 6838
rect 3233 6762 3299 6765
rect 12433 6762 12499 6765
rect 3233 6760 12499 6762
rect 3233 6704 3238 6760
rect 3294 6704 12438 6760
rect 12494 6704 12499 6760
rect 3233 6702 12499 6704
rect 3233 6699 3299 6702
rect 12433 6699 12499 6702
rect 4102 6564 4108 6628
rect 4172 6626 4178 6628
rect 5073 6626 5139 6629
rect 7833 6626 7899 6629
rect 4172 6624 7899 6626
rect 4172 6568 5078 6624
rect 5134 6568 7838 6624
rect 7894 6568 7899 6624
rect 4172 6566 7899 6568
rect 4172 6564 4178 6566
rect 5073 6563 5139 6566
rect 7833 6563 7899 6566
rect 9990 6564 9996 6628
rect 10060 6626 10066 6628
rect 10869 6626 10935 6629
rect 10060 6624 10935 6626
rect 10060 6568 10874 6624
rect 10930 6568 10935 6624
rect 10060 6566 10935 6568
rect 10060 6564 10066 6566
rect 10869 6563 10935 6566
rect 11053 6626 11119 6629
rect 12341 6626 12407 6629
rect 11053 6624 12407 6626
rect 11053 6568 11058 6624
rect 11114 6568 12346 6624
rect 12402 6568 12407 6624
rect 11053 6566 12407 6568
rect 11053 6563 11119 6566
rect 12341 6563 12407 6566
rect 3409 6560 3729 6561
rect 0 6490 800 6520
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 4061 6490 4127 6493
rect 8017 6490 8083 6493
rect 4061 6488 8083 6490
rect 4061 6432 4066 6488
rect 4122 6432 8022 6488
rect 8078 6432 8083 6488
rect 4061 6430 8083 6432
rect 4061 6427 4127 6430
rect 8017 6427 8083 6430
rect 9438 6428 9444 6492
rect 9508 6490 9514 6492
rect 9857 6490 9923 6493
rect 9508 6488 9923 6490
rect 9508 6432 9862 6488
rect 9918 6432 9923 6488
rect 9508 6430 9923 6432
rect 9508 6428 9514 6430
rect 9857 6427 9923 6430
rect 10225 6490 10291 6493
rect 11421 6490 11487 6493
rect 10225 6488 11487 6490
rect 10225 6432 10230 6488
rect 10286 6432 11426 6488
rect 11482 6432 11487 6488
rect 10225 6430 11487 6432
rect 10225 6427 10291 6430
rect 11421 6427 11487 6430
rect 1669 6354 1735 6357
rect 14641 6354 14707 6357
rect 1669 6352 14707 6354
rect 1669 6296 1674 6352
rect 1730 6296 14646 6352
rect 14702 6296 14707 6352
rect 1669 6294 14707 6296
rect 1669 6291 1735 6294
rect 14641 6291 14707 6294
rect 1117 6218 1183 6221
rect 15009 6218 15075 6221
rect 1117 6216 15075 6218
rect 1117 6160 1122 6216
rect 1178 6160 15014 6216
rect 15070 6160 15075 6216
rect 1117 6158 15075 6160
rect 1117 6155 1183 6158
rect 15009 6155 15075 6158
rect 8477 6082 8543 6085
rect 8753 6082 8819 6085
rect 8477 6080 8819 6082
rect 8477 6024 8482 6080
rect 8538 6024 8758 6080
rect 8814 6024 8819 6080
rect 8477 6022 8819 6024
rect 8477 6019 8543 6022
rect 8753 6019 8819 6022
rect 9029 6082 9095 6085
rect 10501 6082 10567 6085
rect 9029 6080 10567 6082
rect 9029 6024 9034 6080
rect 9090 6024 10506 6080
rect 10562 6024 10567 6080
rect 9029 6022 10567 6024
rect 9029 6019 9095 6022
rect 10501 6019 10567 6022
rect 11329 6082 11395 6085
rect 12341 6082 12407 6085
rect 11329 6080 12407 6082
rect 11329 6024 11334 6080
rect 11390 6024 12346 6080
rect 12402 6024 12407 6080
rect 11329 6022 12407 6024
rect 11329 6019 11395 6022
rect 12341 6019 12407 6022
rect 12750 6020 12756 6084
rect 12820 6082 12826 6084
rect 13445 6082 13511 6085
rect 12820 6080 13511 6082
rect 12820 6024 13450 6080
rect 13506 6024 13511 6080
rect 12820 6022 13511 6024
rect 12820 6020 12826 6022
rect 13445 6019 13511 6022
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 11830 5884 11836 5948
rect 11900 5946 11906 5948
rect 13261 5946 13327 5949
rect 11900 5944 13327 5946
rect 11900 5888 13266 5944
rect 13322 5888 13327 5944
rect 11900 5886 13327 5888
rect 11900 5884 11906 5886
rect 13261 5883 13327 5886
rect 5073 5810 5139 5813
rect 7281 5810 7347 5813
rect 14181 5810 14247 5813
rect 5073 5808 7347 5810
rect 5073 5752 5078 5808
rect 5134 5752 7286 5808
rect 7342 5752 7347 5808
rect 5073 5750 7347 5752
rect 5073 5747 5139 5750
rect 7281 5747 7347 5750
rect 7606 5808 14247 5810
rect 7606 5752 14186 5808
rect 14242 5752 14247 5808
rect 7606 5750 14247 5752
rect 1577 5674 1643 5677
rect 7606 5674 7666 5750
rect 14181 5747 14247 5750
rect 1577 5672 7666 5674
rect 1577 5616 1582 5672
rect 1638 5616 7666 5672
rect 1577 5614 7666 5616
rect 7833 5674 7899 5677
rect 9121 5674 9187 5677
rect 9622 5674 9628 5676
rect 7833 5672 8816 5674
rect 7833 5616 7838 5672
rect 7894 5616 8816 5672
rect 7833 5614 8816 5616
rect 1577 5611 1643 5614
rect 7833 5611 7899 5614
rect 5257 5538 5323 5541
rect 8201 5538 8267 5541
rect 5257 5536 8267 5538
rect 5257 5480 5262 5536
rect 5318 5480 8206 5536
rect 8262 5480 8267 5536
rect 5257 5478 8267 5480
rect 8756 5538 8816 5614
rect 9121 5672 9628 5674
rect 9121 5616 9126 5672
rect 9182 5616 9628 5672
rect 9121 5614 9628 5616
rect 9121 5611 9187 5614
rect 9622 5612 9628 5614
rect 9692 5612 9698 5676
rect 10174 5612 10180 5676
rect 10244 5674 10250 5676
rect 12198 5674 12204 5676
rect 10244 5614 12204 5674
rect 10244 5612 10250 5614
rect 12198 5612 12204 5614
rect 12268 5612 12274 5676
rect 13813 5674 13879 5677
rect 13126 5672 13879 5674
rect 13126 5616 13818 5672
rect 13874 5616 13879 5672
rect 13126 5614 13879 5616
rect 9581 5538 9647 5541
rect 13126 5538 13186 5614
rect 13813 5611 13879 5614
rect 8756 5536 13186 5538
rect 8756 5480 9586 5536
rect 9642 5480 13186 5536
rect 8756 5478 13186 5480
rect 5257 5475 5323 5478
rect 8201 5475 8267 5478
rect 9581 5475 9647 5478
rect 13854 5476 13860 5540
rect 13924 5538 13930 5540
rect 13997 5538 14063 5541
rect 13924 5536 14063 5538
rect 13924 5480 14002 5536
rect 14058 5480 14063 5536
rect 13924 5478 14063 5480
rect 13924 5476 13930 5478
rect 13997 5475 14063 5478
rect 3409 5472 3729 5473
rect 0 5402 800 5432
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 4245 5402 4311 5405
rect 9581 5402 9647 5405
rect 10961 5402 11027 5405
rect 0 5342 3296 5402
rect 0 5312 800 5342
rect 3236 5266 3296 5342
rect 4245 5400 8218 5402
rect 4245 5344 4250 5400
rect 4306 5344 8218 5400
rect 4245 5342 8218 5344
rect 4245 5339 4311 5342
rect 7281 5266 7347 5269
rect 3236 5264 7347 5266
rect 3236 5208 7286 5264
rect 7342 5208 7347 5264
rect 3236 5206 7347 5208
rect 7281 5203 7347 5206
rect 7465 5266 7531 5269
rect 8017 5266 8083 5269
rect 7465 5264 8083 5266
rect 7465 5208 7470 5264
rect 7526 5208 8022 5264
rect 8078 5208 8083 5264
rect 7465 5206 8083 5208
rect 8158 5266 8218 5342
rect 9581 5400 11027 5402
rect 9581 5344 9586 5400
rect 9642 5344 10966 5400
rect 11022 5344 11027 5400
rect 9581 5342 11027 5344
rect 9581 5339 9647 5342
rect 10961 5339 11027 5342
rect 12198 5340 12204 5404
rect 12268 5402 12274 5404
rect 12985 5402 13051 5405
rect 12268 5400 13051 5402
rect 12268 5344 12990 5400
rect 13046 5344 13051 5400
rect 12268 5342 13051 5344
rect 12268 5340 12274 5342
rect 12985 5339 13051 5342
rect 10225 5266 10291 5269
rect 8158 5264 10291 5266
rect 8158 5208 10230 5264
rect 10286 5208 10291 5264
rect 8158 5206 10291 5208
rect 7465 5203 7531 5206
rect 8017 5203 8083 5206
rect 10225 5203 10291 5206
rect 10358 5204 10364 5268
rect 10428 5266 10434 5268
rect 11145 5266 11211 5269
rect 10428 5264 11211 5266
rect 10428 5208 11150 5264
rect 11206 5208 11211 5264
rect 10428 5206 11211 5208
rect 10428 5204 10434 5206
rect 11145 5203 11211 5206
rect 11329 5266 11395 5269
rect 12382 5266 12388 5268
rect 11329 5264 12388 5266
rect 11329 5208 11334 5264
rect 11390 5208 12388 5264
rect 11329 5206 12388 5208
rect 11329 5203 11395 5206
rect 12382 5204 12388 5206
rect 12452 5204 12458 5268
rect 749 5130 815 5133
rect 15009 5130 15075 5133
rect 749 5128 15075 5130
rect 749 5072 754 5128
rect 810 5072 15014 5128
rect 15070 5072 15075 5128
rect 749 5070 15075 5072
rect 749 5067 815 5070
rect 15009 5067 15075 5070
rect 2589 4994 2655 4997
rect 3601 4994 3667 4997
rect 2589 4992 3667 4994
rect 2589 4936 2594 4992
rect 2650 4936 3606 4992
rect 3662 4936 3667 4992
rect 2589 4934 3667 4936
rect 2589 4931 2655 4934
rect 3601 4931 3667 4934
rect 4153 4994 4219 4997
rect 5533 4994 5599 4997
rect 4153 4992 5599 4994
rect 4153 4936 4158 4992
rect 4214 4936 5538 4992
rect 5594 4936 5599 4992
rect 4153 4934 5599 4936
rect 4153 4931 4219 4934
rect 5533 4931 5599 4934
rect 8017 4994 8083 4997
rect 9857 4994 9923 4997
rect 8017 4992 9923 4994
rect 8017 4936 8022 4992
rect 8078 4936 9862 4992
rect 9918 4936 9923 4992
rect 8017 4934 9923 4936
rect 8017 4931 8083 4934
rect 9857 4931 9923 4934
rect 10133 4994 10199 4997
rect 10358 4994 10364 4996
rect 10133 4992 10364 4994
rect 10133 4936 10138 4992
rect 10194 4936 10364 4992
rect 10133 4934 10364 4936
rect 10133 4931 10199 4934
rect 10358 4932 10364 4934
rect 10428 4932 10434 4996
rect 11462 4932 11468 4996
rect 11532 4994 11538 4996
rect 12341 4994 12407 4997
rect 11532 4992 12407 4994
rect 11532 4936 12346 4992
rect 12402 4936 12407 4992
rect 11532 4934 12407 4936
rect 11532 4932 11538 4934
rect 12341 4931 12407 4934
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 1945 4858 2011 4861
rect 4245 4858 4311 4861
rect 4613 4858 4679 4861
rect 1945 4856 4679 4858
rect 1945 4800 1950 4856
rect 2006 4800 4250 4856
rect 4306 4800 4618 4856
rect 4674 4800 4679 4856
rect 1945 4798 4679 4800
rect 1945 4795 2011 4798
rect 4245 4795 4311 4798
rect 4613 4795 4679 4798
rect 6637 4858 6703 4861
rect 10501 4858 10567 4861
rect 13721 4860 13787 4861
rect 6637 4856 10567 4858
rect 6637 4800 6642 4856
rect 6698 4800 10506 4856
rect 10562 4800 10567 4856
rect 6637 4798 10567 4800
rect 6637 4795 6703 4798
rect 10501 4795 10567 4798
rect 13670 4796 13676 4860
rect 13740 4858 13787 4860
rect 13740 4856 13832 4858
rect 13782 4800 13832 4856
rect 13740 4798 13832 4800
rect 13740 4796 13787 4798
rect 13721 4795 13787 4796
rect 381 4722 447 4725
rect 3049 4722 3115 4725
rect 4429 4722 4495 4725
rect 381 4720 1042 4722
rect 381 4664 386 4720
rect 442 4664 1042 4720
rect 381 4662 1042 4664
rect 381 4659 447 4662
rect 982 4586 1042 4662
rect 3049 4720 4495 4722
rect 3049 4664 3054 4720
rect 3110 4664 4434 4720
rect 4490 4664 4495 4720
rect 3049 4662 4495 4664
rect 3049 4659 3115 4662
rect 4429 4659 4495 4662
rect 4797 4722 4863 4725
rect 5257 4722 5323 4725
rect 4797 4720 5323 4722
rect 4797 4664 4802 4720
rect 4858 4664 5262 4720
rect 5318 4664 5323 4720
rect 4797 4662 5323 4664
rect 4797 4659 4863 4662
rect 5257 4659 5323 4662
rect 5717 4722 5783 4725
rect 11421 4722 11487 4725
rect 5717 4720 11487 4722
rect 5717 4664 5722 4720
rect 5778 4664 11426 4720
rect 11482 4664 11487 4720
rect 5717 4662 11487 4664
rect 5717 4659 5783 4662
rect 11421 4659 11487 4662
rect 14641 4586 14707 4589
rect 982 4584 14707 4586
rect 982 4528 14646 4584
rect 14702 4528 14707 4584
rect 982 4526 14707 4528
rect 14641 4523 14707 4526
rect 0 4450 800 4480
rect 1393 4450 1459 4453
rect 0 4448 1459 4450
rect 0 4392 1398 4448
rect 1454 4392 1459 4448
rect 0 4390 1459 4392
rect 0 4360 800 4390
rect 1393 4387 1459 4390
rect 5257 4450 5323 4453
rect 5390 4450 5396 4452
rect 5257 4448 5396 4450
rect 5257 4392 5262 4448
rect 5318 4392 5396 4448
rect 5257 4390 5396 4392
rect 5257 4387 5323 4390
rect 5390 4388 5396 4390
rect 5460 4388 5466 4452
rect 5717 4450 5783 4453
rect 6177 4450 6243 4453
rect 5717 4448 6243 4450
rect 5717 4392 5722 4448
rect 5778 4392 6182 4448
rect 6238 4392 6243 4448
rect 5717 4390 6243 4392
rect 5717 4387 5783 4390
rect 6177 4387 6243 4390
rect 9489 4450 9555 4453
rect 12525 4450 12591 4453
rect 9489 4448 12591 4450
rect 9489 4392 9494 4448
rect 9550 4392 12530 4448
rect 12586 4392 12591 4448
rect 9489 4390 12591 4392
rect 9489 4387 9555 4390
rect 12525 4387 12591 4390
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 2129 4314 2195 4317
rect 2086 4312 2195 4314
rect 2086 4256 2134 4312
rect 2190 4256 2195 4312
rect 2086 4251 2195 4256
rect 3877 4314 3943 4317
rect 3877 4312 7482 4314
rect 3877 4256 3882 4312
rect 3938 4256 7482 4312
rect 3877 4254 7482 4256
rect 3877 4251 3943 4254
rect 2086 4042 2146 4251
rect 4061 4180 4127 4181
rect 4061 4178 4108 4180
rect 4016 4176 4108 4178
rect 4016 4120 4066 4176
rect 4016 4118 4108 4120
rect 4061 4116 4108 4118
rect 4172 4116 4178 4180
rect 4245 4178 4311 4181
rect 6913 4178 6979 4181
rect 4245 4176 6979 4178
rect 4245 4120 4250 4176
rect 4306 4120 6918 4176
rect 6974 4120 6979 4176
rect 4245 4118 6979 4120
rect 7422 4178 7482 4254
rect 9254 4252 9260 4316
rect 9324 4314 9330 4316
rect 9489 4314 9555 4317
rect 9324 4312 9555 4314
rect 9324 4256 9494 4312
rect 9550 4256 9555 4312
rect 9324 4254 9555 4256
rect 9324 4252 9330 4254
rect 9489 4251 9555 4254
rect 9622 4252 9628 4316
rect 9692 4314 9698 4316
rect 9857 4314 9923 4317
rect 10685 4314 10751 4317
rect 9692 4312 10751 4314
rect 9692 4256 9862 4312
rect 9918 4256 10690 4312
rect 10746 4256 10751 4312
rect 9692 4254 10751 4256
rect 9692 4252 9698 4254
rect 9857 4251 9923 4254
rect 10685 4251 10751 4254
rect 10961 4314 11027 4317
rect 11421 4314 11487 4317
rect 12801 4314 12867 4317
rect 13118 4314 13124 4316
rect 10961 4312 13124 4314
rect 10961 4256 10966 4312
rect 11022 4256 11426 4312
rect 11482 4256 12806 4312
rect 12862 4256 13124 4312
rect 10961 4254 13124 4256
rect 10961 4251 11027 4254
rect 11421 4251 11487 4254
rect 12801 4251 12867 4254
rect 13118 4252 13124 4254
rect 13188 4252 13194 4316
rect 9673 4178 9739 4181
rect 7422 4176 9739 4178
rect 7422 4120 9678 4176
rect 9734 4120 9739 4176
rect 7422 4118 9739 4120
rect 4061 4115 4127 4116
rect 4245 4115 4311 4118
rect 6913 4115 6979 4118
rect 9673 4115 9739 4118
rect 9990 4116 9996 4180
rect 10060 4178 10066 4180
rect 10133 4178 10199 4181
rect 10060 4176 10199 4178
rect 10060 4120 10138 4176
rect 10194 4120 10199 4176
rect 10060 4118 10199 4120
rect 10060 4116 10066 4118
rect 10133 4115 10199 4118
rect 10501 4178 10567 4181
rect 14273 4178 14339 4181
rect 10501 4176 14339 4178
rect 10501 4120 10506 4176
rect 10562 4120 14278 4176
rect 14334 4120 14339 4176
rect 10501 4118 14339 4120
rect 10501 4115 10567 4118
rect 14273 4115 14339 4118
rect 14733 4042 14799 4045
rect 2086 4040 14799 4042
rect 2086 3984 14738 4040
rect 14794 3984 14799 4040
rect 2086 3982 14799 3984
rect 14733 3979 14799 3982
rect 3325 3906 3391 3909
rect 5165 3906 5231 3909
rect 3325 3904 5231 3906
rect 3325 3848 3330 3904
rect 3386 3848 5170 3904
rect 5226 3848 5231 3904
rect 3325 3846 5231 3848
rect 3325 3843 3391 3846
rect 5165 3843 5231 3846
rect 7097 3906 7163 3909
rect 10501 3906 10567 3909
rect 7097 3904 10567 3906
rect 7097 3848 7102 3904
rect 7158 3848 10506 3904
rect 10562 3848 10567 3904
rect 7097 3846 10567 3848
rect 7097 3843 7163 3846
rect 10501 3843 10567 3846
rect 12934 3844 12940 3908
rect 13004 3906 13010 3908
rect 13721 3906 13787 3909
rect 13004 3904 13787 3906
rect 13004 3848 13726 3904
rect 13782 3848 13787 3904
rect 13004 3846 13787 3848
rect 13004 3844 13010 3846
rect 13721 3843 13787 3846
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 2037 3770 2103 3773
rect 4153 3770 4219 3773
rect 4654 3770 4660 3772
rect 2037 3768 4660 3770
rect 2037 3712 2042 3768
rect 2098 3712 4158 3768
rect 4214 3712 4660 3768
rect 2037 3710 4660 3712
rect 2037 3707 2103 3710
rect 4153 3707 4219 3710
rect 4654 3708 4660 3710
rect 4724 3708 4730 3772
rect 2681 3634 2747 3637
rect 13905 3634 13971 3637
rect 2681 3632 13971 3634
rect 2681 3576 2686 3632
rect 2742 3576 13910 3632
rect 13966 3576 13971 3632
rect 2681 3574 13971 3576
rect 2681 3571 2747 3574
rect 13905 3571 13971 3574
rect 0 3498 800 3528
rect 3141 3498 3207 3501
rect 0 3496 3207 3498
rect 0 3440 3146 3496
rect 3202 3440 3207 3496
rect 0 3438 3207 3440
rect 0 3408 800 3438
rect 3141 3435 3207 3438
rect 3325 3498 3391 3501
rect 14365 3498 14431 3501
rect 3325 3496 14431 3498
rect 3325 3440 3330 3496
rect 3386 3440 14370 3496
rect 14426 3440 14431 3496
rect 3325 3438 14431 3440
rect 3325 3435 3391 3438
rect 14365 3435 14431 3438
rect 3877 3362 3943 3365
rect 3877 3360 8264 3362
rect 3877 3304 3882 3360
rect 3938 3304 8264 3360
rect 3877 3302 8264 3304
rect 3877 3299 3943 3302
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 7097 3226 7163 3229
rect 3926 3224 7163 3226
rect 3926 3168 7102 3224
rect 7158 3168 7163 3224
rect 3926 3166 7163 3168
rect 2773 3090 2839 3093
rect 3926 3090 3986 3166
rect 7097 3163 7163 3166
rect 2773 3088 3986 3090
rect 2773 3032 2778 3088
rect 2834 3032 3986 3088
rect 2773 3030 3986 3032
rect 4429 3090 4495 3093
rect 7925 3090 7991 3093
rect 4429 3088 7991 3090
rect 4429 3032 4434 3088
rect 4490 3032 7930 3088
rect 7986 3032 7991 3088
rect 4429 3030 7991 3032
rect 8204 3090 8264 3302
rect 9806 3300 9812 3364
rect 9876 3362 9882 3364
rect 10501 3362 10567 3365
rect 9876 3360 10567 3362
rect 9876 3304 10506 3360
rect 10562 3304 10567 3360
rect 9876 3302 10567 3304
rect 9876 3300 9882 3302
rect 10501 3299 10567 3302
rect 15101 3362 15167 3365
rect 16200 3362 17000 3392
rect 15101 3360 17000 3362
rect 15101 3304 15106 3360
rect 15162 3304 17000 3360
rect 15101 3302 17000 3304
rect 15101 3299 15167 3302
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 16200 3272 17000 3302
rect 13270 3231 13590 3232
rect 9213 3226 9279 3229
rect 12893 3226 12959 3229
rect 9213 3224 12959 3226
rect 9213 3168 9218 3224
rect 9274 3168 12898 3224
rect 12954 3168 12959 3224
rect 9213 3166 12959 3168
rect 9213 3163 9279 3166
rect 12893 3163 12959 3166
rect 10869 3090 10935 3093
rect 8204 3088 10935 3090
rect 8204 3032 10874 3088
rect 10930 3032 10935 3088
rect 8204 3030 10935 3032
rect 2773 3027 2839 3030
rect 4429 3027 4495 3030
rect 7925 3027 7991 3030
rect 10869 3027 10935 3030
rect 2405 2954 2471 2957
rect 9673 2954 9739 2957
rect 2405 2952 9739 2954
rect 2405 2896 2410 2952
rect 2466 2896 9678 2952
rect 9734 2896 9739 2952
rect 2405 2894 9739 2896
rect 2405 2891 2471 2894
rect 9673 2891 9739 2894
rect 11329 2954 11395 2957
rect 12249 2956 12315 2957
rect 12014 2954 12020 2956
rect 11329 2952 12020 2954
rect 11329 2896 11334 2952
rect 11390 2896 12020 2952
rect 11329 2894 12020 2896
rect 11329 2891 11395 2894
rect 12014 2892 12020 2894
rect 12084 2892 12090 2956
rect 12198 2954 12204 2956
rect 12158 2894 12204 2954
rect 12268 2952 12315 2956
rect 12310 2896 12315 2952
rect 12198 2892 12204 2894
rect 12268 2892 12315 2896
rect 12249 2891 12315 2892
rect 1485 2818 1551 2821
rect 10133 2818 10199 2821
rect 13813 2818 13879 2821
rect 1485 2816 5642 2818
rect 1485 2760 1490 2816
rect 1546 2760 5642 2816
rect 1485 2758 5642 2760
rect 1485 2755 1551 2758
rect 5582 2546 5642 2758
rect 6272 2816 10199 2818
rect 6272 2760 10138 2816
rect 10194 2760 10199 2816
rect 6272 2758 10199 2760
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 6272 2546 6332 2758
rect 10133 2755 10199 2758
rect 11286 2816 13879 2818
rect 11286 2760 13818 2816
rect 13874 2760 13879 2816
rect 11286 2758 13879 2760
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 10133 2682 10199 2685
rect 10542 2682 10548 2684
rect 10133 2680 10548 2682
rect 10133 2624 10138 2680
rect 10194 2624 10548 2680
rect 10133 2622 10548 2624
rect 10133 2619 10199 2622
rect 10542 2620 10548 2622
rect 10612 2620 10618 2684
rect 5582 2486 6332 2546
rect 9673 2546 9739 2549
rect 11286 2546 11346 2758
rect 13813 2755 13879 2758
rect 11973 2682 12039 2685
rect 12198 2682 12204 2684
rect 11973 2680 12204 2682
rect 11973 2624 11978 2680
rect 12034 2624 12204 2680
rect 11973 2622 12204 2624
rect 11973 2619 12039 2622
rect 12198 2620 12204 2622
rect 12268 2620 12274 2684
rect 9673 2544 11346 2546
rect 9673 2488 9678 2544
rect 9734 2488 11346 2544
rect 9673 2486 11346 2488
rect 9673 2483 9739 2486
rect 0 2410 800 2440
rect 1393 2410 1459 2413
rect 0 2408 1459 2410
rect 0 2352 1398 2408
rect 1454 2352 1459 2408
rect 0 2350 1459 2352
rect 0 2320 800 2350
rect 1393 2347 1459 2350
rect 5390 2348 5396 2412
rect 5460 2410 5466 2412
rect 6913 2410 6979 2413
rect 9765 2410 9831 2413
rect 5460 2408 9831 2410
rect 5460 2352 6918 2408
rect 6974 2352 9770 2408
rect 9826 2352 9831 2408
rect 5460 2350 9831 2352
rect 5460 2348 5466 2350
rect 6913 2347 6979 2350
rect 9765 2347 9831 2350
rect 10869 2410 10935 2413
rect 11830 2410 11836 2412
rect 10869 2408 11836 2410
rect 10869 2352 10874 2408
rect 10930 2352 11836 2408
rect 10869 2350 11836 2352
rect 10869 2347 10935 2350
rect 11830 2348 11836 2350
rect 11900 2348 11906 2412
rect 9949 2274 10015 2277
rect 10174 2274 10180 2276
rect 9949 2272 10180 2274
rect 9949 2216 9954 2272
rect 10010 2216 10180 2272
rect 9949 2214 10180 2216
rect 9949 2211 10015 2214
rect 10174 2212 10180 2214
rect 10244 2212 10250 2276
rect 11329 2274 11395 2277
rect 11646 2274 11652 2276
rect 11329 2272 11652 2274
rect 11329 2216 11334 2272
rect 11390 2216 11652 2272
rect 11329 2214 11652 2216
rect 11329 2211 11395 2214
rect 11646 2212 11652 2214
rect 11716 2212 11722 2276
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 11278 2076 11284 2140
rect 11348 2138 11354 2140
rect 12617 2138 12683 2141
rect 11348 2136 12683 2138
rect 11348 2080 12622 2136
rect 12678 2080 12683 2136
rect 11348 2078 12683 2080
rect 11348 2076 11354 2078
rect 12617 2075 12683 2078
rect 3509 2002 3575 2005
rect 3918 2002 3924 2004
rect 3509 2000 3924 2002
rect 3509 1944 3514 2000
rect 3570 1944 3924 2000
rect 3509 1942 3924 1944
rect 3509 1939 3575 1942
rect 3918 1940 3924 1942
rect 3988 1940 3994 2004
rect 0 1458 800 1488
rect 1853 1458 1919 1461
rect 0 1456 1919 1458
rect 0 1400 1858 1456
rect 1914 1400 1919 1456
rect 0 1398 1919 1400
rect 0 1368 800 1398
rect 1853 1395 1919 1398
rect 0 506 800 536
rect 2865 506 2931 509
rect 0 504 2931 506
rect 0 448 2870 504
rect 2926 448 2931 504
rect 0 446 2931 448
rect 0 416 800 446
rect 2865 443 2931 446
<< via3 >>
rect 9076 18532 9140 18596
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 9996 17308 10060 17372
rect 11284 17036 11348 17100
rect 12388 17036 12452 17100
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 9812 16552 9876 16556
rect 9812 16496 9826 16552
rect 9826 16496 9876 16552
rect 9812 16492 9876 16496
rect 10180 16492 10244 16556
rect 8892 16356 8956 16420
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 13124 15948 13188 16012
rect 7236 15812 7300 15876
rect 8892 15812 8956 15876
rect 10180 15812 10244 15876
rect 10548 15872 10612 15876
rect 10548 15816 10562 15872
rect 10562 15816 10612 15872
rect 10548 15812 10612 15816
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 12020 15736 12084 15740
rect 12020 15680 12070 15736
rect 12070 15680 12084 15736
rect 12020 15676 12084 15680
rect 5580 15404 5644 15468
rect 11836 15268 11900 15332
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 9628 15192 9692 15196
rect 9628 15136 9678 15192
rect 9678 15136 9692 15192
rect 9628 15132 9692 15136
rect 11468 15056 11532 15060
rect 11468 15000 11518 15056
rect 11518 15000 11532 15056
rect 11468 14996 11532 15000
rect 9260 14920 9324 14924
rect 9260 14864 9310 14920
rect 9310 14864 9324 14920
rect 9260 14860 9324 14864
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 10364 14648 10428 14652
rect 10364 14592 10378 14648
rect 10378 14592 10428 14648
rect 10364 14588 10428 14592
rect 12756 14512 12820 14516
rect 12756 14456 12806 14512
rect 12806 14456 12820 14512
rect 12756 14452 12820 14456
rect 10180 14180 10244 14244
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 9996 14044 10060 14108
rect 9628 13908 9692 13972
rect 9812 13968 9876 13972
rect 9812 13912 9826 13968
rect 9826 13912 9876 13968
rect 9812 13908 9876 13912
rect 12388 13696 12452 13700
rect 12388 13640 12438 13696
rect 12438 13640 12452 13696
rect 12388 13636 12452 13640
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 11652 13500 11716 13564
rect 12388 13500 12452 13564
rect 12204 13228 12268 13292
rect 9076 13092 9140 13156
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 10548 12956 10612 13020
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 12572 13016 12636 13020
rect 12572 12960 12586 13016
rect 12586 12960 12636 13016
rect 9444 12820 9508 12884
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 9260 12684 9324 12748
rect 12572 12956 12636 12960
rect 11284 12820 11348 12884
rect 12940 12820 13004 12884
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 13124 12548 13188 12612
rect 12020 12472 12084 12476
rect 12020 12416 12034 12472
rect 12034 12416 12084 12472
rect 12020 12412 12084 12416
rect 12756 12412 12820 12476
rect 12756 12276 12820 12340
rect 8892 12200 8956 12204
rect 8892 12144 8942 12200
rect 8942 12144 8956 12200
rect 8892 12140 8956 12144
rect 9628 12140 9692 12204
rect 9996 12140 10060 12204
rect 10364 12140 10428 12204
rect 11652 12004 11716 12068
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 7236 11868 7300 11932
rect 9260 11868 9324 11932
rect 12020 11868 12084 11932
rect 5580 11460 5644 11524
rect 11652 11596 11716 11660
rect 9260 11460 9324 11524
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 10364 11384 10428 11388
rect 10364 11328 10378 11384
rect 10378 11328 10428 11384
rect 10364 11324 10428 11328
rect 11652 11188 11716 11252
rect 13860 11188 13924 11252
rect 10180 10916 10244 10980
rect 13676 11052 13740 11116
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 8892 10644 8956 10708
rect 12204 10644 12268 10708
rect 12388 10432 12452 10436
rect 12388 10376 12438 10432
rect 12438 10376 12452 10432
rect 12388 10372 12452 10376
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 13124 10100 13188 10164
rect 10548 9828 10612 9892
rect 12572 9828 12636 9892
rect 12756 9828 12820 9892
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 8892 9556 8956 9620
rect 10180 9616 10244 9620
rect 10180 9560 10194 9616
rect 10194 9560 10244 9616
rect 10180 9556 10244 9560
rect 11284 9480 11348 9484
rect 11284 9424 11334 9480
rect 11334 9424 11348 9480
rect 11284 9420 11348 9424
rect 9444 9284 9508 9348
rect 11652 9284 11716 9348
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 9996 9148 10060 9212
rect 11652 9208 11716 9212
rect 11652 9152 11666 9208
rect 11666 9152 11716 9208
rect 11652 9148 11716 9152
rect 11468 9012 11532 9076
rect 12572 9556 12636 9620
rect 12020 8876 12084 8940
rect 12388 8936 12452 8940
rect 12388 8880 12402 8936
rect 12402 8880 12452 8936
rect 12388 8876 12452 8880
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 3924 8392 3988 8396
rect 3924 8336 3938 8392
rect 3938 8336 3988 8392
rect 3924 8332 3988 8336
rect 10364 8332 10428 8396
rect 10364 8196 10428 8260
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 9812 8060 9876 8124
rect 11284 8256 11348 8260
rect 11284 8200 11298 8256
rect 11298 8200 11348 8256
rect 11284 8196 11348 8200
rect 12020 8196 12084 8260
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 12388 8060 12452 8124
rect 12756 7788 12820 7852
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 11468 7516 11532 7580
rect 4660 7380 4724 7444
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 9628 6836 9692 6900
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 12572 6972 12636 7036
rect 10364 6836 10428 6900
rect 4108 6564 4172 6628
rect 9996 6564 10060 6628
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 9444 6428 9508 6492
rect 12756 6020 12820 6084
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 11836 5884 11900 5948
rect 9628 5612 9692 5676
rect 10180 5612 10244 5676
rect 12204 5612 12268 5676
rect 13860 5476 13924 5540
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 12204 5340 12268 5404
rect 10364 5204 10428 5268
rect 12388 5204 12452 5268
rect 10364 4932 10428 4996
rect 11468 4932 11532 4996
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 13676 4856 13740 4860
rect 13676 4800 13726 4856
rect 13726 4800 13740 4856
rect 13676 4796 13740 4800
rect 5396 4388 5460 4452
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 4108 4176 4172 4180
rect 4108 4120 4122 4176
rect 4122 4120 4172 4176
rect 4108 4116 4172 4120
rect 9260 4252 9324 4316
rect 9628 4252 9692 4316
rect 13124 4252 13188 4316
rect 9996 4116 10060 4180
rect 12940 3844 13004 3908
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 4660 3708 4724 3772
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 9812 3300 9876 3364
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 12020 2892 12084 2956
rect 12204 2952 12268 2956
rect 12204 2896 12254 2952
rect 12254 2896 12268 2952
rect 12204 2892 12268 2896
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 10548 2620 10612 2684
rect 12204 2620 12268 2684
rect 5396 2348 5460 2412
rect 11836 2348 11900 2412
rect 10180 2212 10244 2276
rect 11652 2212 11716 2276
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
rect 11284 2076 11348 2140
rect 3924 1940 3988 2004
<< metal4 >>
rect 9075 18596 9141 18597
rect 9075 18532 9076 18596
rect 9140 18532 9141 18596
rect 9075 18531 9141 18532
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 15264 3729 16288
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5874 15808 6195 16832
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 8891 16420 8957 16421
rect 8891 16356 8892 16420
rect 8956 16356 8957 16420
rect 8891 16355 8957 16356
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 7235 15876 7301 15877
rect 7235 15812 7236 15876
rect 7300 15812 7301 15876
rect 7235 15811 7301 15812
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5579 15468 5645 15469
rect 5579 15404 5580 15468
rect 5644 15404 5645 15468
rect 5579 15403 5645 15404
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 5582 11525 5642 15403
rect 5874 14720 6195 15744
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5579 11524 5645 11525
rect 5579 11460 5580 11524
rect 5644 11460 5645 11524
rect 5579 11459 5645 11460
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 5874 11456 6195 12480
rect 7238 11933 7298 15811
rect 8340 15264 8660 16288
rect 8894 15877 8954 16355
rect 8891 15876 8957 15877
rect 8891 15812 8892 15876
rect 8956 15812 8957 15876
rect 8891 15811 8957 15812
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8894 12205 8954 15811
rect 9078 13157 9138 18531
rect 9995 17372 10061 17373
rect 9995 17308 9996 17372
rect 10060 17308 10061 17372
rect 9995 17307 10061 17308
rect 9811 16556 9877 16557
rect 9811 16492 9812 16556
rect 9876 16492 9877 16556
rect 9811 16491 9877 16492
rect 9627 15196 9693 15197
rect 9627 15132 9628 15196
rect 9692 15132 9693 15196
rect 9627 15131 9693 15132
rect 9259 14924 9325 14925
rect 9259 14860 9260 14924
rect 9324 14860 9325 14924
rect 9259 14859 9325 14860
rect 9075 13156 9141 13157
rect 9075 13092 9076 13156
rect 9140 13092 9141 13156
rect 9075 13091 9141 13092
rect 9262 12749 9322 14859
rect 9630 13973 9690 15131
rect 9814 13973 9874 16491
rect 9998 14109 10058 17307
rect 10805 16896 11125 17456
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 11283 17100 11349 17101
rect 11283 17036 11284 17100
rect 11348 17036 11349 17100
rect 11283 17035 11349 17036
rect 12387 17100 12453 17101
rect 12387 17036 12388 17100
rect 12452 17036 12453 17100
rect 12387 17035 12453 17036
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10179 16556 10245 16557
rect 10179 16492 10180 16556
rect 10244 16492 10245 16556
rect 10179 16491 10245 16492
rect 10182 15877 10242 16491
rect 10179 15876 10245 15877
rect 10179 15812 10180 15876
rect 10244 15812 10245 15876
rect 10179 15811 10245 15812
rect 10547 15876 10613 15877
rect 10547 15812 10548 15876
rect 10612 15812 10613 15876
rect 10547 15811 10613 15812
rect 10363 14652 10429 14653
rect 10363 14588 10364 14652
rect 10428 14588 10429 14652
rect 10363 14587 10429 14588
rect 10179 14244 10245 14245
rect 10179 14180 10180 14244
rect 10244 14180 10245 14244
rect 10179 14179 10245 14180
rect 9995 14108 10061 14109
rect 9995 14044 9996 14108
rect 10060 14044 10061 14108
rect 9995 14043 10061 14044
rect 9627 13972 9693 13973
rect 9627 13908 9628 13972
rect 9692 13908 9693 13972
rect 9627 13907 9693 13908
rect 9811 13972 9877 13973
rect 9811 13908 9812 13972
rect 9876 13908 9877 13972
rect 9811 13907 9877 13908
rect 9443 12884 9509 12885
rect 9443 12820 9444 12884
rect 9508 12820 9509 12884
rect 9443 12819 9509 12820
rect 9259 12748 9325 12749
rect 9259 12684 9260 12748
rect 9324 12684 9325 12748
rect 9259 12683 9325 12684
rect 8891 12204 8957 12205
rect 8891 12140 8892 12204
rect 8956 12140 8957 12204
rect 8891 12139 8957 12140
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 7235 11932 7301 11933
rect 7235 11868 7236 11932
rect 7300 11868 7301 11932
rect 7235 11867 7301 11868
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 3923 8396 3989 8397
rect 3923 8332 3924 8396
rect 3988 8332 3989 8396
rect 3923 8331 3989 8332
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 3926 2005 3986 8331
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 4659 7444 4725 7445
rect 4659 7380 4660 7444
rect 4724 7380 4725 7444
rect 4659 7379 4725 7380
rect 4107 6628 4173 6629
rect 4107 6564 4108 6628
rect 4172 6564 4173 6628
rect 4107 6563 4173 6564
rect 4110 4181 4170 6563
rect 4107 4180 4173 4181
rect 4107 4116 4108 4180
rect 4172 4116 4173 4180
rect 4107 4115 4173 4116
rect 4662 3773 4722 7379
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5395 4452 5461 4453
rect 5395 4388 5396 4452
rect 5460 4388 5461 4452
rect 5395 4387 5461 4388
rect 4659 3772 4725 3773
rect 4659 3708 4660 3772
rect 4724 3708 4725 3772
rect 4659 3707 4725 3708
rect 5398 2413 5458 4387
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5395 2412 5461 2413
rect 5395 2348 5396 2412
rect 5460 2348 5461 2412
rect 5395 2347 5461 2348
rect 5874 2128 6195 2688
rect 8340 10912 8660 11936
rect 9259 11932 9325 11933
rect 9259 11868 9260 11932
rect 9324 11868 9325 11932
rect 9259 11867 9325 11868
rect 9262 11525 9322 11867
rect 9259 11524 9325 11525
rect 9259 11460 9260 11524
rect 9324 11460 9325 11524
rect 9259 11459 9325 11460
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 8891 10708 8957 10709
rect 8891 10644 8892 10708
rect 8956 10644 8957 10708
rect 8891 10643 8957 10644
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 8894 9621 8954 10643
rect 8891 9620 8957 9621
rect 8891 9556 8892 9620
rect 8956 9556 8957 9620
rect 8891 9555 8957 9556
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 9262 4317 9322 11459
rect 9446 9349 9506 12819
rect 9630 12205 9690 13907
rect 9998 12205 10058 14043
rect 9627 12204 9693 12205
rect 9627 12140 9628 12204
rect 9692 12140 9693 12204
rect 9627 12139 9693 12140
rect 9995 12204 10061 12205
rect 9995 12140 9996 12204
rect 10060 12140 10061 12204
rect 9995 12139 10061 12140
rect 9443 9348 9509 9349
rect 9443 9284 9444 9348
rect 9508 9284 9509 9348
rect 9443 9283 9509 9284
rect 9446 6493 9506 9283
rect 9630 6901 9690 12139
rect 10182 10981 10242 14179
rect 10366 12205 10426 14587
rect 10550 13021 10610 15811
rect 10805 15808 11125 16832
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10547 13020 10613 13021
rect 10547 12956 10548 13020
rect 10612 12956 10613 13020
rect 10547 12955 10613 12956
rect 10805 12544 11125 13568
rect 11286 12885 11346 17035
rect 12019 15740 12085 15741
rect 12019 15676 12020 15740
rect 12084 15676 12085 15740
rect 12019 15675 12085 15676
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11467 15060 11533 15061
rect 11467 14996 11468 15060
rect 11532 14996 11533 15060
rect 11467 14995 11533 14996
rect 11283 12884 11349 12885
rect 11283 12820 11284 12884
rect 11348 12820 11349 12884
rect 11283 12819 11349 12820
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10363 12204 10429 12205
rect 10363 12140 10364 12204
rect 10428 12140 10429 12204
rect 10363 12139 10429 12140
rect 10805 11456 11125 12480
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10363 11388 10429 11389
rect 10363 11324 10364 11388
rect 10428 11324 10429 11388
rect 10363 11323 10429 11324
rect 10179 10980 10245 10981
rect 10179 10916 10180 10980
rect 10244 10916 10245 10980
rect 10179 10915 10245 10916
rect 10179 9620 10245 9621
rect 10179 9556 10180 9620
rect 10244 9556 10245 9620
rect 10179 9555 10245 9556
rect 9995 9212 10061 9213
rect 9995 9148 9996 9212
rect 10060 9148 10061 9212
rect 9995 9147 10061 9148
rect 9811 8124 9877 8125
rect 9811 8060 9812 8124
rect 9876 8060 9877 8124
rect 9811 8059 9877 8060
rect 9627 6900 9693 6901
rect 9627 6836 9628 6900
rect 9692 6836 9693 6900
rect 9627 6835 9693 6836
rect 9443 6492 9509 6493
rect 9443 6428 9444 6492
rect 9508 6428 9509 6492
rect 9443 6427 9509 6428
rect 9627 5676 9693 5677
rect 9627 5612 9628 5676
rect 9692 5612 9693 5676
rect 9627 5611 9693 5612
rect 9630 4317 9690 5611
rect 9259 4316 9325 4317
rect 9259 4252 9260 4316
rect 9324 4252 9325 4316
rect 9259 4251 9325 4252
rect 9627 4316 9693 4317
rect 9627 4252 9628 4316
rect 9692 4252 9693 4316
rect 9627 4251 9693 4252
rect 9814 3365 9874 8059
rect 9998 6629 10058 9147
rect 9995 6628 10061 6629
rect 9995 6564 9996 6628
rect 10060 6564 10061 6628
rect 9995 6563 10061 6564
rect 9998 4181 10058 6563
rect 10182 5677 10242 9555
rect 10366 8397 10426 11323
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10547 9892 10613 9893
rect 10547 9828 10548 9892
rect 10612 9828 10613 9892
rect 10547 9827 10613 9828
rect 10363 8396 10429 8397
rect 10363 8332 10364 8396
rect 10428 8332 10429 8396
rect 10363 8331 10429 8332
rect 10363 8260 10429 8261
rect 10363 8196 10364 8260
rect 10428 8196 10429 8260
rect 10363 8195 10429 8196
rect 10366 6901 10426 8195
rect 10363 6900 10429 6901
rect 10363 6836 10364 6900
rect 10428 6836 10429 6900
rect 10363 6835 10429 6836
rect 10179 5676 10245 5677
rect 10179 5612 10180 5676
rect 10244 5612 10245 5676
rect 10179 5611 10245 5612
rect 9995 4180 10061 4181
rect 9995 4116 9996 4180
rect 10060 4116 10061 4180
rect 9995 4115 10061 4116
rect 9811 3364 9877 3365
rect 9811 3300 9812 3364
rect 9876 3300 9877 3364
rect 9811 3299 9877 3300
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 10182 2277 10242 5611
rect 10363 5268 10429 5269
rect 10363 5204 10364 5268
rect 10428 5204 10429 5268
rect 10363 5203 10429 5204
rect 10366 4997 10426 5203
rect 10363 4996 10429 4997
rect 10363 4932 10364 4996
rect 10428 4932 10429 4996
rect 10363 4931 10429 4932
rect 10550 2685 10610 9827
rect 10805 9280 11125 10304
rect 11283 9484 11349 9485
rect 11283 9420 11284 9484
rect 11348 9420 11349 9484
rect 11283 9419 11349 9420
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 11286 8261 11346 9419
rect 11470 9077 11530 14995
rect 11651 13564 11717 13565
rect 11651 13500 11652 13564
rect 11716 13500 11717 13564
rect 11651 13499 11717 13500
rect 11654 12069 11714 13499
rect 11651 12068 11717 12069
rect 11651 12004 11652 12068
rect 11716 12004 11717 12068
rect 11651 12003 11717 12004
rect 11654 11661 11714 12003
rect 11651 11660 11717 11661
rect 11651 11596 11652 11660
rect 11716 11596 11717 11660
rect 11651 11595 11717 11596
rect 11651 11252 11717 11253
rect 11651 11188 11652 11252
rect 11716 11188 11717 11252
rect 11651 11187 11717 11188
rect 11654 9349 11714 11187
rect 11651 9348 11717 9349
rect 11651 9284 11652 9348
rect 11716 9284 11717 9348
rect 11651 9283 11717 9284
rect 11651 9212 11717 9213
rect 11651 9148 11652 9212
rect 11716 9148 11717 9212
rect 11651 9147 11717 9148
rect 11467 9076 11533 9077
rect 11467 9012 11468 9076
rect 11532 9012 11533 9076
rect 11467 9011 11533 9012
rect 11283 8260 11349 8261
rect 11283 8196 11284 8260
rect 11348 8196 11349 8260
rect 11283 8195 11349 8196
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10547 2684 10613 2685
rect 10547 2620 10548 2684
rect 10612 2620 10613 2684
rect 10547 2619 10613 2620
rect 10179 2276 10245 2277
rect 10179 2212 10180 2276
rect 10244 2212 10245 2276
rect 10179 2211 10245 2212
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 2128 11125 2688
rect 11286 2141 11346 8195
rect 11467 7580 11533 7581
rect 11467 7516 11468 7580
rect 11532 7516 11533 7580
rect 11467 7515 11533 7516
rect 11470 4997 11530 7515
rect 11467 4996 11533 4997
rect 11467 4932 11468 4996
rect 11532 4932 11533 4996
rect 11467 4931 11533 4932
rect 11654 2277 11714 9147
rect 11838 5949 11898 15267
rect 12022 12477 12082 15675
rect 12390 13701 12450 17035
rect 13270 16352 13590 17376
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13123 16012 13189 16013
rect 13123 15948 13124 16012
rect 13188 15948 13189 16012
rect 13123 15947 13189 15948
rect 12755 14516 12821 14517
rect 12755 14452 12756 14516
rect 12820 14452 12821 14516
rect 12755 14451 12821 14452
rect 12387 13700 12453 13701
rect 12387 13636 12388 13700
rect 12452 13636 12453 13700
rect 12387 13635 12453 13636
rect 12387 13564 12453 13565
rect 12387 13500 12388 13564
rect 12452 13500 12453 13564
rect 12387 13499 12453 13500
rect 12203 13292 12269 13293
rect 12203 13228 12204 13292
rect 12268 13228 12269 13292
rect 12203 13227 12269 13228
rect 12019 12476 12085 12477
rect 12019 12412 12020 12476
rect 12084 12412 12085 12476
rect 12019 12411 12085 12412
rect 12019 11932 12085 11933
rect 12019 11868 12020 11932
rect 12084 11868 12085 11932
rect 12019 11867 12085 11868
rect 12022 8941 12082 11867
rect 12206 10709 12266 13227
rect 12203 10708 12269 10709
rect 12203 10644 12204 10708
rect 12268 10644 12269 10708
rect 12203 10643 12269 10644
rect 12390 10437 12450 13499
rect 12571 13020 12637 13021
rect 12571 12956 12572 13020
rect 12636 12956 12637 13020
rect 12571 12955 12637 12956
rect 12387 10436 12453 10437
rect 12387 10372 12388 10436
rect 12452 10372 12453 10436
rect 12387 10371 12453 10372
rect 12574 9893 12634 12955
rect 12758 12477 12818 14451
rect 12939 12884 13005 12885
rect 12939 12820 12940 12884
rect 13004 12820 13005 12884
rect 12939 12819 13005 12820
rect 12755 12476 12821 12477
rect 12755 12412 12756 12476
rect 12820 12412 12821 12476
rect 12755 12411 12821 12412
rect 12755 12340 12821 12341
rect 12755 12276 12756 12340
rect 12820 12276 12821 12340
rect 12755 12275 12821 12276
rect 12758 9893 12818 12275
rect 12571 9892 12637 9893
rect 12571 9828 12572 9892
rect 12636 9828 12637 9892
rect 12571 9827 12637 9828
rect 12755 9892 12821 9893
rect 12755 9828 12756 9892
rect 12820 9828 12821 9892
rect 12755 9827 12821 9828
rect 12571 9620 12637 9621
rect 12571 9556 12572 9620
rect 12636 9556 12637 9620
rect 12571 9555 12637 9556
rect 12019 8940 12085 8941
rect 12019 8876 12020 8940
rect 12084 8876 12085 8940
rect 12019 8875 12085 8876
rect 12387 8940 12453 8941
rect 12387 8876 12388 8940
rect 12452 8876 12453 8940
rect 12387 8875 12453 8876
rect 12019 8260 12085 8261
rect 12019 8196 12020 8260
rect 12084 8196 12085 8260
rect 12019 8195 12085 8196
rect 11835 5948 11901 5949
rect 11835 5884 11836 5948
rect 11900 5884 11901 5948
rect 11835 5883 11901 5884
rect 11838 2413 11898 5883
rect 12022 2957 12082 8195
rect 12390 8125 12450 8875
rect 12387 8124 12453 8125
rect 12387 8060 12388 8124
rect 12452 8060 12453 8124
rect 12387 8059 12453 8060
rect 12203 5676 12269 5677
rect 12203 5612 12204 5676
rect 12268 5612 12269 5676
rect 12203 5611 12269 5612
rect 12206 5405 12266 5611
rect 12203 5404 12269 5405
rect 12203 5340 12204 5404
rect 12268 5340 12269 5404
rect 12203 5339 12269 5340
rect 12390 5269 12450 8059
rect 12574 7037 12634 9555
rect 12755 7852 12821 7853
rect 12755 7788 12756 7852
rect 12820 7788 12821 7852
rect 12755 7787 12821 7788
rect 12571 7036 12637 7037
rect 12571 6972 12572 7036
rect 12636 6972 12637 7036
rect 12571 6971 12637 6972
rect 12758 6085 12818 7787
rect 12755 6084 12821 6085
rect 12755 6020 12756 6084
rect 12820 6020 12821 6084
rect 12755 6019 12821 6020
rect 12387 5268 12453 5269
rect 12387 5204 12388 5268
rect 12452 5204 12453 5268
rect 12387 5203 12453 5204
rect 12942 3909 13002 12819
rect 13126 12613 13186 15947
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13123 12612 13189 12613
rect 13123 12548 13124 12612
rect 13188 12548 13189 12612
rect 13123 12547 13189 12548
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13859 11252 13925 11253
rect 13859 11188 13860 11252
rect 13924 11188 13925 11252
rect 13859 11187 13925 11188
rect 13675 11116 13741 11117
rect 13675 11052 13676 11116
rect 13740 11052 13741 11116
rect 13675 11051 13741 11052
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13123 10164 13189 10165
rect 13123 10100 13124 10164
rect 13188 10100 13189 10164
rect 13123 10099 13189 10100
rect 13126 4317 13186 10099
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13678 4861 13738 11051
rect 13862 5541 13922 11187
rect 13859 5540 13925 5541
rect 13859 5476 13860 5540
rect 13924 5476 13925 5540
rect 13859 5475 13925 5476
rect 13675 4860 13741 4861
rect 13675 4796 13676 4860
rect 13740 4796 13741 4860
rect 13675 4795 13741 4796
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13123 4316 13189 4317
rect 13123 4252 13124 4316
rect 13188 4252 13189 4316
rect 13123 4251 13189 4252
rect 12939 3908 13005 3909
rect 12939 3844 12940 3908
rect 13004 3844 13005 3908
rect 12939 3843 13005 3844
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 12019 2956 12085 2957
rect 12019 2892 12020 2956
rect 12084 2892 12085 2956
rect 12019 2891 12085 2892
rect 12203 2956 12269 2957
rect 12203 2892 12204 2956
rect 12268 2892 12269 2956
rect 12203 2891 12269 2892
rect 12206 2685 12266 2891
rect 12203 2684 12269 2685
rect 12203 2620 12204 2684
rect 12268 2620 12269 2684
rect 12203 2619 12269 2620
rect 11835 2412 11901 2413
rect 11835 2348 11836 2412
rect 11900 2348 11901 2412
rect 11835 2347 11901 2348
rect 11651 2276 11717 2277
rect 11651 2212 11652 2276
rect 11716 2212 11717 2276
rect 11651 2211 11717 2212
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 11283 2140 11349 2141
rect 11283 2076 11284 2140
rect 11348 2076 11349 2140
rect 13270 2128 13590 2144
rect 11283 2075 11349 2076
rect 3923 2004 3989 2005
rect 3923 1940 3924 2004
rect 3988 1940 3989 2004
rect 3923 1939 3989 1940
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608764397
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608764397
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608764397
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608764397
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1608764397
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1608764397
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 1608764397
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1608764397
transform 1 0 15456 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608764397
transform 1 0 13340 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1608764397
transform 1 0 12972 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_137
timestamp 1608764397
transform 1 0 13708 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_129
timestamp 1608764397
transform 1 0 12972 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_141
timestamp 1608764397
transform 1 0 14076 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608764397
transform 1 0 12604 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608764397
transform 1 0 12604 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608764397
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_122
timestamp 1608764397
transform 1 0 12328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608764397
transform 1 0 11868 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1608764397
transform 1 0 12236 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1608764397
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608764397
transform 1 0 11132 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608764397
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1608764397
transform 1 0 10764 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1608764397
transform 1 0 11500 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_106
timestamp 1608764397
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608764397
transform 1 0 10396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608764397
transform 1 0 10488 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 1608764397
transform 1 0 10120 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608764397
transform 1 0 9752 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1608764397
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608764397
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608764397
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608764397
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1608764397
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608764397
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608764397
transform 1 0 8832 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1608764397
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1608764397
transform 1 0 9200 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608764397
transform 1 0 8096 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1608764397
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1608764397
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1608764397
transform 1 0 7268 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1608764397
transform 1 0 8464 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1608764397
transform 1 0 7728 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_80
timestamp 1608764397
transform 1 0 8464 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608764397
transform 1 0 4968 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1608764397
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1608764397
transform 1 0 5244 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1608764397
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608764397
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 4968 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1608764397
transform 1 0 6072 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1608764397
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1608764397
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1608764397
transform 1 0 4048 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608764397
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608764397
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1608764397
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1608764397
transform 1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_26
timestamp 1608764397
transform 1 0 3496 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_30
timestamp 1608764397
transform 1 0 3864 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_38
timestamp 1608764397
transform 1 0 4600 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 2668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1608764397
transform 1 0 2944 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1608764397
transform 1 0 2576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1608764397
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1748 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_13
timestamp 1608764397
transform 1 0 2300 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_9
timestamp 1608764397
transform 1 0 1932 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608764397
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608764397
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1608764397
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1608764397
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608764397
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1608764397
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608764397
transform 1 0 13156 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608764397
transform 1 0 13892 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1608764397
transform 1 0 12788 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1608764397
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_143
timestamp 1608764397
transform 1 0 14260 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608764397
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608764397
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608764397
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_105
timestamp 1608764397
transform 1 0 10764 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1608764397
transform 1 0 11500 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1608764397
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608764397
transform 1 0 10396 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1608764397
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1608764397
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1608764397
transform 1 0 10028 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1608764397
transform 1 0 8004 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1608764397
transform 1 0 7636 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1608764397
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1608764397
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608764397
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_53
timestamp 1608764397
transform 1 0 5980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1608764397
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1608764397
transform 1 0 3956 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_23
timestamp 1608764397
transform 1 0 3220 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_40
timestamp 1608764397
transform 1 0 4784 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 2668 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1748 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608764397
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1608764397
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_13
timestamp 1608764397
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608764397
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608764397
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1608764397
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1608764397
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1608764397
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608764397
transform 1 0 13064 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1608764397
transform 1 0 12696 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_134
timestamp 1608764397
transform 1 0 13432 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608764397
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608764397
transform 1 0 11592 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608764397
transform 1 0 12328 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1608764397
transform 1 0 11224 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1608764397
transform 1 0 11960 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1608764397
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608764397
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1608764397
transform 1 0 8924 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1608764397
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608764397
transform 1 0 8556 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1608764397
transform 1 0 7360 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1608764397
transform 1 0 6992 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1608764397
transform 1 0 8188 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 5520 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp 1608764397
transform 1 0 5152 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1608764397
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608764397
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_22
timestamp 1608764397
transform 1 0 3128 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1608764397
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 2576 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1656 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608764397
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1608764397
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1608764397
transform 1 0 2208 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608764397
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_146
timestamp 1608764397
transform 1 0 14536 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_154
timestamp 1608764397
transform 1 0 15272 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608764397
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1608764397
transform 1 0 12788 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_134
timestamp 1608764397
transform 1 0 13432 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608764397
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1608764397
transform 1 0 11040 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608764397
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1608764397
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1608764397
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1608764397
transform 1 0 9844 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1608764397
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_104
timestamp 1608764397
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1608764397
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1608764397
transform 1 0 8280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608764397
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1608764397
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1608764397
transform 1 0 3680 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_24
timestamp 1608764397
transform 1 0 3312 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_37
timestamp 1608764397
transform 1 0 4508 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1564 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1608764397
transform 1 0 2484 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608764397
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1608764397
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1608764397
transform 1 0 2116 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608764397
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608764397
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1608764397
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608764397
transform 1 0 13524 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608764397
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608764397
transform 1 0 12788 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1608764397
transform 1 0 13156 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_138
timestamp 1608764397
transform 1 0 13800 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1608764397
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608764397
transform 1 0 12052 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1608764397
transform 1 0 10856 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1608764397
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_123
timestamp 1608764397
transform 1 0 12420 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1608764397
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608764397
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1608764397
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1608764397
transform 1 0 10488 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_63
timestamp 1608764397
transform 1 0 6900 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_83
timestamp 1608764397
transform 1 0 8740 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 5428 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1608764397
transform 1 0 5060 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1608764397
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608764397
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608764397
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1608764397
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1840 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1608764397
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608764397
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608764397
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1608764397
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1608764397
transform 1 0 2392 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1608764397
transform 1 0 14628 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608764397
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1608764397
transform 1 0 15180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608764397
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1608764397
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_139
timestamp 1608764397
transform 1 0 13892 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608764397
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1608764397
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608764397
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1608764397
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1608764397
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1608764397
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1608764397
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 8648 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1608764397
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608764397
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1608764397
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 3036 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1608764397
transform 1 0 4508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1608764397
transform 1 0 1840 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608764397
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1608764397
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1608764397
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_17
timestamp 1608764397
transform 1 0 2668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1608764397
transform 1 0 14536 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608764397
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608764397
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608764397
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1608764397
transform 1 0 15088 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_156
timestamp 1608764397
transform 1 0 15456 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1608764397
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1608764397
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1608764397
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608764397
transform 1 0 14444 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1608764397
transform 1 0 13248 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1608764397
transform 1 0 13616 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1608764397
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1608764397
transform 1 0 14168 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_128
timestamp 1608764397
transform 1 0 12880 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1608764397
transform 1 0 14076 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608764397
transform 1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1608764397
transform 1 0 10856 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1608764397
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1608764397
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608764397
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_111
timestamp 1608764397
transform 1 0 11316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1608764397
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1608764397
transform 1 0 11684 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1608764397
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1608764397
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608764397
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1608764397
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1608764397
transform 1 0 8924 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1608764397
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7452 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 8648 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1608764397
transform 1 0 8280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1608764397
transform 1 0 7084 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 5612 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608764397
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1608764397
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1608764397
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1608764397
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1608764397
transform 1 0 3680 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608764397
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1608764397
transform 1 0 3312 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1608764397
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608764397
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1608764397
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1608764397
transform 1 0 2484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_11
timestamp 1608764397
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1608764397
transform 1 0 2392 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1564 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608764397
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608764397
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1608764397
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1608764397
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608764397
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608764397
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1608764397
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1608764397
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608764397
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1608764397
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1608764397
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1608764397
transform 1 0 14076 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1608764397
transform 1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1608764397
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1608764397
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1608764397
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608764397
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_84
timestamp 1608764397
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608764397
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1608764397
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7360 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1608764397
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1608764397
transform 1 0 5152 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1608764397
transform 1 0 4324 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608764397
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608764397
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1608764397
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608764397
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1608764397
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1608764397
transform 1 0 2392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608764397
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608764397
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1608764397
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1608764397
transform 1 0 13616 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1608764397
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1608764397
transform 1 0 14444 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608764397
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1608764397
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608764397
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_111
timestamp 1608764397
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1608764397
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1608764397
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1608764397
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 8648 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1608764397
transform 1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608764397
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1608764397
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 3036 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_37
timestamp 1608764397
transform 1 0 4508 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1608764397
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608764397
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1608764397
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1608764397
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1608764397
transform 1 0 2668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608764397
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608764397
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1608764397
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1608764397
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608764397
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1608764397
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1608764397
transform 1 0 12880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1608764397
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1608764397
transform 1 0 10856 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1608764397
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1608764397
transform 1 0 11684 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608764397
transform 1 0 8924 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1608764397
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608764397
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1608764397
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1608764397
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 7084 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_81
timestamp 1608764397
transform 1 0 8556 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 5244 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_61
timestamp 1608764397
transform 1 0 6716 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1608764397
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608764397
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608764397
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1608764397
transform 1 0 4876 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608764397
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1608764397
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1608764397
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_14
timestamp 1608764397
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608764397
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608764397
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1608764397
transform 1 0 15180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1608764397
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1608764397
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1608764397
transform 1 0 14444 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1608764397
transform 1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1608764397
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608764397
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_111
timestamp 1608764397
transform 1 0 11316 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1608764397
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1608764397
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1608764397
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 8648 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1608764397
transform 1 0 8280 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 5244 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608764397
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 4968 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 3036 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1608764397
transform 1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_41
timestamp 1608764397
transform 1 0 4876 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1608764397
transform 1 0 1840 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608764397
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1608764397
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1608764397
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1608764397
transform 1 0 2668 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608764397
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608764397
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608764397
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608764397
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1608764397
transform 1 0 15180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1608764397
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1608764397
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608764397
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1608764397
transform 1 0 13616 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1608764397
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1608764397
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1608764397
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 1608764397
transform 1 0 12880 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1608764397
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1608764397
transform 1 0 10856 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1608764397
transform 1 0 11040 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1608764397
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1608764397
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608764397
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1608764397
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1608764397
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1608764397
transform 1 0 11684 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1608764397
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1608764397
transform 1 0 9844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608764397
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1608764397
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1608764397
transform 1 0 10672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1608764397
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1608764397
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1608764397
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7636 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1608764397
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1608764397
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_68
timestamp 1608764397
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 5888 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608764397
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1608764397
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 4416 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1608764397
transform 1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1608764397
transform 1 0 3220 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608764397
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608764397
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1608764397
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1608764397
transform 1 0 2392 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1608764397
transform 1 0 2760 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_11
timestamp 1608764397
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1608764397
transform 1 0 2392 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1564 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1608764397
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608764397
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608764397
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1608764397
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1608764397
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608764397
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608764397
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1608764397
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1608764397
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608764397
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1608764397
transform 1 0 13248 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1608764397
transform 1 0 12880 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1608764397
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1608764397
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1608764397
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1608764397
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1608764397
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608764397
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1608764397
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1608764397
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 7728 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 5888 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1608764397
transform 1 0 5520 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608764397
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608764397
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608764397
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1608764397
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1608764397
transform 1 0 2392 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608764397
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608764397
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1608764397
transform 1 0 15180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1608764397
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1608764397
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1608764397
transform 1 0 14444 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1608764397
transform 1 0 11040 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1608764397
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608764397
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1608764397
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608764397
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1608764397
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1608764397
transform 1 0 9476 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 1608764397
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1608764397
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1608764397
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608764397
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1608764397
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1608764397
transform 1 0 3680 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1608764397
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1608764397
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1564 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1608764397
transform 1 0 2484 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608764397
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1608764397
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1608764397
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608764397
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608764397
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1608764397
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1608764397
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608764397
transform 1 0 14444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1608764397
transform 1 0 13248 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1608764397
transform 1 0 12880 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1608764397
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1608764397
transform 1 0 10856 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1608764397
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1608764397
transform 1 0 11684 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1608764397
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608764397
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1608764397
transform 1 0 8924 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1608764397
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7452 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1608764397
transform 1 0 7084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 5612 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_45
timestamp 1608764397
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1608764397
transform 1 0 4416 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608764397
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608764397
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1608764397
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608764397
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1608764397
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1608764397
transform 1 0 2392 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608764397
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608764397
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1608764397
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1608764397
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1608764397
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1608764397
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608764397
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1608764397
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608764397
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1608764397
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1608764397
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1608764397
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1608764397
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1608764397
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608764397
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1608764397
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1608764397
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1608764397
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608764397
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1608764397
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1608764397
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1608764397
transform 1 0 2668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608764397
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608764397
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1608764397
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1608764397
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1608764397
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1608764397
transform 1 0 12696 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1608764397
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1608764397
transform 1 0 13524 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1608764397
transform 1 0 11500 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1608764397
transform 1 0 11132 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1608764397
transform 1 0 12328 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608764397
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1608764397
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1608764397
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7636 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1608764397
transform 1 0 7268 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 5796 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_47
timestamp 1608764397
transform 1 0 5428 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1608764397
transform 1 0 4600 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608764397
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608764397
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1608764397
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608764397
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1608764397
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1608764397
transform 1 0 2392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608764397
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608764397
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608764397
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608764397
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608764397
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1608764397
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1608764397
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1608764397
transform 1 0 13524 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1608764397
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1608764397
transform 1 0 13156 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1608764397
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1608764397
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1608764397
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608764397
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1608764397
transform 1 0 11132 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1608764397
transform 1 0 12328 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1608764397
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608764397
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp 1608764397
transform 1 0 10764 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_118
timestamp 1608764397
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1608764397
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1608764397
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1608764397
transform 1 0 8924 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1608764397
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608764397
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608764397
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1608764397
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1608764397
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7084 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_81
timestamp 1608764397
transform 1 0 8556 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1608764397
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 5244 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608764397
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_61
timestamp 1608764397
transform 1 0 6716 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1608764397
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1608764397
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608764397
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608764397
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1608764397
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1608764397
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1608764397
transform 1 0 2392 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1608764397
transform 1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1608764397
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608764397
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608764397
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1608764397
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1608764397
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1608764397
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608764397
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608764397
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1608764397
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1608764397
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1608764397
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1608764397
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608764397
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1608764397
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608764397
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_111
timestamp 1608764397
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1608764397
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1608764397
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1608764397
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 8648 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1608764397
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608764397
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1608764397
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 3036 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1608764397
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1608764397
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608764397
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1608764397
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1608764397
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1608764397
transform 1 0 2668 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608764397
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608764397
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1608764397
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1608764397
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608764397
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1608764397
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1608764397
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1608764397
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1608764397
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1608764397
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1608764397
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1608764397
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608764397
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1608764397
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1608764397
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 7268 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1608764397
transform 1 0 6900 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_83
timestamp 1608764397
transform 1 0 8740 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 5428 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_43
timestamp 1608764397
transform 1 0 5060 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1608764397
transform 1 0 4232 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608764397
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608764397
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1608764397
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1608764397
transform 1 0 2760 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1608764397
transform 1 0 1564 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608764397
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1608764397
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_14
timestamp 1608764397
transform 1 0 2392 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1608764397
transform 1 0 14536 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608764397
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_152
timestamp 1608764397
transform 1 0 15088 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_156
timestamp 1608764397
transform 1 0 15456 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1608764397
transform 1 0 13616 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1608764397
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1608764397
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608764397
transform 1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1608764397
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608764397
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_111
timestamp 1608764397
transform 1 0 11316 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1608764397
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1608764397
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1608764397
transform 1 0 10120 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 8648 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1608764397
transform 1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608764397
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1608764397
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764397
transform 1 0 4876 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1608764397
transform 1 0 3680 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1608764397
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1608764397
transform 1 0 4508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1608764397
transform 1 0 2484 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1564 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608764397
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1608764397
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1608764397
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608764397
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608764397
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1608764397
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1608764397
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 13248 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1608764397
transform 1 0 14260 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1608764397
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_138
timestamp 1608764397
transform 1 0 13800 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1608764397
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1608764397
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1608764397
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1608764397
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1608764397
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608764397
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9016 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1608764397
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1608764397
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 7176 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1608764397
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764397
transform 1 0 5336 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1608764397
transform 1 0 4968 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1608764397
transform 1 0 6808 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1608764397
transform 1 0 4140 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608764397
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608764397
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1608764397
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1608764397
transform 1 0 2760 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1608764397
transform 1 0 1564 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608764397
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1608764397
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1608764397
transform 1 0 2392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608764397
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608764397
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608764397
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608764397
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1608764397
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_149
timestamp 1608764397
transform 1 0 14812 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1608764397
transform 1 0 13892 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1608764397
transform 1 0 14260 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1608764397
transform 1 0 13340 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1608764397
transform 1 0 13156 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145
timestamp 1608764397
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1608764397
transform 1 0 12972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1608764397
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608764397
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1608764397
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608764397
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 12144 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116
timestamp 1608764397
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1608764397
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1608764397
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608764397
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1608764397
transform 1 0 11040 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1608764397
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1608764397
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1608764397
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608764397
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_right_ipin_0.prog_clk
timestamp 1608764397
transform 1 0 9292 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1608764397
transform 1 0 8924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1608764397
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1608764397
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 1608764397
transform 1 0 9476 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1608764397
transform 1 0 10672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1608764397
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1608764397
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1608764397
transform 1 0 8648 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1608764397
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1608764397
transform 1 0 8280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764397
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1608764397
transform 1 0 5612 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608764397
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608764397
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1608764397
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1608764397
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1608764397
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 4876 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1608764397
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1608764397
transform 1 0 4416 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608764397
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608764397
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1608764397
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1608764397
transform 1 0 3312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1608764397
transform 1 0 4508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608764397
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764397
transform 1 0 2116 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764397
transform 1 0 1564 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1608764397
transform 1 0 2484 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608764397
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608764397
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7
timestamp 1608764397
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1608764397
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1608764397
transform 1 0 2116 0 1 2720
box -38 -48 406 592
<< labels >>
rlabel metal3 s 16200 16600 17000 16720 4 Test_en_E_in
port 1 nsew
rlabel metal3 s 16200 9936 17000 10056 4 Test_en_E_out
port 2 nsew
rlabel metal2 s 3146 19200 3202 20000 4 Test_en_N_out
port 3 nsew
rlabel metal2 s 13726 0 13782 800 4 Test_en_S_in
port 4 nsew
rlabel metal3 s 0 17280 800 17400 4 Test_en_W_in
port 5 nsew
rlabel metal3 s 0 18368 800 18488 4 Test_en_W_out
port 6 nsew
rlabel metal3 s 0 416 800 536 4 ccff_head
port 7 nsew
rlabel metal3 s 16200 3272 17000 3392 4 ccff_tail
port 8 nsew
rlabel metal2 s 6918 0 6974 800 4 chany_bottom_in[0]
port 9 nsew
rlabel metal2 s 10322 0 10378 800 4 chany_bottom_in[10]
port 10 nsew
rlabel metal2 s 10598 0 10654 800 4 chany_bottom_in[11]
port 11 nsew
rlabel metal2 s 10966 0 11022 800 4 chany_bottom_in[12]
port 12 nsew
rlabel metal2 s 11334 0 11390 800 4 chany_bottom_in[13]
port 13 nsew
rlabel metal2 s 11610 0 11666 800 4 chany_bottom_in[14]
port 14 nsew
rlabel metal2 s 11978 0 12034 800 4 chany_bottom_in[15]
port 15 nsew
rlabel metal2 s 12346 0 12402 800 4 chany_bottom_in[16]
port 16 nsew
rlabel metal2 s 12622 0 12678 800 4 chany_bottom_in[17]
port 17 nsew
rlabel metal2 s 12990 0 13046 800 4 chany_bottom_in[18]
port 18 nsew
rlabel metal2 s 13358 0 13414 800 4 chany_bottom_in[19]
port 19 nsew
rlabel metal2 s 7194 0 7250 800 4 chany_bottom_in[1]
port 20 nsew
rlabel metal2 s 7562 0 7618 800 4 chany_bottom_in[2]
port 21 nsew
rlabel metal2 s 7930 0 7986 800 4 chany_bottom_in[3]
port 22 nsew
rlabel metal2 s 8206 0 8262 800 4 chany_bottom_in[4]
port 23 nsew
rlabel metal2 s 8574 0 8630 800 4 chany_bottom_in[5]
port 24 nsew
rlabel metal2 s 8942 0 8998 800 4 chany_bottom_in[6]
port 25 nsew
rlabel metal2 s 9218 0 9274 800 4 chany_bottom_in[7]
port 26 nsew
rlabel metal2 s 9586 0 9642 800 4 chany_bottom_in[8]
port 27 nsew
rlabel metal2 s 9954 0 10010 800 4 chany_bottom_in[9]
port 28 nsew
rlabel metal2 s 110 0 166 800 4 chany_bottom_out[0]
port 29 nsew
rlabel metal2 s 3514 0 3570 800 4 chany_bottom_out[10]
port 30 nsew
rlabel metal2 s 3790 0 3846 800 4 chany_bottom_out[11]
port 31 nsew
rlabel metal2 s 4158 0 4214 800 4 chany_bottom_out[12]
port 32 nsew
rlabel metal2 s 4526 0 4582 800 4 chany_bottom_out[13]
port 33 nsew
rlabel metal2 s 4802 0 4858 800 4 chany_bottom_out[14]
port 34 nsew
rlabel metal2 s 5170 0 5226 800 4 chany_bottom_out[15]
port 35 nsew
rlabel metal2 s 5538 0 5594 800 4 chany_bottom_out[16]
port 36 nsew
rlabel metal2 s 5814 0 5870 800 4 chany_bottom_out[17]
port 37 nsew
rlabel metal2 s 6182 0 6238 800 4 chany_bottom_out[18]
port 38 nsew
rlabel metal2 s 6550 0 6606 800 4 chany_bottom_out[19]
port 39 nsew
rlabel metal2 s 386 0 442 800 4 chany_bottom_out[1]
port 40 nsew
rlabel metal2 s 754 0 810 800 4 chany_bottom_out[2]
port 41 nsew
rlabel metal2 s 1122 0 1178 800 4 chany_bottom_out[3]
port 42 nsew
rlabel metal2 s 1398 0 1454 800 4 chany_bottom_out[4]
port 43 nsew
rlabel metal2 s 1766 0 1822 800 4 chany_bottom_out[5]
port 44 nsew
rlabel metal2 s 2134 0 2190 800 4 chany_bottom_out[6]
port 45 nsew
rlabel metal2 s 2410 0 2466 800 4 chany_bottom_out[7]
port 46 nsew
rlabel metal2 s 2778 0 2834 800 4 chany_bottom_out[8]
port 47 nsew
rlabel metal2 s 3146 0 3202 800 4 chany_bottom_out[9]
port 48 nsew
rlabel metal2 s 10322 19200 10378 20000 4 chany_top_in[0]
port 49 nsew
rlabel metal2 s 13726 19200 13782 20000 4 chany_top_in[10]
port 50 nsew
rlabel metal2 s 14002 19200 14058 20000 4 chany_top_in[11]
port 51 nsew
rlabel metal2 s 14370 19200 14426 20000 4 chany_top_in[12]
port 52 nsew
rlabel metal2 s 14738 19200 14794 20000 4 chany_top_in[13]
port 53 nsew
rlabel metal2 s 15014 19200 15070 20000 4 chany_top_in[14]
port 54 nsew
rlabel metal2 s 15382 19200 15438 20000 4 chany_top_in[15]
port 55 nsew
rlabel metal2 s 15750 19200 15806 20000 4 chany_top_in[16]
port 56 nsew
rlabel metal2 s 16026 19200 16082 20000 4 chany_top_in[17]
port 57 nsew
rlabel metal2 s 16394 19200 16450 20000 4 chany_top_in[18]
port 58 nsew
rlabel metal2 s 16762 19200 16818 20000 4 chany_top_in[19]
port 59 nsew
rlabel metal2 s 10598 19200 10654 20000 4 chany_top_in[1]
port 60 nsew
rlabel metal2 s 10966 19200 11022 20000 4 chany_top_in[2]
port 61 nsew
rlabel metal2 s 11334 19200 11390 20000 4 chany_top_in[3]
port 62 nsew
rlabel metal2 s 11610 19200 11666 20000 4 chany_top_in[4]
port 63 nsew
rlabel metal2 s 11978 19200 12034 20000 4 chany_top_in[5]
port 64 nsew
rlabel metal2 s 12346 19200 12402 20000 4 chany_top_in[6]
port 65 nsew
rlabel metal2 s 12622 19200 12678 20000 4 chany_top_in[7]
port 66 nsew
rlabel metal2 s 12990 19200 13046 20000 4 chany_top_in[8]
port 67 nsew
rlabel metal2 s 13358 19200 13414 20000 4 chany_top_in[9]
port 68 nsew
rlabel metal2 s 3514 19200 3570 20000 4 chany_top_out[0]
port 69 nsew
rlabel metal2 s 6918 19200 6974 20000 4 chany_top_out[10]
port 70 nsew
rlabel metal2 s 7194 19200 7250 20000 4 chany_top_out[11]
port 71 nsew
rlabel metal2 s 7562 19200 7618 20000 4 chany_top_out[12]
port 72 nsew
rlabel metal2 s 7930 19200 7986 20000 4 chany_top_out[13]
port 73 nsew
rlabel metal2 s 8206 19200 8262 20000 4 chany_top_out[14]
port 74 nsew
rlabel metal2 s 8574 19200 8630 20000 4 chany_top_out[15]
port 75 nsew
rlabel metal2 s 8942 19200 8998 20000 4 chany_top_out[16]
port 76 nsew
rlabel metal2 s 9218 19200 9274 20000 4 chany_top_out[17]
port 77 nsew
rlabel metal2 s 9586 19200 9642 20000 4 chany_top_out[18]
port 78 nsew
rlabel metal2 s 9954 19200 10010 20000 4 chany_top_out[19]
port 79 nsew
rlabel metal2 s 3790 19200 3846 20000 4 chany_top_out[1]
port 80 nsew
rlabel metal2 s 4158 19200 4214 20000 4 chany_top_out[2]
port 81 nsew
rlabel metal2 s 4526 19200 4582 20000 4 chany_top_out[3]
port 82 nsew
rlabel metal2 s 4802 19200 4858 20000 4 chany_top_out[4]
port 83 nsew
rlabel metal2 s 5170 19200 5226 20000 4 chany_top_out[5]
port 84 nsew
rlabel metal2 s 5538 19200 5594 20000 4 chany_top_out[6]
port 85 nsew
rlabel metal2 s 5814 19200 5870 20000 4 chany_top_out[7]
port 86 nsew
rlabel metal2 s 6182 19200 6238 20000 4 chany_top_out[8]
port 87 nsew
rlabel metal2 s 6550 19200 6606 20000 4 chany_top_out[9]
port 88 nsew
rlabel metal2 s 110 19200 166 20000 4 clk_2_N_in
port 89 nsew
rlabel metal2 s 1398 19200 1454 20000 4 clk_2_N_out
port 90 nsew
rlabel metal2 s 14002 0 14058 800 4 clk_2_S_in
port 91 nsew
rlabel metal2 s 15382 0 15438 800 4 clk_2_S_out
port 92 nsew
rlabel metal2 s 386 19200 442 20000 4 clk_3_N_in
port 93 nsew
rlabel metal2 s 1766 19200 1822 20000 4 clk_3_N_out
port 94 nsew
rlabel metal2 s 14370 0 14426 800 4 clk_3_S_in
port 95 nsew
rlabel metal2 s 15750 0 15806 800 4 clk_3_S_out
port 96 nsew
rlabel metal3 s 0 1368 800 1488 4 left_grid_pin_16_
port 97 nsew
rlabel metal3 s 0 2320 800 2440 4 left_grid_pin_17_
port 98 nsew
rlabel metal3 s 0 3408 800 3528 4 left_grid_pin_18_
port 99 nsew
rlabel metal3 s 0 4360 800 4480 4 left_grid_pin_19_
port 100 nsew
rlabel metal3 s 0 5312 800 5432 4 left_grid_pin_20_
port 101 nsew
rlabel metal3 s 0 6400 800 6520 4 left_grid_pin_21_
port 102 nsew
rlabel metal3 s 0 7352 800 7472 4 left_grid_pin_22_
port 103 nsew
rlabel metal3 s 0 8304 800 8424 4 left_grid_pin_23_
port 104 nsew
rlabel metal3 s 0 9392 800 9512 4 left_grid_pin_24_
port 105 nsew
rlabel metal3 s 0 10344 800 10464 4 left_grid_pin_25_
port 106 nsew
rlabel metal3 s 0 11296 800 11416 4 left_grid_pin_26_
port 107 nsew
rlabel metal3 s 0 12384 800 12504 4 left_grid_pin_27_
port 108 nsew
rlabel metal3 s 0 13336 800 13456 4 left_grid_pin_28_
port 109 nsew
rlabel metal3 s 0 14288 800 14408 4 left_grid_pin_29_
port 110 nsew
rlabel metal3 s 0 15376 800 15496 4 left_grid_pin_30_
port 111 nsew
rlabel metal3 s 0 16328 800 16448 4 left_grid_pin_31_
port 112 nsew
rlabel metal2 s 2134 19200 2190 20000 4 prog_clk_0_N_out
port 113 nsew
rlabel metal2 s 16026 0 16082 800 4 prog_clk_0_S_out
port 114 nsew
rlabel metal3 s 0 19320 800 19440 4 prog_clk_0_W_in
port 115 nsew
rlabel metal2 s 754 19200 810 20000 4 prog_clk_2_N_in
port 116 nsew
rlabel metal2 s 2410 19200 2466 20000 4 prog_clk_2_N_out
port 117 nsew
rlabel metal2 s 14738 0 14794 800 4 prog_clk_2_S_in
port 118 nsew
rlabel metal2 s 16394 0 16450 800 4 prog_clk_2_S_out
port 119 nsew
rlabel metal2 s 1122 19200 1178 20000 4 prog_clk_3_N_in
port 120 nsew
rlabel metal2 s 2778 19200 2834 20000 4 prog_clk_3_N_out
port 121 nsew
rlabel metal2 s 15014 0 15070 800 4 prog_clk_3_S_in
port 122 nsew
rlabel metal2 s 16762 0 16818 800 4 prog_clk_3_S_out
port 123 nsew
rlabel metal4 s 3409 2128 3729 17456 4 VPWR
port 124 nsew
rlabel metal4 s 5875 2128 6195 17456 4 VGND
port 125 nsew
<< properties >>
string FIXED_BBOX 0 0 17000 20000
string GDS_FILE /ef/openfpga/openlane/runs/cby_1__1_/results/magic/cby_1__1_.gds
string GDS_END 1148986
string GDS_START 81920
<< end >>
