magic
tech sky130A
magscale 1 2
timestamp 1606474019
<< locali >>
rect 10057 19227 10091 19397
rect 12265 18071 12299 18241
rect 12909 18207 12943 18309
rect 13829 18071 13863 18173
rect 12909 17527 12943 17833
rect 12541 16983 12575 17085
rect 13921 15895 13955 15997
rect 16497 15895 16531 16201
rect 10333 15555 10367 15657
rect 14105 15487 14139 15657
rect 16221 13719 16255 13957
rect 15025 5695 15059 5865
rect 11345 5015 11379 5321
<< viali >>
rect 8769 20009 8803 20043
rect 11897 20009 11931 20043
rect 13001 20009 13035 20043
rect 14565 20009 14599 20043
rect 16313 20009 16347 20043
rect 16865 20009 16899 20043
rect 17417 20009 17451 20043
rect 18521 20009 18555 20043
rect 19073 20009 19107 20043
rect 19625 20009 19659 20043
rect 20177 20009 20211 20043
rect 20729 20009 20763 20043
rect 10517 19941 10551 19975
rect 8585 19873 8619 19907
rect 9137 19873 9171 19907
rect 10425 19873 10459 19907
rect 11069 19873 11103 19907
rect 11989 19873 12023 19907
rect 12817 19873 12851 19907
rect 13829 19873 13863 19907
rect 14381 19873 14415 19907
rect 15577 19873 15611 19907
rect 16129 19873 16163 19907
rect 16681 19873 16715 19907
rect 17233 19873 17267 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 10609 19805 10643 19839
rect 12081 19805 12115 19839
rect 9321 19737 9355 19771
rect 14013 19737 14047 19771
rect 15761 19737 15795 19771
rect 10057 19669 10091 19703
rect 11529 19669 11563 19703
rect 9965 19397 9999 19431
rect 10057 19397 10091 19431
rect 8585 19261 8619 19295
rect 16405 19329 16439 19363
rect 10241 19261 10275 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 14749 19261 14783 19295
rect 15025 19261 15059 19295
rect 17049 19261 17083 19295
rect 18245 19261 18279 19295
rect 18521 19261 18555 19295
rect 19073 19261 19107 19295
rect 19625 19261 19659 19295
rect 8852 19193 8886 19227
rect 10057 19193 10091 19227
rect 10486 19193 10520 19227
rect 12694 19193 12728 19227
rect 17325 19193 17359 19227
rect 20453 19193 20487 19227
rect 11621 19125 11655 19159
rect 13829 19125 13863 19159
rect 14289 19125 14323 19159
rect 15761 19125 15795 19159
rect 16129 19125 16163 19159
rect 16221 19125 16255 19159
rect 19257 19125 19291 19159
rect 9229 18921 9263 18955
rect 10241 18921 10275 18955
rect 11989 18921 12023 18955
rect 14749 18921 14783 18955
rect 16681 18921 16715 18955
rect 17141 18921 17175 18955
rect 17785 18921 17819 18955
rect 18521 18921 18555 18955
rect 10876 18853 10910 18887
rect 12992 18853 13026 18887
rect 19993 18853 20027 18887
rect 7849 18785 7883 18819
rect 8116 18785 8150 18819
rect 10057 18785 10091 18819
rect 12725 18785 12759 18819
rect 14565 18785 14599 18819
rect 15557 18785 15591 18819
rect 16957 18785 16991 18819
rect 17601 18785 17635 18819
rect 19165 18785 19199 18819
rect 19717 18785 19751 18819
rect 10609 18717 10643 18751
rect 15301 18717 15335 18751
rect 18613 18717 18647 18751
rect 18797 18717 18831 18751
rect 14105 18581 14139 18615
rect 18153 18581 18187 18615
rect 19349 18581 19383 18615
rect 11989 18377 12023 18411
rect 12633 18377 12667 18411
rect 15393 18377 15427 18411
rect 15945 18377 15979 18411
rect 17693 18377 17727 18411
rect 19349 18377 19383 18411
rect 8861 18309 8895 18343
rect 12909 18309 12943 18343
rect 13001 18309 13035 18343
rect 18061 18309 18095 18343
rect 9413 18241 9447 18275
rect 10701 18241 10735 18275
rect 12265 18241 12299 18275
rect 9321 18173 9355 18207
rect 10425 18173 10459 18207
rect 11069 18173 11103 18207
rect 11805 18173 11839 18207
rect 9229 18105 9263 18139
rect 10517 18105 10551 18139
rect 11345 18105 11379 18139
rect 13461 18241 13495 18275
rect 13645 18241 13679 18275
rect 16313 18241 16347 18275
rect 18613 18241 18647 18275
rect 20729 18241 20763 18275
rect 12449 18173 12483 18207
rect 12909 18173 12943 18207
rect 13829 18173 13863 18207
rect 14013 18173 14047 18207
rect 14269 18173 14303 18207
rect 15761 18173 15795 18207
rect 18429 18173 18463 18207
rect 19165 18173 19199 18207
rect 19717 18173 19751 18207
rect 20453 18173 20487 18207
rect 16580 18105 16614 18139
rect 19993 18105 20027 18139
rect 10057 18037 10091 18071
rect 12265 18037 12299 18071
rect 13369 18037 13403 18071
rect 13829 18037 13863 18071
rect 18521 18037 18555 18071
rect 8861 17833 8895 17867
rect 9689 17833 9723 17867
rect 10149 17833 10183 17867
rect 12909 17833 12943 17867
rect 13001 17833 13035 17867
rect 13461 17833 13495 17867
rect 15761 17833 15795 17867
rect 18797 17833 18831 17867
rect 19257 17833 19291 17867
rect 20913 17833 20947 17867
rect 11989 17765 12023 17799
rect 7481 17697 7515 17731
rect 7748 17697 7782 17731
rect 10057 17697 10091 17731
rect 10793 17697 10827 17731
rect 11897 17697 11931 17731
rect 10241 17629 10275 17663
rect 11069 17629 11103 17663
rect 12081 17629 12115 17663
rect 12541 17629 12575 17663
rect 13369 17765 13403 17799
rect 14749 17765 14783 17799
rect 14013 17697 14047 17731
rect 15301 17697 15335 17731
rect 16129 17697 16163 17731
rect 17141 17697 17175 17731
rect 17408 17697 17442 17731
rect 19165 17697 19199 17731
rect 19809 17697 19843 17731
rect 13553 17629 13587 17663
rect 14289 17629 14323 17663
rect 16221 17629 16255 17663
rect 16405 17629 16439 17663
rect 19349 17629 19383 17663
rect 19993 17629 20027 17663
rect 18521 17561 18555 17595
rect 11529 17493 11563 17527
rect 12909 17493 12943 17527
rect 8401 17289 8435 17323
rect 12633 17289 12667 17323
rect 15761 17289 15795 17323
rect 11989 17221 12023 17255
rect 15393 17221 15427 17255
rect 17049 17221 17083 17255
rect 9229 17153 9263 17187
rect 10241 17153 10275 17187
rect 11161 17153 11195 17187
rect 11345 17153 11379 17187
rect 13093 17153 13127 17187
rect 13277 17153 13311 17187
rect 14565 17153 14599 17187
rect 16313 17153 16347 17187
rect 20545 17153 20579 17187
rect 7021 17085 7055 17119
rect 10149 17085 10183 17119
rect 11069 17085 11103 17119
rect 11805 17085 11839 17119
rect 12541 17085 12575 17119
rect 13001 17085 13035 17119
rect 15209 17085 15243 17119
rect 16865 17085 16899 17119
rect 17417 17085 17451 17119
rect 18061 17085 18095 17119
rect 18328 17085 18362 17119
rect 7288 17017 7322 17051
rect 10057 17017 10091 17051
rect 14381 17017 14415 17051
rect 20453 17017 20487 17051
rect 8677 16949 8711 16983
rect 9045 16949 9079 16983
rect 9137 16949 9171 16983
rect 9689 16949 9723 16983
rect 10701 16949 10735 16983
rect 12541 16949 12575 16983
rect 13921 16949 13955 16983
rect 14289 16949 14323 16983
rect 16129 16949 16163 16983
rect 16221 16949 16255 16983
rect 17601 16949 17635 16983
rect 19441 16949 19475 16983
rect 19993 16949 20027 16983
rect 20361 16949 20395 16983
rect 7389 16745 7423 16779
rect 7481 16745 7515 16779
rect 8217 16745 8251 16779
rect 9689 16745 9723 16779
rect 11621 16745 11655 16779
rect 15301 16745 15335 16779
rect 17141 16745 17175 16779
rect 19625 16745 19659 16779
rect 20085 16745 20119 16779
rect 8677 16677 8711 16711
rect 17233 16677 17267 16711
rect 18153 16677 18187 16711
rect 8585 16609 8619 16643
rect 9505 16609 9539 16643
rect 10241 16609 10275 16643
rect 10508 16609 10542 16643
rect 11897 16609 11931 16643
rect 12164 16609 12198 16643
rect 13553 16609 13587 16643
rect 13820 16609 13854 16643
rect 16129 16609 16163 16643
rect 17877 16609 17911 16643
rect 18981 16609 19015 16643
rect 19993 16609 20027 16643
rect 7665 16541 7699 16575
rect 8769 16541 8803 16575
rect 16221 16541 16255 16575
rect 16405 16541 16439 16575
rect 17325 16541 17359 16575
rect 19073 16541 19107 16575
rect 19257 16541 19291 16575
rect 20177 16541 20211 16575
rect 7021 16473 7055 16507
rect 9321 16473 9355 16507
rect 13277 16405 13311 16439
rect 14933 16405 14967 16439
rect 15761 16405 15795 16439
rect 16773 16405 16807 16439
rect 18613 16405 18647 16439
rect 8217 16201 8251 16235
rect 12449 16201 12483 16235
rect 16497 16201 16531 16235
rect 9413 16065 9447 16099
rect 11529 16065 11563 16099
rect 11713 16065 11747 16099
rect 13093 16065 13127 16099
rect 14013 16065 14047 16099
rect 16129 16065 16163 16099
rect 16221 16065 16255 16099
rect 6837 15997 6871 16031
rect 8677 15997 8711 16031
rect 12817 15997 12851 16031
rect 12909 15997 12943 16031
rect 13461 15997 13495 16031
rect 13921 15997 13955 16031
rect 7104 15929 7138 15963
rect 8953 15929 8987 15963
rect 9680 15929 9714 15963
rect 11437 15929 11471 15963
rect 14280 15929 14314 15963
rect 16037 15929 16071 15963
rect 17141 16065 17175 16099
rect 17325 16065 17359 16099
rect 20361 16065 20395 16099
rect 17049 15997 17083 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 20821 15997 20855 16031
rect 18328 15929 18362 15963
rect 20177 15929 20211 15963
rect 20269 15929 20303 15963
rect 10793 15861 10827 15895
rect 11069 15861 11103 15895
rect 13645 15861 13679 15895
rect 13921 15861 13955 15895
rect 15393 15861 15427 15895
rect 15669 15861 15703 15895
rect 16497 15861 16531 15895
rect 16681 15861 16715 15895
rect 17693 15861 17727 15895
rect 19441 15861 19475 15895
rect 19809 15861 19843 15895
rect 21005 15861 21039 15895
rect 10333 15657 10367 15691
rect 10425 15657 10459 15691
rect 10793 15657 10827 15691
rect 13185 15657 13219 15691
rect 14105 15657 14139 15691
rect 15301 15657 15335 15691
rect 15669 15657 15703 15691
rect 17785 15657 17819 15691
rect 18061 15657 18095 15691
rect 19901 15657 19935 15691
rect 20453 15657 20487 15691
rect 6460 15589 6494 15623
rect 6193 15521 6227 15555
rect 8861 15521 8895 15555
rect 9689 15521 9723 15555
rect 10333 15521 10367 15555
rect 11529 15521 11563 15555
rect 11796 15521 11830 15555
rect 13553 15521 13587 15555
rect 14565 15589 14599 15623
rect 18788 15589 18822 15623
rect 16672 15521 16706 15555
rect 18521 15521 18555 15555
rect 20269 15521 20303 15555
rect 9137 15453 9171 15487
rect 9965 15453 9999 15487
rect 10885 15453 10919 15487
rect 10977 15453 11011 15487
rect 13645 15453 13679 15487
rect 13737 15453 13771 15487
rect 14105 15453 14139 15487
rect 14657 15453 14691 15487
rect 14841 15453 14875 15487
rect 15761 15453 15795 15487
rect 15853 15453 15887 15487
rect 16405 15453 16439 15487
rect 14197 15385 14231 15419
rect 7573 15317 7607 15351
rect 12909 15317 12943 15351
rect 5733 15113 5767 15147
rect 10333 15113 10367 15147
rect 18521 15113 18555 15147
rect 19625 15113 19659 15147
rect 20821 15113 20855 15147
rect 9045 15045 9079 15079
rect 12817 15045 12851 15079
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 9781 14977 9815 15011
rect 9873 14977 9907 15011
rect 10793 14977 10827 15011
rect 10977 14977 11011 15011
rect 11897 14977 11931 15011
rect 13645 14977 13679 15011
rect 14289 14977 14323 15011
rect 17233 14977 17267 15011
rect 19073 14977 19107 15011
rect 20085 14977 20119 15011
rect 20269 14977 20303 15011
rect 6101 14909 6135 14943
rect 7665 14909 7699 14943
rect 7932 14909 7966 14943
rect 13001 14909 13035 14943
rect 14556 14909 14590 14943
rect 16129 14909 16163 14943
rect 18889 14909 18923 14943
rect 20637 14909 20671 14943
rect 10701 14841 10735 14875
rect 17049 14841 17083 14875
rect 18981 14841 19015 14875
rect 9321 14773 9355 14807
rect 9689 14773 9723 14807
rect 11345 14773 11379 14807
rect 11713 14773 11747 14807
rect 11805 14773 11839 14807
rect 13093 14773 13127 14807
rect 13461 14773 13495 14807
rect 13553 14773 13587 14807
rect 15669 14773 15703 14807
rect 16313 14773 16347 14807
rect 16681 14773 16715 14807
rect 17141 14773 17175 14807
rect 19993 14773 20027 14807
rect 8493 14569 8527 14603
rect 8953 14569 8987 14603
rect 11345 14569 11379 14603
rect 13001 14569 13035 14603
rect 13645 14569 13679 14603
rect 13737 14569 13771 14603
rect 17509 14569 17543 14603
rect 20453 14569 20487 14603
rect 7104 14501 7138 14535
rect 9956 14501 9990 14535
rect 14565 14501 14599 14535
rect 16396 14501 16430 14535
rect 6837 14433 6871 14467
rect 8861 14433 8895 14467
rect 11529 14433 11563 14467
rect 11888 14433 11922 14467
rect 14289 14433 14323 14467
rect 15301 14433 15335 14467
rect 16129 14433 16163 14467
rect 18153 14433 18187 14467
rect 19073 14433 19107 14467
rect 19340 14433 19374 14467
rect 9045 14365 9079 14399
rect 9689 14365 9723 14399
rect 11621 14365 11655 14399
rect 13829 14365 13863 14399
rect 15577 14365 15611 14399
rect 18245 14365 18279 14399
rect 18337 14365 18371 14399
rect 20913 14365 20947 14399
rect 8217 14229 8251 14263
rect 11069 14229 11103 14263
rect 13277 14229 13311 14263
rect 17785 14229 17819 14263
rect 8493 14025 8527 14059
rect 12449 14025 12483 14059
rect 13645 14025 13679 14059
rect 14657 14025 14691 14059
rect 17693 14025 17727 14059
rect 18061 14025 18095 14059
rect 19809 14025 19843 14059
rect 21005 14025 21039 14059
rect 11345 13957 11379 13991
rect 16221 13957 16255 13991
rect 9137 13889 9171 13923
rect 10793 13889 10827 13923
rect 11897 13889 11931 13923
rect 13093 13889 13127 13923
rect 14105 13889 14139 13923
rect 14289 13889 14323 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 8953 13821 8987 13855
rect 10609 13821 10643 13855
rect 11805 13821 11839 13855
rect 12817 13821 12851 13855
rect 15761 13821 15795 13855
rect 8861 13753 8895 13787
rect 9505 13753 9539 13787
rect 15025 13753 15059 13787
rect 18613 13889 18647 13923
rect 20361 13889 20395 13923
rect 16313 13821 16347 13855
rect 18521 13821 18555 13855
rect 19073 13821 19107 13855
rect 20177 13821 20211 13855
rect 20821 13821 20855 13855
rect 16580 13753 16614 13787
rect 19349 13753 19383 13787
rect 20269 13753 20303 13787
rect 10149 13685 10183 13719
rect 10517 13685 10551 13719
rect 11713 13685 11747 13719
rect 12909 13685 12943 13719
rect 14013 13685 14047 13719
rect 15945 13685 15979 13719
rect 16221 13685 16255 13719
rect 18429 13685 18463 13719
rect 9321 13481 9355 13515
rect 11345 13481 11379 13515
rect 11713 13481 11747 13515
rect 12725 13481 12759 13515
rect 14013 13481 14047 13515
rect 16313 13481 16347 13515
rect 17141 13481 17175 13515
rect 17233 13481 17267 13515
rect 18245 13481 18279 13515
rect 18981 13481 19015 13515
rect 19809 13481 19843 13515
rect 11805 13413 11839 13447
rect 9505 13345 9539 13379
rect 9689 13345 9723 13379
rect 9956 13345 9990 13379
rect 12909 13345 12943 13379
rect 13093 13345 13127 13379
rect 14657 13345 14691 13379
rect 15669 13345 15703 13379
rect 18153 13345 18187 13379
rect 18797 13345 18831 13379
rect 19717 13345 19751 13379
rect 11897 13277 11931 13311
rect 13369 13277 13403 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 17417 13277 17451 13311
rect 18429 13277 18463 13311
rect 19993 13277 20027 13311
rect 14841 13209 14875 13243
rect 15301 13209 15335 13243
rect 17785 13209 17819 13243
rect 11069 13141 11103 13175
rect 16773 13141 16807 13175
rect 19349 13141 19383 13175
rect 10609 12937 10643 12971
rect 16589 12937 16623 12971
rect 16865 12937 16899 12971
rect 20177 12937 20211 12971
rect 12449 12869 12483 12903
rect 11069 12801 11103 12835
rect 11161 12801 11195 12835
rect 13093 12801 13127 12835
rect 17509 12801 17543 12835
rect 18337 12801 18371 12835
rect 20729 12801 20763 12835
rect 8953 12733 8987 12767
rect 11621 12733 11655 12767
rect 13553 12733 13587 12767
rect 15209 12733 15243 12767
rect 18061 12733 18095 12767
rect 18797 12733 18831 12767
rect 20453 12733 20487 12767
rect 9220 12665 9254 12699
rect 11897 12665 11931 12699
rect 13820 12665 13854 12699
rect 15476 12665 15510 12699
rect 17233 12665 17267 12699
rect 19064 12665 19098 12699
rect 10333 12597 10367 12631
rect 10977 12597 11011 12631
rect 12817 12597 12851 12631
rect 12909 12597 12943 12631
rect 14933 12597 14967 12631
rect 17325 12597 17359 12631
rect 12817 12393 12851 12427
rect 17601 12393 17635 12427
rect 19993 12393 20027 12427
rect 8024 12325 8058 12359
rect 13338 12325 13372 12359
rect 16190 12325 16224 12359
rect 17969 12325 18003 12359
rect 20913 12325 20947 12359
rect 7757 12257 7791 12291
rect 10701 12257 10735 12291
rect 10793 12257 10827 12291
rect 11704 12257 11738 12291
rect 13093 12257 13127 12291
rect 18880 12257 18914 12291
rect 20269 12257 20303 12291
rect 10885 12189 10919 12223
rect 11437 12189 11471 12223
rect 15301 12189 15335 12223
rect 15945 12189 15979 12223
rect 18061 12189 18095 12223
rect 18245 12189 18279 12223
rect 18613 12189 18647 12223
rect 10333 12121 10367 12155
rect 9137 12053 9171 12087
rect 14473 12053 14507 12087
rect 17325 12053 17359 12087
rect 20453 12053 20487 12087
rect 11529 11849 11563 11883
rect 12541 11849 12575 11883
rect 15485 11849 15519 11883
rect 16497 11849 16531 11883
rect 19349 11849 19383 11883
rect 21097 11849 21131 11883
rect 13461 11781 13495 11815
rect 10609 11713 10643 11747
rect 12081 11713 12115 11747
rect 13093 11713 13127 11747
rect 14105 11713 14139 11747
rect 14933 11713 14967 11747
rect 16037 11713 16071 11747
rect 17509 11713 17543 11747
rect 18613 11713 18647 11747
rect 19717 11713 19751 11747
rect 9413 11645 9447 11679
rect 11253 11645 11287 11679
rect 11897 11645 11931 11679
rect 15945 11645 15979 11679
rect 16681 11645 16715 11679
rect 19165 11645 19199 11679
rect 9689 11577 9723 11611
rect 15853 11577 15887 11611
rect 17233 11577 17267 11611
rect 17325 11577 17359 11611
rect 18429 11577 18463 11611
rect 19984 11577 20018 11611
rect 8953 11509 8987 11543
rect 11989 11509 12023 11543
rect 12909 11509 12943 11543
rect 13001 11509 13035 11543
rect 13829 11509 13863 11543
rect 13921 11509 13955 11543
rect 14289 11509 14323 11543
rect 14657 11509 14691 11543
rect 14749 11509 14783 11543
rect 16865 11509 16899 11543
rect 18061 11509 18095 11543
rect 18521 11509 18555 11543
rect 9689 11305 9723 11339
rect 10057 11305 10091 11339
rect 12265 11305 12299 11339
rect 14289 11305 14323 11339
rect 15669 11305 15703 11339
rect 20085 11305 20119 11339
rect 8208 11237 8242 11271
rect 16405 11237 16439 11271
rect 16948 11237 16982 11271
rect 18797 11237 18831 11271
rect 7941 11169 7975 11203
rect 10885 11169 10919 11203
rect 11152 11169 11186 11203
rect 13001 11169 13035 11203
rect 16129 11169 16163 11203
rect 18705 11169 18739 11203
rect 19993 11169 20027 11203
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 16681 11101 16715 11135
rect 18889 11101 18923 11135
rect 20177 11101 20211 11135
rect 9321 11033 9355 11067
rect 18337 11033 18371 11067
rect 15301 10965 15335 10999
rect 18061 10965 18095 10999
rect 19625 10965 19659 10999
rect 8769 10761 8803 10795
rect 12449 10761 12483 10795
rect 13461 10761 13495 10795
rect 15393 10761 15427 10795
rect 11345 10693 11379 10727
rect 9321 10625 9355 10659
rect 10057 10625 10091 10659
rect 11897 10625 11931 10659
rect 13093 10625 13127 10659
rect 14013 10625 14047 10659
rect 15117 10625 15151 10659
rect 15853 10625 15887 10659
rect 16037 10625 16071 10659
rect 18061 10625 18095 10659
rect 19257 10625 19291 10659
rect 9781 10557 9815 10591
rect 12817 10557 12851 10591
rect 13829 10557 13863 10591
rect 15025 10557 15059 10591
rect 15761 10557 15795 10591
rect 16313 10557 16347 10591
rect 19073 10557 19107 10591
rect 19625 10557 19659 10591
rect 11805 10489 11839 10523
rect 14933 10489 14967 10523
rect 16580 10489 16614 10523
rect 19870 10489 19904 10523
rect 9137 10421 9171 10455
rect 9229 10421 9263 10455
rect 11713 10421 11747 10455
rect 12909 10421 12943 10455
rect 13921 10421 13955 10455
rect 14565 10421 14599 10455
rect 17693 10421 17727 10455
rect 18613 10421 18647 10455
rect 18981 10421 19015 10455
rect 21005 10421 21039 10455
rect 11989 10217 12023 10251
rect 13645 10217 13679 10251
rect 14197 10217 14231 10251
rect 16681 10217 16715 10251
rect 16957 10217 16991 10251
rect 17325 10217 17359 10251
rect 18153 10217 18187 10251
rect 18613 10217 18647 10251
rect 20545 10217 20579 10251
rect 8208 10149 8242 10183
rect 13553 10149 13587 10183
rect 14657 10149 14691 10183
rect 18521 10149 18555 10183
rect 10517 10081 10551 10115
rect 10876 10081 10910 10115
rect 14565 10081 14599 10115
rect 15568 10081 15602 10115
rect 19165 10081 19199 10115
rect 19432 10081 19466 10115
rect 7941 10013 7975 10047
rect 9689 10013 9723 10047
rect 10609 10013 10643 10047
rect 13737 10013 13771 10047
rect 14749 10013 14783 10047
rect 15301 10013 15335 10047
rect 17417 10013 17451 10047
rect 17601 10013 17635 10047
rect 18797 10013 18831 10047
rect 10333 9945 10367 9979
rect 9321 9877 9355 9911
rect 13185 9877 13219 9911
rect 14565 9673 14599 9707
rect 15577 9673 15611 9707
rect 16957 9673 16991 9707
rect 11345 9605 11379 9639
rect 11897 9537 11931 9571
rect 15209 9537 15243 9571
rect 16221 9537 16255 9571
rect 17509 9537 17543 9571
rect 20637 9537 20671 9571
rect 8217 9469 8251 9503
rect 8484 9469 8518 9503
rect 9965 9469 9999 9503
rect 11621 9469 11655 9503
rect 12449 9469 12483 9503
rect 14289 9469 14323 9503
rect 14933 9469 14967 9503
rect 17325 9469 17359 9503
rect 17417 9469 17451 9503
rect 18061 9469 18095 9503
rect 20545 9469 20579 9503
rect 10232 9401 10266 9435
rect 12716 9401 12750 9435
rect 18306 9401 18340 9435
rect 9597 9333 9631 9367
rect 13829 9333 13863 9367
rect 14105 9333 14139 9367
rect 15025 9333 15059 9367
rect 15945 9333 15979 9367
rect 16037 9333 16071 9367
rect 19441 9333 19475 9367
rect 20085 9333 20119 9367
rect 20453 9333 20487 9367
rect 8585 9129 8619 9163
rect 8953 9129 8987 9163
rect 11437 9129 11471 9163
rect 12449 9129 12483 9163
rect 15301 9129 15335 9163
rect 17141 9129 17175 9163
rect 17693 9129 17727 9163
rect 18061 9129 18095 9163
rect 20361 9129 20395 9163
rect 13268 9061 13302 9095
rect 18972 9061 19006 9095
rect 10048 8993 10082 9027
rect 11805 8993 11839 9027
rect 12633 8993 12667 9027
rect 13001 8993 13035 9027
rect 15761 8993 15795 9027
rect 16028 8993 16062 9027
rect 17601 8993 17635 9027
rect 18705 8993 18739 9027
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 9781 8925 9815 8959
rect 11897 8925 11931 8959
rect 11989 8925 12023 8959
rect 18153 8925 18187 8959
rect 18337 8925 18371 8959
rect 11161 8857 11195 8891
rect 17417 8857 17451 8891
rect 20085 8857 20119 8891
rect 14381 8789 14415 8823
rect 8217 8585 8251 8619
rect 10609 8585 10643 8619
rect 10885 8585 10919 8619
rect 15209 8585 15243 8619
rect 12449 8517 12483 8551
rect 18613 8517 18647 8551
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 11437 8449 11471 8483
rect 13001 8449 13035 8483
rect 14381 8449 14415 8483
rect 16405 8449 16439 8483
rect 17233 8449 17267 8483
rect 17417 8449 17451 8483
rect 19165 8449 19199 8483
rect 20269 8449 20303 8483
rect 9229 8381 9263 8415
rect 11345 8381 11379 8415
rect 15393 8381 15427 8415
rect 18981 8381 19015 8415
rect 8585 8313 8619 8347
rect 9496 8313 9530 8347
rect 11253 8313 11287 8347
rect 11897 8313 11931 8347
rect 12817 8313 12851 8347
rect 14197 8313 14231 8347
rect 17141 8313 17175 8347
rect 12909 8245 12943 8279
rect 13829 8245 13863 8279
rect 14289 8245 14323 8279
rect 15761 8245 15795 8279
rect 16129 8245 16163 8279
rect 16221 8245 16255 8279
rect 16773 8245 16807 8279
rect 19073 8245 19107 8279
rect 19625 8245 19659 8279
rect 19993 8245 20027 8279
rect 20085 8245 20119 8279
rect 9873 8041 9907 8075
rect 12541 8041 12575 8075
rect 15669 8041 15703 8075
rect 20269 8041 20303 8075
rect 20913 8041 20947 8075
rect 9137 7973 9171 8007
rect 19156 7973 19190 8007
rect 8861 7905 8895 7939
rect 10241 7905 10275 7939
rect 11152 7905 11186 7939
rect 12909 7905 12943 7939
rect 13820 7905 13854 7939
rect 16037 7905 16071 7939
rect 16129 7905 16163 7939
rect 16948 7905 16982 7939
rect 18889 7905 18923 7939
rect 10333 7837 10367 7871
rect 10517 7837 10551 7871
rect 10885 7837 10919 7871
rect 13001 7837 13035 7871
rect 13185 7837 13219 7871
rect 13553 7837 13587 7871
rect 16313 7837 16347 7871
rect 16681 7837 16715 7871
rect 12265 7701 12299 7735
rect 14933 7701 14967 7735
rect 18061 7701 18095 7735
rect 9781 7497 9815 7531
rect 10333 7497 10367 7531
rect 11345 7497 11379 7531
rect 12817 7497 12851 7531
rect 13829 7497 13863 7531
rect 16865 7497 16899 7531
rect 10885 7361 10919 7395
rect 11897 7361 11931 7395
rect 13369 7361 13403 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 15485 7361 15519 7395
rect 18613 7361 18647 7395
rect 20453 7361 20487 7395
rect 8401 7293 8435 7327
rect 11713 7293 11747 7327
rect 13277 7293 13311 7327
rect 14197 7293 14231 7327
rect 15752 7293 15786 7327
rect 17141 7293 17175 7327
rect 18429 7293 18463 7327
rect 20361 7293 20395 7327
rect 8668 7225 8702 7259
rect 10793 7225 10827 7259
rect 13185 7225 13219 7259
rect 14841 7225 14875 7259
rect 10701 7157 10735 7191
rect 11805 7157 11839 7191
rect 18061 7157 18095 7191
rect 18521 7157 18555 7191
rect 19901 7157 19935 7191
rect 20269 7157 20303 7191
rect 9689 6953 9723 6987
rect 11069 6953 11103 6987
rect 13829 6953 13863 6987
rect 14289 6953 14323 6987
rect 16865 6953 16899 6987
rect 17233 6953 17267 6987
rect 18245 6953 18279 6987
rect 20545 6953 20579 6987
rect 15669 6885 15703 6919
rect 10057 6817 10091 6851
rect 11161 6817 11195 6851
rect 11969 6817 12003 6851
rect 14197 6817 14231 6851
rect 15761 6817 15795 6851
rect 16497 6817 16531 6851
rect 18337 6817 18371 6851
rect 19432 6817 19466 6851
rect 9137 6749 9171 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11253 6749 11287 6783
rect 11713 6749 11747 6783
rect 14381 6749 14415 6783
rect 15853 6749 15887 6783
rect 17325 6749 17359 6783
rect 17509 6749 17543 6783
rect 18521 6749 18555 6783
rect 19165 6749 19199 6783
rect 17877 6681 17911 6715
rect 10701 6613 10735 6647
rect 13093 6613 13127 6647
rect 15301 6613 15335 6647
rect 16313 6613 16347 6647
rect 9873 6409 9907 6443
rect 10149 6409 10183 6443
rect 18245 6409 18279 6443
rect 20637 6409 20671 6443
rect 10701 6273 10735 6307
rect 11713 6273 11747 6307
rect 13093 6273 13127 6307
rect 14105 6273 14139 6307
rect 15025 6273 15059 6307
rect 16313 6273 16347 6307
rect 17233 6273 17267 6307
rect 18889 6273 18923 6307
rect 6837 6205 6871 6239
rect 8493 6205 8527 6239
rect 10517 6205 10551 6239
rect 11621 6205 11655 6239
rect 13921 6205 13955 6239
rect 16129 6205 16163 6239
rect 19257 6205 19291 6239
rect 19524 6205 19558 6239
rect 7082 6137 7116 6171
rect 8738 6137 8772 6171
rect 11529 6137 11563 6171
rect 12817 6137 12851 6171
rect 14841 6137 14875 6171
rect 16037 6137 16071 6171
rect 17141 6137 17175 6171
rect 18613 6137 18647 6171
rect 8217 6069 8251 6103
rect 10609 6069 10643 6103
rect 11161 6069 11195 6103
rect 12449 6069 12483 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 13829 6069 13863 6103
rect 14473 6069 14507 6103
rect 14933 6069 14967 6103
rect 15669 6069 15703 6103
rect 16681 6069 16715 6103
rect 17049 6069 17083 6103
rect 18705 6069 18739 6103
rect 9781 5865 9815 5899
rect 10149 5865 10183 5899
rect 13093 5865 13127 5899
rect 14197 5865 14231 5899
rect 14565 5865 14599 5899
rect 15025 5865 15059 5899
rect 16681 5865 16715 5899
rect 18613 5865 18647 5899
rect 20913 5865 20947 5899
rect 11244 5797 11278 5831
rect 10977 5729 11011 5763
rect 13001 5729 13035 5763
rect 14657 5729 14691 5763
rect 15568 5797 15602 5831
rect 19134 5797 19168 5831
rect 15301 5729 15335 5763
rect 17500 5729 17534 5763
rect 10241 5661 10275 5695
rect 10333 5661 10367 5695
rect 13277 5661 13311 5695
rect 13645 5661 13679 5695
rect 14841 5661 14875 5695
rect 15025 5661 15059 5695
rect 17233 5661 17267 5695
rect 18889 5661 18923 5695
rect 12357 5593 12391 5627
rect 12633 5525 12667 5559
rect 20269 5525 20303 5559
rect 10425 5321 10459 5355
rect 11345 5321 11379 5355
rect 11437 5321 11471 5355
rect 12541 5321 12575 5355
rect 15117 5321 15151 5355
rect 17325 5321 17359 5355
rect 19901 5321 19935 5355
rect 10977 5185 11011 5219
rect 10885 5117 10919 5151
rect 10793 5049 10827 5083
rect 20177 5253 20211 5287
rect 13093 5185 13127 5219
rect 15945 5185 15979 5219
rect 18521 5185 18555 5219
rect 20729 5185 20763 5219
rect 11621 5117 11655 5151
rect 12909 5117 12943 5151
rect 13737 5117 13771 5151
rect 15393 5117 15427 5151
rect 16212 5117 16246 5151
rect 18788 5117 18822 5151
rect 13982 5049 14016 5083
rect 20545 5049 20579 5083
rect 11345 4981 11379 5015
rect 13001 4981 13035 5015
rect 15577 4981 15611 5015
rect 20637 4981 20671 5015
rect 13645 4777 13679 4811
rect 15301 4777 15335 4811
rect 15669 4777 15703 4811
rect 16313 4777 16347 4811
rect 17785 4777 17819 4811
rect 19165 4777 19199 4811
rect 20177 4777 20211 4811
rect 12532 4709 12566 4743
rect 12265 4641 12299 4675
rect 13921 4641 13955 4675
rect 14565 4641 14599 4675
rect 15761 4641 15795 4675
rect 17325 4641 17359 4675
rect 18153 4641 18187 4675
rect 19257 4641 19291 4675
rect 15945 4573 15979 4607
rect 18245 4573 18279 4607
rect 18337 4573 18371 4607
rect 19441 4573 19475 4607
rect 20269 4573 20303 4607
rect 20361 4573 20395 4607
rect 14105 4437 14139 4471
rect 14749 4437 14783 4471
rect 18797 4437 18831 4471
rect 19809 4437 19843 4471
rect 12817 4233 12851 4267
rect 19717 4233 19751 4267
rect 14013 4165 14047 4199
rect 11437 4097 11471 4131
rect 13369 4097 13403 4131
rect 14565 4097 14599 4131
rect 20269 4097 20303 4131
rect 9137 4029 9171 4063
rect 9393 4029 9427 4063
rect 13185 4029 13219 4063
rect 15025 4029 15059 4063
rect 15761 4029 15795 4063
rect 16037 4029 16071 4063
rect 16497 4029 16531 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 20085 4029 20119 4063
rect 20177 4029 20211 4063
rect 20729 4029 20763 4063
rect 11161 3961 11195 3995
rect 11805 3961 11839 3995
rect 13277 3961 13311 3995
rect 14473 3961 14507 3995
rect 18328 3961 18362 3995
rect 10517 3893 10551 3927
rect 10793 3893 10827 3927
rect 11253 3893 11287 3927
rect 14381 3893 14415 3927
rect 15209 3893 15243 3927
rect 16681 3893 16715 3927
rect 17601 3893 17635 3927
rect 19441 3893 19475 3927
rect 20913 3893 20947 3927
rect 11437 3689 11471 3723
rect 14749 3689 14783 3723
rect 16957 3689 16991 3723
rect 18613 3689 18647 3723
rect 11958 3621 11992 3655
rect 17478 3621 17512 3655
rect 10324 3553 10358 3587
rect 13369 3553 13403 3587
rect 13625 3553 13659 3587
rect 15577 3553 15611 3587
rect 15844 3553 15878 3587
rect 17233 3553 17267 3587
rect 19073 3553 19107 3587
rect 19809 3553 19843 3587
rect 10057 3485 10091 3519
rect 11713 3485 11747 3519
rect 19349 3485 19383 3519
rect 20085 3485 20119 3519
rect 13093 3417 13127 3451
rect 10425 3145 10459 3179
rect 13369 3145 13403 3179
rect 16497 3145 16531 3179
rect 18061 3145 18095 3179
rect 15761 3077 15795 3111
rect 19625 3077 19659 3111
rect 10977 3009 11011 3043
rect 13921 3009 13955 3043
rect 14381 3009 14415 3043
rect 16037 3009 16071 3043
rect 17141 3009 17175 3043
rect 18613 3009 18647 3043
rect 10885 2941 10919 2975
rect 11621 2941 11655 2975
rect 12449 2941 12483 2975
rect 13737 2941 13771 2975
rect 18429 2941 18463 2975
rect 18889 2941 18923 2975
rect 19441 2941 19475 2975
rect 19993 2941 20027 2975
rect 20545 2941 20579 2975
rect 11897 2873 11931 2907
rect 12725 2873 12759 2907
rect 14626 2873 14660 2907
rect 16865 2873 16899 2907
rect 17509 2873 17543 2907
rect 18521 2873 18555 2907
rect 10793 2805 10827 2839
rect 13829 2805 13863 2839
rect 16957 2805 16991 2839
rect 20177 2805 20211 2839
rect 20729 2805 20763 2839
rect 14473 2601 14507 2635
rect 15577 2601 15611 2635
rect 13829 2533 13863 2567
rect 15945 2533 15979 2567
rect 11345 2465 11379 2499
rect 11897 2465 11931 2499
rect 12817 2465 12851 2499
rect 13553 2465 13587 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 16589 2465 16623 2499
rect 17325 2465 17359 2499
rect 18429 2465 18463 2499
rect 18981 2465 19015 2499
rect 19533 2465 19567 2499
rect 20361 2465 20395 2499
rect 13093 2397 13127 2431
rect 16037 2397 16071 2431
rect 16129 2397 16163 2431
rect 11529 2329 11563 2363
rect 15025 2329 15059 2363
rect 19717 2329 19751 2363
rect 12081 2261 12115 2295
rect 16773 2261 16807 2295
rect 17509 2261 17543 2295
rect 18613 2261 18647 2295
rect 19165 2261 19199 2295
rect 20545 2261 20579 2295
<< metal1 >>
rect 7466 20272 7472 20324
rect 7524 20312 7530 20324
rect 11882 20312 11888 20324
rect 7524 20284 11888 20312
rect 7524 20272 7530 20284
rect 11882 20272 11888 20284
rect 11940 20272 11946 20324
rect 8754 20204 8760 20256
rect 8812 20244 8818 20256
rect 22462 20244 22468 20256
rect 8812 20216 22468 20244
rect 8812 20204 8818 20216
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 8754 20040 8760 20052
rect 8715 20012 8760 20040
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 10594 20040 10600 20052
rect 10336 20012 10600 20040
rect 10336 19972 10364 20012
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11388 20012 11897 20040
rect 11388 20000 11394 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 12989 20043 13047 20049
rect 12989 20009 13001 20043
rect 13035 20040 13047 20043
rect 13078 20040 13084 20052
rect 13035 20012 13084 20040
rect 13035 20009 13047 20012
rect 12989 20003 13047 20009
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 14182 20000 14188 20052
rect 14240 20040 14246 20052
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 14240 20012 14565 20040
rect 14240 20000 14246 20012
rect 14553 20009 14565 20012
rect 14599 20009 14611 20043
rect 14553 20003 14611 20009
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 15896 20012 16313 20040
rect 15896 20000 15902 20012
rect 16301 20009 16313 20012
rect 16347 20009 16359 20043
rect 16301 20003 16359 20009
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16632 20012 16865 20040
rect 16632 20000 16638 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 17405 20043 17463 20049
rect 17405 20009 17417 20043
rect 17451 20040 17463 20043
rect 17494 20040 17500 20052
rect 17451 20012 17500 20040
rect 17451 20009 17463 20012
rect 17405 20003 17463 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18506 20040 18512 20052
rect 18467 20012 18512 20040
rect 18506 20000 18512 20012
rect 18564 20000 18570 20052
rect 18598 20000 18604 20052
rect 18656 20040 18662 20052
rect 19061 20043 19119 20049
rect 19061 20040 19073 20043
rect 18656 20012 19073 20040
rect 18656 20000 18662 20012
rect 19061 20009 19073 20012
rect 19107 20009 19119 20043
rect 19061 20003 19119 20009
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 19613 20043 19671 20049
rect 19613 20040 19625 20043
rect 19392 20012 19625 20040
rect 19392 20000 19398 20012
rect 19613 20009 19625 20012
rect 19659 20009 19671 20043
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 19613 20003 19671 20009
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 8588 19944 10364 19972
rect 10505 19975 10563 19981
rect 8588 19913 8616 19944
rect 10505 19941 10517 19975
rect 10551 19972 10563 19975
rect 17310 19972 17316 19984
rect 10551 19944 17316 19972
rect 10551 19941 10563 19944
rect 10505 19935 10563 19941
rect 17310 19932 17316 19944
rect 17368 19932 17374 19984
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 10226 19904 10232 19916
rect 9171 19876 10232 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 10226 19864 10232 19876
rect 10284 19864 10290 19916
rect 10413 19907 10471 19913
rect 10413 19873 10425 19907
rect 10459 19904 10471 19907
rect 11057 19907 11115 19913
rect 11057 19904 11069 19907
rect 10459 19876 11069 19904
rect 10459 19873 10471 19876
rect 10413 19867 10471 19873
rect 11057 19873 11069 19876
rect 11103 19873 11115 19907
rect 11057 19867 11115 19873
rect 11882 19864 11888 19916
rect 11940 19904 11946 19916
rect 11977 19907 12035 19913
rect 11977 19904 11989 19907
rect 11940 19876 11989 19904
rect 11940 19864 11946 19876
rect 11977 19873 11989 19876
rect 12023 19873 12035 19907
rect 12802 19904 12808 19916
rect 12763 19876 12808 19904
rect 11977 19867 12035 19873
rect 12802 19864 12808 19876
rect 12860 19864 12866 19916
rect 13814 19904 13820 19916
rect 13775 19876 13820 19904
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 14366 19904 14372 19916
rect 14327 19876 14372 19904
rect 14366 19864 14372 19876
rect 14424 19864 14430 19916
rect 15562 19904 15568 19916
rect 15523 19876 15568 19904
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 16117 19907 16175 19913
rect 16117 19904 16129 19907
rect 15804 19876 16129 19904
rect 15804 19864 15810 19876
rect 16117 19873 16129 19876
rect 16163 19873 16175 19907
rect 16117 19867 16175 19873
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 16448 19876 16681 19904
rect 16448 19864 16454 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 17221 19907 17279 19913
rect 17221 19904 17233 19907
rect 16816 19876 17233 19904
rect 16816 19864 16822 19876
rect 17221 19873 17233 19876
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18598 19904 18604 19916
rect 18371 19876 18604 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 18874 19904 18880 19916
rect 18835 19876 18880 19904
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19978 19904 19984 19916
rect 19939 19876 19984 19904
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 20220 19876 20545 19904
rect 20220 19864 20226 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 10502 19796 10508 19848
rect 10560 19836 10566 19848
rect 10597 19839 10655 19845
rect 10597 19836 10609 19839
rect 10560 19808 10609 19836
rect 10560 19796 10566 19808
rect 10597 19805 10609 19808
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12124 19808 12169 19836
rect 12124 19796 12130 19808
rect 19242 19796 19248 19848
rect 19300 19836 19306 19848
rect 21358 19836 21364 19848
rect 19300 19808 21364 19836
rect 19300 19796 19306 19808
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 9766 19768 9772 19780
rect 9355 19740 9772 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 9766 19728 9772 19740
rect 9824 19728 9830 19780
rect 14001 19771 14059 19777
rect 14001 19737 14013 19771
rect 14047 19768 14059 19771
rect 15286 19768 15292 19780
rect 14047 19740 15292 19768
rect 14047 19737 14059 19740
rect 14001 19731 14059 19737
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 15749 19771 15807 19777
rect 15749 19737 15761 19771
rect 15795 19768 15807 19771
rect 18138 19768 18144 19780
rect 15795 19740 18144 19768
rect 15795 19737 15807 19740
rect 15749 19731 15807 19737
rect 18138 19728 18144 19740
rect 18196 19728 18202 19780
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 12250 19700 12256 19712
rect 11563 19672 12256 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 8588 19468 9720 19496
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 8588 19301 8616 19468
rect 9692 19360 9720 19468
rect 10226 19456 10232 19508
rect 10284 19496 10290 19508
rect 15930 19496 15936 19508
rect 10284 19468 15936 19496
rect 10284 19456 10290 19468
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 9953 19431 10011 19437
rect 9953 19397 9965 19431
rect 9999 19428 10011 19431
rect 10045 19431 10103 19437
rect 10045 19428 10057 19431
rect 9999 19400 10057 19428
rect 9999 19397 10011 19400
rect 9953 19391 10011 19397
rect 10045 19397 10057 19400
rect 10091 19397 10103 19431
rect 10045 19391 10103 19397
rect 16393 19363 16451 19369
rect 9692 19332 10272 19360
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 7800 19264 8585 19292
rect 7800 19252 7806 19264
rect 8573 19261 8585 19264
rect 8619 19261 8631 19295
rect 10134 19292 10140 19304
rect 8573 19255 8631 19261
rect 8772 19264 10140 19292
rect 1946 19184 1952 19236
rect 2004 19224 2010 19236
rect 2958 19224 2964 19236
rect 2004 19196 2964 19224
rect 2004 19184 2010 19196
rect 2958 19184 2964 19196
rect 3016 19184 3022 19236
rect 3050 19184 3056 19236
rect 3108 19224 3114 19236
rect 8772 19224 8800 19264
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 10244 19301 10272 19332
rect 16393 19329 16405 19363
rect 16439 19360 16451 19363
rect 16666 19360 16672 19372
rect 16439 19332 16672 19360
rect 16439 19329 16451 19332
rect 16393 19323 16451 19329
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 10229 19295 10287 19301
rect 10229 19261 10241 19295
rect 10275 19292 10287 19295
rect 10318 19292 10324 19304
rect 10275 19264 10324 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 12158 19292 12164 19304
rect 10704 19264 12164 19292
rect 10704 19236 10732 19264
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14182 19292 14188 19304
rect 14139 19264 14188 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14332 19264 14412 19292
rect 14332 19252 14338 19264
rect 3108 19196 8800 19224
rect 8840 19227 8898 19233
rect 3108 19184 3114 19196
rect 8840 19193 8852 19227
rect 8886 19224 8898 19227
rect 9214 19224 9220 19236
rect 8886 19196 9220 19224
rect 8886 19193 8898 19196
rect 8840 19187 8898 19193
rect 9214 19184 9220 19196
rect 9272 19184 9278 19236
rect 10045 19227 10103 19233
rect 10045 19193 10057 19227
rect 10091 19224 10103 19227
rect 10410 19224 10416 19236
rect 10091 19196 10416 19224
rect 10091 19193 10103 19196
rect 10045 19187 10103 19193
rect 10410 19184 10416 19196
rect 10468 19233 10474 19236
rect 10468 19227 10532 19233
rect 10468 19193 10486 19227
rect 10520 19193 10532 19227
rect 10468 19187 10532 19193
rect 10468 19184 10474 19187
rect 10686 19184 10692 19236
rect 10744 19184 10750 19236
rect 10870 19184 10876 19236
rect 10928 19224 10934 19236
rect 10928 19196 11928 19224
rect 10928 19184 10934 19196
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 8478 19156 8484 19168
rect 1452 19128 8484 19156
rect 1452 19116 1458 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 10778 19156 10784 19168
rect 8628 19128 10784 19156
rect 8628 19116 8634 19128
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11606 19156 11612 19168
rect 11567 19128 11612 19156
rect 11606 19116 11612 19128
rect 11664 19116 11670 19168
rect 11900 19156 11928 19196
rect 11974 19184 11980 19236
rect 12032 19224 12038 19236
rect 12682 19227 12740 19233
rect 12682 19224 12694 19227
rect 12032 19196 12694 19224
rect 12032 19184 12038 19196
rect 12682 19193 12694 19196
rect 12728 19193 12740 19227
rect 12682 19187 12740 19193
rect 13630 19184 13636 19236
rect 13688 19224 13694 19236
rect 14384 19224 14412 19264
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 14516 19264 14749 19292
rect 14516 19252 14522 19264
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 14737 19255 14795 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15562 19292 15568 19304
rect 15059 19264 15568 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 16850 19292 16856 19304
rect 15672 19264 16856 19292
rect 15672 19224 15700 19264
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 17034 19292 17040 19304
rect 16995 19264 17040 19292
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 18233 19295 18291 19301
rect 18233 19261 18245 19295
rect 18279 19292 18291 19295
rect 18414 19292 18420 19304
rect 18279 19264 18420 19292
rect 18279 19261 18291 19264
rect 18233 19255 18291 19261
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19292 18567 19295
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 18555 19264 19073 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 17218 19224 17224 19236
rect 13688 19196 14320 19224
rect 14384 19196 15700 19224
rect 15764 19196 17224 19224
rect 13688 19184 13694 19196
rect 12066 19156 12072 19168
rect 11900 19128 12072 19156
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12342 19116 12348 19168
rect 12400 19156 12406 19168
rect 12526 19156 12532 19168
rect 12400 19128 12532 19156
rect 12400 19116 12406 19128
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13538 19156 13544 19168
rect 13044 19128 13544 19156
rect 13044 19116 13050 19128
rect 13538 19116 13544 19128
rect 13596 19156 13602 19168
rect 14292 19165 14320 19196
rect 15764 19165 15792 19196
rect 17218 19184 17224 19196
rect 17276 19184 17282 19236
rect 17313 19227 17371 19233
rect 17313 19193 17325 19227
rect 17359 19224 17371 19227
rect 18598 19224 18604 19236
rect 17359 19196 18604 19224
rect 17359 19193 17371 19196
rect 17313 19187 17371 19193
rect 18598 19184 18604 19196
rect 18656 19184 18662 19236
rect 18966 19184 18972 19236
rect 19024 19224 19030 19236
rect 19628 19224 19656 19255
rect 19024 19196 19656 19224
rect 19024 19184 19030 19196
rect 19794 19184 19800 19236
rect 19852 19224 19858 19236
rect 20441 19227 20499 19233
rect 20441 19224 20453 19227
rect 19852 19196 20453 19224
rect 19852 19184 19858 19196
rect 20441 19193 20453 19196
rect 20487 19193 20499 19227
rect 20441 19187 20499 19193
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13596 19128 13829 19156
rect 13596 19116 13602 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 13817 19119 13875 19125
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19125 14335 19159
rect 14277 19119 14335 19125
rect 15749 19159 15807 19165
rect 15749 19125 15761 19159
rect 15795 19125 15807 19159
rect 16114 19156 16120 19168
rect 16075 19128 16120 19156
rect 15749 19119 15807 19125
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16206 19116 16212 19168
rect 16264 19156 16270 19168
rect 16264 19128 16309 19156
rect 16264 19116 16270 19128
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 19245 19159 19303 19165
rect 19245 19156 19257 19159
rect 19116 19128 19257 19156
rect 19116 19116 19122 19128
rect 19245 19125 19257 19128
rect 19291 19125 19303 19159
rect 19245 19119 19303 19125
rect 19334 19116 19340 19168
rect 19392 19156 19398 19168
rect 21910 19156 21916 19168
rect 19392 19128 21916 19156
rect 19392 19116 19398 19128
rect 21910 19116 21916 19128
rect 21968 19116 21974 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2958 18912 2964 18964
rect 3016 18952 3022 18964
rect 9214 18952 9220 18964
rect 3016 18924 9076 18952
rect 9175 18924 9220 18952
rect 3016 18912 3022 18924
rect 9048 18884 9076 18924
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 10229 18955 10287 18961
rect 10229 18921 10241 18955
rect 10275 18952 10287 18955
rect 11790 18952 11796 18964
rect 10275 18924 11796 18952
rect 10275 18921 10287 18924
rect 10229 18915 10287 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 11974 18952 11980 18964
rect 11935 18924 11980 18952
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 14274 18952 14280 18964
rect 12216 18924 14280 18952
rect 12216 18912 12222 18924
rect 14274 18912 14280 18924
rect 14332 18912 14338 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 14608 18924 14749 18952
rect 14608 18912 14614 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 14737 18915 14795 18921
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 16482 18952 16488 18964
rect 15988 18924 16488 18952
rect 15988 18912 15994 18924
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 16666 18952 16672 18964
rect 16627 18924 16672 18952
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 16942 18912 16948 18964
rect 17000 18952 17006 18964
rect 17129 18955 17187 18961
rect 17129 18952 17141 18955
rect 17000 18924 17141 18952
rect 17000 18912 17006 18924
rect 17129 18921 17141 18924
rect 17175 18921 17187 18955
rect 17129 18915 17187 18921
rect 17773 18955 17831 18961
rect 17773 18921 17785 18955
rect 17819 18952 17831 18955
rect 17954 18952 17960 18964
rect 17819 18924 17960 18952
rect 17819 18921 17831 18924
rect 17773 18915 17831 18921
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 18509 18955 18567 18961
rect 18509 18921 18521 18955
rect 18555 18952 18567 18955
rect 20898 18952 20904 18964
rect 18555 18924 20904 18952
rect 18555 18921 18567 18924
rect 18509 18915 18567 18921
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 9766 18884 9772 18896
rect 9048 18856 9772 18884
rect 9766 18844 9772 18856
rect 9824 18844 9830 18896
rect 10686 18844 10692 18896
rect 10744 18884 10750 18896
rect 10864 18887 10922 18893
rect 10864 18884 10876 18887
rect 10744 18856 10876 18884
rect 10744 18844 10750 18856
rect 10864 18853 10876 18856
rect 10910 18884 10922 18887
rect 11606 18884 11612 18896
rect 10910 18856 11612 18884
rect 10910 18853 10922 18856
rect 10864 18847 10922 18853
rect 11606 18844 11612 18856
rect 11664 18844 11670 18896
rect 12986 18893 12992 18896
rect 12980 18884 12992 18893
rect 12947 18856 12992 18884
rect 12980 18847 12992 18856
rect 12986 18844 12992 18847
rect 13044 18844 13050 18896
rect 13078 18844 13084 18896
rect 13136 18884 13142 18896
rect 19978 18884 19984 18896
rect 13136 18856 19840 18884
rect 19939 18856 19984 18884
rect 13136 18844 13142 18856
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7800 18788 7849 18816
rect 7800 18776 7806 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 8104 18819 8162 18825
rect 8104 18785 8116 18819
rect 8150 18816 8162 18819
rect 8846 18816 8852 18828
rect 8150 18788 8852 18816
rect 8150 18785 8162 18788
rect 8104 18779 8162 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 9950 18776 9956 18828
rect 10008 18816 10014 18828
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 10008 18788 10057 18816
rect 10008 18776 10014 18788
rect 10045 18785 10057 18788
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 12713 18819 12771 18825
rect 12713 18816 12725 18819
rect 12584 18788 12725 18816
rect 12584 18776 12590 18788
rect 12713 18785 12725 18788
rect 12759 18785 12771 18819
rect 12713 18779 12771 18785
rect 14274 18776 14280 18828
rect 14332 18816 14338 18828
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14332 18788 14565 18816
rect 14332 18776 14338 18788
rect 14553 18785 14565 18788
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 15378 18776 15384 18828
rect 15436 18816 15442 18828
rect 15545 18819 15603 18825
rect 15545 18816 15557 18819
rect 15436 18788 15557 18816
rect 15436 18776 15442 18788
rect 15545 18785 15557 18788
rect 15591 18785 15603 18819
rect 15545 18779 15603 18785
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 15896 18788 16344 18816
rect 15896 18776 15902 18788
rect 10502 18708 10508 18760
rect 10560 18748 10566 18760
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10560 18720 10609 18748
rect 10560 18708 10566 18720
rect 10597 18717 10609 18720
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 15102 18748 15108 18760
rect 13964 18720 15108 18748
rect 13964 18708 13970 18720
rect 15102 18708 15108 18720
rect 15160 18748 15166 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 15160 18720 15301 18748
rect 15160 18708 15166 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 16316 18748 16344 18788
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 16945 18819 17003 18825
rect 16945 18816 16957 18819
rect 16632 18788 16957 18816
rect 16632 18776 16638 18788
rect 16945 18785 16957 18788
rect 16991 18785 17003 18819
rect 16945 18779 17003 18785
rect 17310 18776 17316 18828
rect 17368 18816 17374 18828
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 17368 18788 17601 18816
rect 17368 18776 17374 18788
rect 17589 18785 17601 18788
rect 17635 18785 17647 18819
rect 17589 18779 17647 18785
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18785 19211 18819
rect 19702 18816 19708 18828
rect 19663 18788 19708 18816
rect 19153 18779 19211 18785
rect 18601 18751 18659 18757
rect 18601 18748 18613 18751
rect 16316 18720 18613 18748
rect 15289 18711 15347 18717
rect 18601 18717 18613 18720
rect 18647 18717 18659 18751
rect 18782 18748 18788 18760
rect 18743 18720 18788 18748
rect 18601 18711 18659 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19168 18748 19196 18779
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 19812 18816 19840 18856
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 20254 18816 20260 18828
rect 19812 18788 20260 18816
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 20714 18748 20720 18760
rect 19168 18720 20720 18748
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 290 18640 296 18692
rect 348 18680 354 18692
rect 7650 18680 7656 18692
rect 348 18652 7656 18680
rect 348 18640 354 18652
rect 7650 18640 7656 18652
rect 7708 18640 7714 18692
rect 13924 18652 15148 18680
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 13924 18612 13952 18652
rect 14090 18612 14096 18624
rect 8260 18584 13952 18612
rect 14051 18584 14096 18612
rect 8260 18572 8266 18584
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 15010 18612 15016 18624
rect 14240 18584 15016 18612
rect 14240 18572 14246 18584
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15120 18612 15148 18652
rect 16298 18640 16304 18692
rect 16356 18680 16362 18692
rect 19610 18680 19616 18692
rect 16356 18652 19616 18680
rect 16356 18640 16362 18652
rect 19610 18640 19616 18652
rect 19668 18640 19674 18692
rect 16022 18612 16028 18624
rect 15120 18584 16028 18612
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 17770 18612 17776 18624
rect 16908 18584 17776 18612
rect 16908 18572 16914 18584
rect 17770 18572 17776 18584
rect 17828 18572 17834 18624
rect 18141 18615 18199 18621
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18506 18612 18512 18624
rect 18187 18584 18512 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 19242 18572 19248 18624
rect 19300 18612 19306 18624
rect 19337 18615 19395 18621
rect 19337 18612 19349 18615
rect 19300 18584 19349 18612
rect 19300 18572 19306 18584
rect 19337 18581 19349 18584
rect 19383 18581 19395 18615
rect 19337 18575 19395 18581
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 10502 18408 10508 18420
rect 2556 18380 10508 18408
rect 2556 18368 2562 18380
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 11977 18411 12035 18417
rect 11977 18377 11989 18411
rect 12023 18408 12035 18411
rect 12434 18408 12440 18420
rect 12023 18380 12440 18408
rect 12023 18377 12035 18380
rect 11977 18371 12035 18377
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12621 18411 12679 18417
rect 12621 18377 12633 18411
rect 12667 18408 12679 18411
rect 13078 18408 13084 18420
rect 12667 18380 13084 18408
rect 12667 18377 12679 18380
rect 12621 18371 12679 18377
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 15378 18408 15384 18420
rect 13228 18380 14964 18408
rect 15339 18380 15384 18408
rect 13228 18368 13234 18380
rect 4154 18300 4160 18352
rect 4212 18340 4218 18352
rect 8849 18343 8907 18349
rect 4212 18312 8800 18340
rect 4212 18300 4218 18312
rect 4706 18232 4712 18284
rect 4764 18272 4770 18284
rect 6178 18272 6184 18284
rect 4764 18244 6184 18272
rect 4764 18232 4770 18244
rect 6178 18232 6184 18244
rect 6236 18232 6242 18284
rect 8570 18272 8576 18284
rect 6288 18244 8576 18272
rect 3602 18164 3608 18216
rect 3660 18204 3666 18216
rect 6288 18204 6316 18244
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 8772 18272 8800 18312
rect 8849 18309 8861 18343
rect 8895 18340 8907 18343
rect 10134 18340 10140 18352
rect 8895 18312 10140 18340
rect 8895 18309 8907 18312
rect 8849 18303 8907 18309
rect 10134 18300 10140 18312
rect 10192 18300 10198 18352
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 12897 18343 12955 18349
rect 12897 18340 12909 18343
rect 10284 18312 12909 18340
rect 10284 18300 10290 18312
rect 12897 18309 12909 18312
rect 12943 18309 12955 18343
rect 12897 18303 12955 18309
rect 12989 18343 13047 18349
rect 12989 18309 13001 18343
rect 13035 18340 13047 18343
rect 13998 18340 14004 18352
rect 13035 18312 14004 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 13998 18300 14004 18312
rect 14056 18300 14062 18352
rect 14936 18340 14964 18380
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 15933 18411 15991 18417
rect 15933 18377 15945 18411
rect 15979 18408 15991 18411
rect 16298 18408 16304 18420
rect 15979 18380 16304 18408
rect 15979 18377 15991 18380
rect 15933 18371 15991 18377
rect 16298 18368 16304 18380
rect 16356 18368 16362 18420
rect 17681 18411 17739 18417
rect 17681 18377 17693 18411
rect 17727 18408 17739 18411
rect 18782 18408 18788 18420
rect 17727 18380 18788 18408
rect 17727 18377 17739 18380
rect 17681 18371 17739 18377
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 19150 18368 19156 18420
rect 19208 18408 19214 18420
rect 19337 18411 19395 18417
rect 19337 18408 19349 18411
rect 19208 18380 19349 18408
rect 19208 18368 19214 18380
rect 19337 18377 19349 18380
rect 19383 18377 19395 18411
rect 19337 18371 19395 18377
rect 15838 18340 15844 18352
rect 14936 18312 15844 18340
rect 15838 18300 15844 18312
rect 15896 18300 15902 18352
rect 18049 18343 18107 18349
rect 18049 18309 18061 18343
rect 18095 18340 18107 18343
rect 18095 18312 19748 18340
rect 18095 18309 18107 18312
rect 18049 18303 18107 18309
rect 9030 18272 9036 18284
rect 8772 18244 9036 18272
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 9401 18275 9459 18281
rect 9401 18272 9413 18275
rect 9272 18244 9413 18272
rect 9272 18232 9278 18244
rect 9401 18241 9413 18244
rect 9447 18241 9459 18275
rect 10686 18272 10692 18284
rect 10647 18244 10692 18272
rect 9401 18235 9459 18241
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 10778 18232 10784 18284
rect 10836 18272 10842 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 10836 18244 12265 18272
rect 10836 18232 10842 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 13170 18272 13176 18284
rect 12253 18235 12311 18241
rect 12452 18244 13176 18272
rect 3660 18176 6316 18204
rect 3660 18164 3666 18176
rect 6362 18164 6368 18216
rect 6420 18204 6426 18216
rect 8662 18204 8668 18216
rect 6420 18176 8668 18204
rect 6420 18164 6426 18176
rect 8662 18164 8668 18176
rect 8720 18204 8726 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 8720 18176 9321 18204
rect 8720 18164 8726 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 10042 18164 10048 18216
rect 10100 18204 10106 18216
rect 10413 18207 10471 18213
rect 10413 18204 10425 18207
rect 10100 18176 10425 18204
rect 10100 18164 10106 18176
rect 10413 18173 10425 18176
rect 10459 18173 10471 18207
rect 11054 18204 11060 18216
rect 11015 18176 11060 18204
rect 10413 18167 10471 18173
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18204 11851 18207
rect 11974 18204 11980 18216
rect 11839 18176 11980 18204
rect 11839 18173 11851 18176
rect 11793 18167 11851 18173
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12452 18213 12480 18244
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13446 18272 13452 18284
rect 13407 18244 13452 18272
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 13679 18244 14136 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 14108 18216 14136 18244
rect 15102 18232 15108 18284
rect 15160 18272 15166 18284
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 15160 18244 16313 18272
rect 15160 18232 15166 18244
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 18598 18272 18604 18284
rect 18559 18244 18604 18272
rect 16301 18235 16359 18241
rect 12437 18207 12495 18213
rect 12176 18176 12388 18204
rect 9122 18096 9128 18148
rect 9180 18136 9186 18148
rect 9217 18139 9275 18145
rect 9217 18136 9229 18139
rect 9180 18108 9229 18136
rect 9180 18096 9186 18108
rect 9217 18105 9229 18108
rect 9263 18105 9275 18139
rect 9217 18099 9275 18105
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 10505 18139 10563 18145
rect 10505 18136 10517 18139
rect 9732 18108 10517 18136
rect 9732 18096 9738 18108
rect 10505 18105 10517 18108
rect 10551 18105 10563 18139
rect 10505 18099 10563 18105
rect 11333 18139 11391 18145
rect 11333 18105 11345 18139
rect 11379 18136 11391 18139
rect 12176 18136 12204 18176
rect 11379 18108 12204 18136
rect 12360 18136 12388 18176
rect 12437 18173 12449 18207
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18204 12955 18207
rect 13817 18207 13875 18213
rect 13817 18204 13829 18207
rect 12943 18176 13829 18204
rect 12943 18173 12955 18176
rect 12897 18167 12955 18173
rect 13817 18173 13829 18176
rect 13863 18173 13875 18207
rect 13817 18167 13875 18173
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 13964 18176 14013 18204
rect 13964 18164 13970 18176
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14257 18207 14315 18213
rect 14257 18204 14269 18207
rect 14148 18176 14269 18204
rect 14148 18164 14154 18176
rect 14257 18173 14269 18176
rect 14303 18173 14315 18207
rect 14257 18167 14315 18173
rect 15654 18164 15660 18216
rect 15712 18204 15718 18216
rect 15749 18207 15807 18213
rect 15749 18204 15761 18207
rect 15712 18176 15761 18204
rect 15712 18164 15718 18176
rect 15749 18173 15761 18176
rect 15795 18173 15807 18207
rect 16316 18204 16344 18235
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 16850 18204 16856 18216
rect 16316 18176 16856 18204
rect 15749 18167 15807 18173
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 18417 18207 18475 18213
rect 18417 18173 18429 18207
rect 18463 18204 18475 18207
rect 18506 18204 18512 18216
rect 18463 18176 18512 18204
rect 18463 18173 18475 18176
rect 18417 18167 18475 18173
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 19720 18213 19748 18312
rect 20714 18272 20720 18284
rect 20675 18244 20720 18272
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18173 19211 18207
rect 19153 18167 19211 18173
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 16568 18139 16626 18145
rect 12360 18108 16068 18136
rect 11379 18105 11391 18108
rect 11333 18099 11391 18105
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 7466 18068 7472 18080
rect 5868 18040 7472 18068
rect 5868 18028 5874 18040
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7650 18028 7656 18080
rect 7708 18068 7714 18080
rect 9858 18068 9864 18080
rect 7708 18040 9864 18068
rect 7708 18028 7714 18040
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 10045 18071 10103 18077
rect 10045 18037 10057 18071
rect 10091 18068 10103 18071
rect 10318 18068 10324 18080
rect 10091 18040 10324 18068
rect 10091 18037 10103 18040
rect 10045 18031 10103 18037
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 12253 18071 12311 18077
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 13078 18068 13084 18080
rect 12299 18040 13084 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13357 18071 13415 18077
rect 13357 18068 13369 18071
rect 13320 18040 13369 18068
rect 13320 18028 13326 18040
rect 13357 18037 13369 18040
rect 13403 18037 13415 18071
rect 13357 18031 13415 18037
rect 13817 18071 13875 18077
rect 13817 18037 13829 18071
rect 13863 18068 13875 18071
rect 14182 18068 14188 18080
rect 13863 18040 14188 18068
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 16040 18068 16068 18108
rect 16568 18105 16580 18139
rect 16614 18136 16626 18139
rect 16666 18136 16672 18148
rect 16614 18108 16672 18136
rect 16614 18105 16626 18108
rect 16568 18099 16626 18105
rect 16666 18096 16672 18108
rect 16724 18096 16730 18148
rect 19168 18136 19196 18167
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 20128 18176 20453 18204
rect 20128 18164 20134 18176
rect 20441 18173 20453 18176
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 16776 18108 19196 18136
rect 19981 18139 20039 18145
rect 16776 18068 16804 18108
rect 19981 18105 19993 18139
rect 20027 18136 20039 18139
rect 20530 18136 20536 18148
rect 20027 18108 20536 18136
rect 20027 18105 20039 18108
rect 19981 18099 20039 18105
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 18506 18068 18512 18080
rect 16040 18040 16804 18068
rect 18467 18040 18512 18068
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 7742 17864 7748 17876
rect 7484 17836 7748 17864
rect 7484 17737 7512 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 8846 17864 8852 17876
rect 8807 17836 8852 17864
rect 8846 17824 8852 17836
rect 8904 17864 8910 17876
rect 9490 17864 9496 17876
rect 8904 17836 9496 17864
rect 8904 17824 8910 17836
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 10134 17864 10140 17876
rect 10095 17836 10140 17864
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 10888 17836 12909 17864
rect 9122 17756 9128 17808
rect 9180 17796 9186 17808
rect 10888 17796 10916 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 12897 17827 12955 17833
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13262 17864 13268 17876
rect 13035 17836 13268 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 13630 17864 13636 17876
rect 13495 17836 13636 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 13630 17824 13636 17836
rect 13688 17864 13694 17876
rect 15470 17864 15476 17876
rect 13688 17836 15476 17864
rect 13688 17824 13694 17836
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 15749 17867 15807 17873
rect 15749 17833 15761 17867
rect 15795 17864 15807 17867
rect 16114 17864 16120 17876
rect 15795 17836 16120 17864
rect 15795 17833 15807 17836
rect 15749 17827 15807 17833
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 18506 17824 18512 17876
rect 18564 17864 18570 17876
rect 18785 17867 18843 17873
rect 18785 17864 18797 17867
rect 18564 17836 18797 17864
rect 18564 17824 18570 17836
rect 18785 17833 18797 17836
rect 18831 17833 18843 17867
rect 18785 17827 18843 17833
rect 18966 17824 18972 17876
rect 19024 17864 19030 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 19024 17836 19257 17864
rect 19024 17824 19030 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 20898 17864 20904 17876
rect 20859 17836 20904 17864
rect 19245 17827 19303 17833
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 9180 17768 10916 17796
rect 11977 17799 12035 17805
rect 9180 17756 9186 17768
rect 11977 17765 11989 17799
rect 12023 17796 12035 17799
rect 13170 17796 13176 17808
rect 12023 17768 13176 17796
rect 12023 17765 12035 17768
rect 11977 17759 12035 17765
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 13357 17799 13415 17805
rect 13357 17765 13369 17799
rect 13403 17796 13415 17799
rect 14737 17799 14795 17805
rect 14737 17796 14749 17799
rect 13403 17768 14749 17796
rect 13403 17765 13415 17768
rect 13357 17759 13415 17765
rect 14737 17765 14749 17768
rect 14783 17765 14795 17799
rect 16942 17796 16948 17808
rect 14737 17759 14795 17765
rect 14844 17768 16948 17796
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17697 7527 17731
rect 7469 17691 7527 17697
rect 7736 17731 7794 17737
rect 7736 17697 7748 17731
rect 7782 17728 7794 17731
rect 8294 17728 8300 17740
rect 7782 17700 8300 17728
rect 7782 17697 7794 17700
rect 7736 17691 7794 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 10042 17728 10048 17740
rect 10003 17700 10048 17728
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 10318 17688 10324 17740
rect 10376 17728 10382 17740
rect 10781 17731 10839 17737
rect 10781 17728 10793 17731
rect 10376 17700 10793 17728
rect 10376 17688 10382 17700
rect 10781 17697 10793 17700
rect 10827 17697 10839 17731
rect 10781 17691 10839 17697
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 12618 17728 12624 17740
rect 11931 17700 12624 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 13998 17728 14004 17740
rect 13372 17700 13768 17728
rect 13959 17700 14004 17728
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17660 10287 17663
rect 10410 17660 10416 17672
rect 10275 17632 10416 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 12066 17660 12072 17672
rect 12027 17632 12072 17660
rect 11057 17623 11115 17629
rect 11072 17592 11100 17623
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12526 17660 12532 17672
rect 12487 17632 12532 17660
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 12894 17620 12900 17672
rect 12952 17660 12958 17672
rect 13372 17660 13400 17700
rect 12952 17632 13400 17660
rect 12952 17620 12958 17632
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 13740 17660 13768 17700
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 14844 17728 14872 17768
rect 16942 17756 16948 17768
rect 17000 17756 17006 17808
rect 17218 17756 17224 17808
rect 17276 17796 17282 17808
rect 17276 17768 19840 17796
rect 17276 17756 17282 17768
rect 14108 17700 14872 17728
rect 15289 17731 15347 17737
rect 14108 17660 14136 17700
rect 15289 17697 15301 17731
rect 15335 17728 15347 17731
rect 16117 17731 16175 17737
rect 16117 17728 16129 17731
rect 15335 17700 16129 17728
rect 15335 17697 15347 17700
rect 15289 17691 15347 17697
rect 16117 17697 16129 17700
rect 16163 17697 16175 17731
rect 16117 17691 16175 17697
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17129 17731 17187 17737
rect 17129 17728 17141 17731
rect 16908 17700 17141 17728
rect 16908 17688 16914 17700
rect 17129 17697 17141 17700
rect 17175 17697 17187 17731
rect 17129 17691 17187 17697
rect 17396 17731 17454 17737
rect 17396 17697 17408 17731
rect 17442 17728 17454 17731
rect 18782 17728 18788 17740
rect 17442 17700 18788 17728
rect 17442 17697 17454 17700
rect 17396 17691 17454 17697
rect 18782 17688 18788 17700
rect 18840 17688 18846 17740
rect 19150 17728 19156 17740
rect 19111 17700 19156 17728
rect 19150 17688 19156 17700
rect 19208 17688 19214 17740
rect 19812 17737 19840 17768
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 13596 17632 13641 17660
rect 13740 17632 14136 17660
rect 14277 17663 14335 17669
rect 13596 17620 13602 17632
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 15470 17660 15476 17672
rect 14323 17632 15476 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 16209 17663 16267 17669
rect 16209 17660 16221 17663
rect 15712 17632 16221 17660
rect 15712 17620 15718 17632
rect 16209 17629 16221 17632
rect 16255 17629 16267 17663
rect 16209 17623 16267 17629
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 16356 17632 16405 17660
rect 16356 17620 16362 17632
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 19337 17663 19395 17669
rect 19337 17629 19349 17663
rect 19383 17629 19395 17663
rect 19337 17623 19395 17629
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17629 20039 17663
rect 19981 17623 20039 17629
rect 15194 17592 15200 17604
rect 11072 17564 15200 17592
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 18509 17595 18567 17601
rect 18509 17561 18521 17595
rect 18555 17592 18567 17595
rect 18598 17592 18604 17604
rect 18555 17564 18604 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 18782 17552 18788 17604
rect 18840 17592 18846 17604
rect 19352 17592 19380 17623
rect 18840 17564 19380 17592
rect 18840 17552 18846 17564
rect 842 17484 848 17536
rect 900 17524 906 17536
rect 8478 17524 8484 17536
rect 900 17496 8484 17524
rect 900 17484 906 17496
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 11517 17527 11575 17533
rect 11517 17524 11529 17527
rect 11204 17496 11529 17524
rect 11204 17484 11210 17496
rect 11517 17493 11529 17496
rect 11563 17493 11575 17527
rect 11517 17487 11575 17493
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12342 17524 12348 17536
rect 11756 17496 12348 17524
rect 11756 17484 11762 17496
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 12897 17527 12955 17533
rect 12897 17493 12909 17527
rect 12943 17524 12955 17527
rect 16758 17524 16764 17536
rect 12943 17496 16764 17524
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 16850 17484 16856 17536
rect 16908 17524 16914 17536
rect 17126 17524 17132 17536
rect 16908 17496 17132 17524
rect 16908 17484 16914 17496
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 19996 17524 20024 17623
rect 17460 17496 20024 17524
rect 17460 17484 17466 17496
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 8389 17323 8447 17329
rect 8389 17320 8401 17323
rect 8352 17292 8401 17320
rect 8352 17280 8358 17292
rect 8389 17289 8401 17292
rect 8435 17289 8447 17323
rect 8389 17283 8447 17289
rect 8404 17184 8432 17283
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 12621 17323 12679 17329
rect 9088 17292 10456 17320
rect 9088 17280 9094 17292
rect 8478 17212 8484 17264
rect 8536 17252 8542 17264
rect 8536 17224 10364 17252
rect 8536 17212 8542 17224
rect 8754 17184 8760 17196
rect 8404 17156 8760 17184
rect 8754 17144 8760 17156
rect 8812 17184 8818 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8812 17156 9229 17184
rect 8812 17144 8818 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 9490 17144 9496 17196
rect 9548 17184 9554 17196
rect 10229 17187 10287 17193
rect 10229 17184 10241 17187
rect 9548 17156 10241 17184
rect 9548 17144 9554 17156
rect 10229 17153 10241 17156
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 7742 17116 7748 17128
rect 7055 17088 7748 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8202 17076 8208 17128
rect 8260 17116 8266 17128
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 8260 17088 10149 17116
rect 8260 17076 8266 17088
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 10137 17079 10195 17085
rect 7276 17051 7334 17057
rect 7276 17017 7288 17051
rect 7322 17048 7334 17051
rect 7650 17048 7656 17060
rect 7322 17020 7656 17048
rect 7322 17017 7334 17020
rect 7276 17011 7334 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 8680 17020 10057 17048
rect 8680 16989 8708 17020
rect 10045 17017 10057 17020
rect 10091 17017 10103 17051
rect 10336 17048 10364 17224
rect 10428 17116 10456 17292
rect 12621 17289 12633 17323
rect 12667 17320 12679 17323
rect 13446 17320 13452 17332
rect 12667 17292 13452 17320
rect 12667 17289 12679 17292
rect 12621 17283 12679 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 15654 17320 15660 17332
rect 14476 17292 15660 17320
rect 11977 17255 12035 17261
rect 11256 17224 11928 17252
rect 10502 17144 10508 17196
rect 10560 17184 10566 17196
rect 11149 17187 11207 17193
rect 11149 17184 11161 17187
rect 10560 17156 11161 17184
rect 10560 17144 10566 17156
rect 11149 17153 11161 17156
rect 11195 17153 11207 17187
rect 11149 17147 11207 17153
rect 11057 17119 11115 17125
rect 11057 17116 11069 17119
rect 10428 17088 11069 17116
rect 11057 17085 11069 17088
rect 11103 17116 11115 17119
rect 11256 17116 11284 17224
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 11698 17184 11704 17196
rect 11379 17156 11704 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 11103 17088 11284 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11606 17076 11612 17128
rect 11664 17116 11670 17128
rect 11793 17119 11851 17125
rect 11793 17116 11805 17119
rect 11664 17088 11805 17116
rect 11664 17076 11670 17088
rect 11793 17085 11805 17088
rect 11839 17085 11851 17119
rect 11900 17116 11928 17224
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 12894 17252 12900 17264
rect 12023 17224 12900 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 12894 17212 12900 17224
rect 12952 17212 12958 17264
rect 12986 17212 12992 17264
rect 13044 17252 13050 17264
rect 14476 17252 14504 17292
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 16206 17320 16212 17332
rect 15795 17292 16212 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 16942 17280 16948 17332
rect 17000 17320 17006 17332
rect 19334 17320 19340 17332
rect 17000 17292 19340 17320
rect 17000 17280 17006 17292
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 15286 17252 15292 17264
rect 13044 17224 14504 17252
rect 14568 17224 15292 17252
rect 13044 17212 13050 17224
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12308 17156 13093 17184
rect 12308 17144 12314 17156
rect 13081 17153 13093 17156
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17184 13323 17187
rect 13538 17184 13544 17196
rect 13311 17156 13544 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 14568 17193 14596 17224
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 15381 17255 15439 17261
rect 15381 17221 15393 17255
rect 15427 17252 15439 17255
rect 16758 17252 16764 17264
rect 15427 17224 16764 17252
rect 15427 17221 15439 17224
rect 15381 17215 15439 17221
rect 16758 17212 16764 17224
rect 16816 17212 16822 17264
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 18046 17252 18052 17264
rect 17083 17224 18052 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 16298 17184 16304 17196
rect 16259 17156 16304 17184
rect 14553 17147 14611 17153
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 16540 17156 17264 17184
rect 16540 17144 16546 17156
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 11900 17088 12541 17116
rect 11793 17079 11851 17085
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 12989 17119 13047 17125
rect 12989 17116 13001 17119
rect 12768 17088 13001 17116
rect 12768 17076 12774 17088
rect 12989 17085 13001 17088
rect 13035 17116 13047 17119
rect 15194 17116 15200 17128
rect 13035 17088 14504 17116
rect 15155 17088 15200 17116
rect 13035 17085 13047 17088
rect 12989 17079 13047 17085
rect 14369 17051 14427 17057
rect 14369 17048 14381 17051
rect 10336 17020 14381 17048
rect 10045 17011 10103 17017
rect 14369 17017 14381 17020
rect 14415 17017 14427 17051
rect 14476 17048 14504 17088
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 15528 17088 16865 17116
rect 15528 17076 15534 17088
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 17126 17048 17132 17060
rect 14476 17020 17132 17048
rect 14369 17011 14427 17017
rect 17126 17008 17132 17020
rect 17184 17008 17190 17060
rect 17236 17048 17264 17156
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 20533 17187 20591 17193
rect 20533 17184 20545 17187
rect 19668 17156 20545 17184
rect 19668 17144 19674 17156
rect 20533 17153 20545 17156
rect 20579 17153 20591 17187
rect 20533 17147 20591 17153
rect 17402 17116 17408 17128
rect 17363 17088 17408 17116
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17920 17088 18061 17116
rect 17920 17076 17926 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 18316 17119 18374 17125
rect 18316 17085 18328 17119
rect 18362 17116 18374 17119
rect 18598 17116 18604 17128
rect 18362 17088 18604 17116
rect 18362 17085 18374 17088
rect 18316 17079 18374 17085
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 19886 17116 19892 17128
rect 19444 17088 19892 17116
rect 19444 17048 19472 17088
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 17236 17020 19472 17048
rect 19518 17008 19524 17060
rect 19576 17048 19582 17060
rect 20441 17051 20499 17057
rect 20441 17048 20453 17051
rect 19576 17020 20453 17048
rect 19576 17008 19582 17020
rect 20441 17017 20453 17020
rect 20487 17017 20499 17051
rect 20441 17011 20499 17017
rect 8665 16983 8723 16989
rect 8665 16949 8677 16983
rect 8711 16949 8723 16983
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 8665 16943 8723 16949
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9674 16980 9680 16992
rect 9180 16952 9225 16980
rect 9635 16952 9680 16980
rect 9180 16940 9186 16952
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 10502 16980 10508 16992
rect 9916 16952 10508 16980
rect 9916 16940 9922 16952
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 10686 16980 10692 16992
rect 10647 16952 10692 16980
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 12529 16983 12587 16989
rect 12529 16949 12541 16983
rect 12575 16980 12587 16983
rect 13262 16980 13268 16992
rect 12575 16952 13268 16980
rect 12575 16949 12587 16952
rect 12529 16943 12587 16949
rect 13262 16940 13268 16952
rect 13320 16940 13326 16992
rect 13906 16980 13912 16992
rect 13867 16952 13912 16980
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 14277 16983 14335 16989
rect 14277 16980 14289 16983
rect 14240 16952 14289 16980
rect 14240 16940 14246 16952
rect 14277 16949 14289 16952
rect 14323 16949 14335 16983
rect 14277 16943 14335 16949
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 15528 16952 16129 16980
rect 15528 16940 15534 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 16117 16943 16175 16949
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 16298 16980 16304 16992
rect 16255 16952 16304 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 17954 16980 17960 16992
rect 17635 16952 17960 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 19392 16952 19441 16980
rect 19392 16940 19398 16952
rect 19429 16949 19441 16952
rect 19475 16949 19487 16983
rect 19978 16980 19984 16992
rect 19939 16952 19984 16980
rect 19429 16943 19487 16949
rect 19978 16940 19984 16952
rect 20036 16940 20042 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 6972 16748 7389 16776
rect 6972 16736 6978 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 7377 16739 7435 16745
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 8202 16776 8208 16788
rect 7524 16748 7569 16776
rect 8163 16748 8208 16776
rect 7524 16736 7530 16748
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 9030 16736 9036 16788
rect 9088 16776 9094 16788
rect 9677 16779 9735 16785
rect 9677 16776 9689 16779
rect 9088 16748 9689 16776
rect 9088 16736 9094 16748
rect 9677 16745 9689 16748
rect 9723 16745 9735 16779
rect 10870 16776 10876 16788
rect 9677 16739 9735 16745
rect 10152 16748 10876 16776
rect 8665 16711 8723 16717
rect 8665 16708 8677 16711
rect 7024 16680 8677 16708
rect 7024 16513 7052 16680
rect 8665 16677 8677 16680
rect 8711 16677 8723 16711
rect 10152 16708 10180 16748
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11609 16779 11667 16785
rect 11609 16776 11621 16779
rect 11020 16748 11621 16776
rect 11020 16736 11026 16748
rect 11609 16745 11621 16748
rect 11655 16776 11667 16779
rect 12066 16776 12072 16788
rect 11655 16748 12072 16776
rect 11655 16745 11667 16748
rect 11609 16739 11667 16745
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 13262 16736 13268 16788
rect 13320 16776 13326 16788
rect 14090 16776 14096 16788
rect 13320 16748 14096 16776
rect 13320 16736 13326 16748
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 16942 16776 16948 16788
rect 15335 16748 16948 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 17126 16776 17132 16788
rect 17087 16748 17132 16776
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 18874 16736 18880 16788
rect 18932 16776 18938 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 18932 16748 19625 16776
rect 18932 16736 18938 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 19886 16736 19892 16788
rect 19944 16776 19950 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 19944 16748 20085 16776
rect 19944 16736 19950 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 20073 16739 20131 16745
rect 8665 16671 8723 16677
rect 9232 16680 10180 16708
rect 10244 16680 11928 16708
rect 9232 16652 9260 16680
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 9214 16640 9220 16652
rect 8619 16612 9220 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9490 16640 9496 16652
rect 9451 16612 9496 16640
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 10244 16649 10272 16680
rect 11900 16652 11928 16680
rect 12434 16668 12440 16720
rect 12492 16708 12498 16720
rect 17221 16711 17279 16717
rect 17221 16708 17233 16711
rect 12492 16680 17233 16708
rect 12492 16668 12498 16680
rect 17221 16677 17233 16680
rect 17267 16677 17279 16711
rect 17221 16671 17279 16677
rect 18141 16711 18199 16717
rect 18141 16677 18153 16711
rect 18187 16708 18199 16711
rect 20254 16708 20260 16720
rect 18187 16680 20260 16708
rect 18187 16677 18199 16680
rect 18141 16671 18199 16677
rect 20254 16668 20260 16680
rect 20312 16668 20318 16720
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 9600 16612 10241 16640
rect 7650 16572 7656 16584
rect 7563 16544 7656 16572
rect 7650 16532 7656 16544
rect 7708 16572 7714 16584
rect 8202 16572 8208 16584
rect 7708 16544 8208 16572
rect 7708 16532 7714 16544
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8754 16572 8760 16584
rect 8715 16544 8760 16572
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 9600 16572 9628 16612
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 10496 16643 10554 16649
rect 10496 16609 10508 16643
rect 10542 16640 10554 16643
rect 11698 16640 11704 16652
rect 10542 16612 11704 16640
rect 10542 16609 10554 16612
rect 10496 16603 10554 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 12152 16643 12210 16649
rect 11940 16612 12033 16640
rect 11940 16600 11946 16612
rect 12152 16609 12164 16643
rect 12198 16640 12210 16643
rect 12894 16640 12900 16652
rect 12198 16612 12900 16640
rect 12198 16609 12210 16612
rect 12152 16603 12210 16609
rect 12894 16600 12900 16612
rect 12952 16600 12958 16652
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13630 16640 13636 16652
rect 13587 16612 13636 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 13808 16643 13866 16649
rect 13808 16609 13820 16643
rect 13854 16640 13866 16643
rect 15286 16640 15292 16652
rect 13854 16612 15292 16640
rect 13854 16609 13866 16612
rect 13808 16603 13866 16609
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 15620 16612 15976 16640
rect 15620 16600 15626 16612
rect 15194 16572 15200 16584
rect 9324 16544 9628 16572
rect 14559 16544 15200 16572
rect 7009 16507 7067 16513
rect 7009 16473 7021 16507
rect 7055 16473 7067 16507
rect 7009 16467 7067 16473
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 9324 16513 9352 16544
rect 9309 16507 9367 16513
rect 9309 16504 9321 16507
rect 7800 16476 9321 16504
rect 7800 16464 7806 16476
rect 9309 16473 9321 16476
rect 9355 16504 9367 16507
rect 9398 16504 9404 16516
rect 9355 16476 9404 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 13262 16436 13268 16448
rect 13223 16408 13268 16436
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 14559 16436 14587 16544
rect 15194 16532 15200 16544
rect 15252 16572 15258 16584
rect 15746 16572 15752 16584
rect 15252 16544 15752 16572
rect 15252 16532 15258 16544
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 15948 16572 15976 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 16080 16612 16129 16640
rect 16080 16600 16086 16612
rect 16117 16609 16129 16612
rect 16163 16640 16175 16643
rect 17586 16640 17592 16652
rect 16163 16612 17592 16640
rect 16163 16609 16175 16612
rect 16117 16603 16175 16609
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 17862 16640 17868 16652
rect 17823 16612 17868 16640
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 18969 16643 19027 16649
rect 18969 16640 18981 16643
rect 18564 16612 18981 16640
rect 18564 16600 18570 16612
rect 18969 16609 18981 16612
rect 19015 16609 19027 16643
rect 18969 16603 19027 16609
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19484 16612 19993 16640
rect 19484 16600 19490 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 16206 16572 16212 16584
rect 15948 16544 16212 16572
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16572 16451 16575
rect 17310 16572 17316 16584
rect 16439 16544 17316 16572
rect 16439 16541 16451 16544
rect 16393 16535 16451 16541
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 16408 16504 16436 16535
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 19061 16575 19119 16581
rect 19061 16572 19073 16575
rect 17736 16544 19073 16572
rect 17736 16532 17742 16544
rect 19061 16541 19073 16544
rect 19107 16541 19119 16575
rect 19061 16535 19119 16541
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16572 19303 16575
rect 19334 16572 19340 16584
rect 19291 16544 19340 16572
rect 19291 16541 19303 16544
rect 19245 16535 19303 16541
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 20165 16575 20223 16581
rect 20165 16541 20177 16575
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 15344 16476 16436 16504
rect 15344 16464 15350 16476
rect 16482 16464 16488 16516
rect 16540 16504 16546 16516
rect 19352 16504 19380 16532
rect 20180 16504 20208 16535
rect 16540 16476 18736 16504
rect 19352 16476 20208 16504
rect 16540 16464 16546 16476
rect 13412 16408 14587 16436
rect 14921 16439 14979 16445
rect 13412 16396 13418 16408
rect 14921 16405 14933 16439
rect 14967 16436 14979 16439
rect 15010 16436 15016 16448
rect 14967 16408 15016 16436
rect 14967 16405 14979 16408
rect 14921 16399 14979 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 15746 16436 15752 16448
rect 15707 16408 15752 16436
rect 15746 16396 15752 16408
rect 15804 16396 15810 16448
rect 15838 16396 15844 16448
rect 15896 16436 15902 16448
rect 16761 16439 16819 16445
rect 16761 16436 16773 16439
rect 15896 16408 16773 16436
rect 15896 16396 15902 16408
rect 16761 16405 16773 16408
rect 16807 16405 16819 16439
rect 18598 16436 18604 16448
rect 18559 16408 18604 16436
rect 16761 16399 16819 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 18708 16436 18736 16476
rect 20714 16436 20720 16448
rect 18708 16408 20720 16436
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 8202 16232 8208 16244
rect 8163 16204 8208 16232
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9674 16232 9680 16244
rect 9232 16204 9680 16232
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 6914 16028 6920 16040
rect 6871 16000 6920 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 6914 15988 6920 16000
rect 6972 16028 6978 16040
rect 7650 16028 7656 16040
rect 6972 16000 7656 16028
rect 6972 15988 6978 16000
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 9232 16028 9260 16204
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 12250 16232 12256 16244
rect 11532 16204 12256 16232
rect 9398 16096 9404 16108
rect 9359 16068 9404 16096
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11532 16105 11560 16204
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12618 16232 12624 16244
rect 12483 16204 12624 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 14274 16192 14280 16244
rect 14332 16232 14338 16244
rect 16485 16235 16543 16241
rect 14332 16204 16344 16232
rect 14332 16192 14338 16204
rect 12158 16124 12164 16176
rect 12216 16164 12222 16176
rect 12710 16164 12716 16176
rect 12216 16136 12716 16164
rect 12216 16124 12222 16136
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 13630 16124 13636 16176
rect 13688 16164 13694 16176
rect 13688 16136 14044 16164
rect 13688 16124 13694 16136
rect 14016 16108 14044 16136
rect 15010 16124 15016 16176
rect 15068 16164 15074 16176
rect 15068 16136 16252 16164
rect 15068 16124 15074 16136
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 10928 16068 11529 16096
rect 10928 16056 10934 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11698 16096 11704 16108
rect 11611 16068 11704 16096
rect 11517 16059 11575 16065
rect 11698 16056 11704 16068
rect 11756 16096 11762 16108
rect 13081 16099 13139 16105
rect 13081 16096 13093 16099
rect 11756 16068 13093 16096
rect 11756 16056 11762 16068
rect 13081 16065 13093 16068
rect 13127 16096 13139 16099
rect 13262 16096 13268 16108
rect 13127 16068 13268 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13262 16056 13268 16068
rect 13320 16096 13326 16108
rect 13722 16096 13728 16108
rect 13320 16068 13728 16096
rect 13320 16056 13326 16068
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 13998 16096 14004 16108
rect 13959 16068 14004 16096
rect 13998 16056 14004 16068
rect 14056 16056 14062 16108
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 16224 16105 16252 16136
rect 16117 16099 16175 16105
rect 16117 16096 16129 16099
rect 15804 16068 16129 16096
rect 15804 16056 15810 16068
rect 16117 16065 16129 16068
rect 16163 16065 16175 16099
rect 16117 16059 16175 16065
rect 16209 16099 16267 16105
rect 16209 16065 16221 16099
rect 16255 16065 16267 16099
rect 16316 16096 16344 16204
rect 16485 16201 16497 16235
rect 16531 16232 16543 16235
rect 20714 16232 20720 16244
rect 16531 16204 20720 16232
rect 16531 16201 16543 16204
rect 16485 16195 16543 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 17129 16099 17187 16105
rect 17129 16096 17141 16099
rect 16316 16068 17141 16096
rect 16209 16059 16267 16065
rect 17129 16065 17141 16068
rect 17175 16065 17187 16099
rect 17310 16096 17316 16108
rect 17271 16068 17316 16096
rect 17129 16059 17187 16065
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 19886 16056 19892 16108
rect 19944 16096 19950 16108
rect 20349 16099 20407 16105
rect 20349 16096 20361 16099
rect 19944 16068 20361 16096
rect 19944 16056 19950 16068
rect 20349 16065 20361 16068
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 8711 16000 9260 16028
rect 9324 16000 12480 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 8846 15960 8852 15972
rect 7138 15932 8852 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 8941 15963 8999 15969
rect 8941 15929 8953 15963
rect 8987 15960 8999 15963
rect 9324 15960 9352 16000
rect 8987 15932 9352 15960
rect 9668 15963 9726 15969
rect 8987 15929 8999 15932
rect 8941 15923 8999 15929
rect 9668 15929 9680 15963
rect 9714 15960 9726 15963
rect 10962 15960 10968 15972
rect 9714 15932 10968 15960
rect 9714 15929 9726 15932
rect 9668 15923 9726 15929
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 11425 15963 11483 15969
rect 11425 15929 11437 15963
rect 11471 15960 11483 15963
rect 12158 15960 12164 15972
rect 11471 15932 12164 15960
rect 11471 15929 11483 15932
rect 11425 15923 11483 15929
rect 12158 15920 12164 15932
rect 12216 15920 12222 15972
rect 12452 15960 12480 16000
rect 12526 15988 12532 16040
rect 12584 16028 12590 16040
rect 12805 16031 12863 16037
rect 12805 16028 12817 16031
rect 12584 16000 12817 16028
rect 12584 15988 12590 16000
rect 12805 15997 12817 16000
rect 12851 15997 12863 16031
rect 12805 15991 12863 15997
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 16028 12955 16031
rect 13354 16028 13360 16040
rect 12943 16000 13360 16028
rect 12943 15997 12955 16000
rect 12897 15991 12955 15997
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 13449 16031 13507 16037
rect 13449 15997 13461 16031
rect 13495 16028 13507 16031
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 13495 16000 13921 16028
rect 13495 15997 13507 16000
rect 13449 15991 13507 15997
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 14016 16000 16804 16028
rect 14016 15960 14044 16000
rect 12452 15932 14044 15960
rect 14268 15963 14326 15969
rect 14268 15929 14280 15963
rect 14314 15960 14326 15963
rect 15010 15960 15016 15972
rect 14314 15932 15016 15960
rect 14314 15929 14326 15932
rect 14268 15923 14326 15929
rect 15010 15920 15016 15932
rect 15068 15920 15074 15972
rect 16025 15963 16083 15969
rect 15212 15932 15976 15960
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11054 15892 11060 15904
rect 11015 15864 11060 15892
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 12986 15892 12992 15904
rect 12308 15864 12992 15892
rect 12308 15852 12314 15864
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 13630 15892 13636 15904
rect 13591 15864 13636 15892
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 13909 15895 13967 15901
rect 13909 15861 13921 15895
rect 13955 15892 13967 15895
rect 15212 15892 15240 15932
rect 15378 15892 15384 15904
rect 13955 15864 15240 15892
rect 15339 15864 15384 15892
rect 13955 15861 13967 15864
rect 13909 15855 13967 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 15654 15892 15660 15904
rect 15615 15864 15660 15892
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 15948 15892 15976 15932
rect 16025 15929 16037 15963
rect 16071 15960 16083 15963
rect 16776 15960 16804 16000
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17037 16031 17095 16037
rect 17037 16028 17049 16031
rect 17000 16000 17049 16028
rect 17000 15988 17006 16000
rect 17037 15997 17049 16000
rect 17083 15997 17095 16031
rect 17037 15991 17095 15997
rect 17678 15988 17684 16040
rect 17736 16028 17742 16040
rect 17865 16031 17923 16037
rect 17865 16028 17877 16031
rect 17736 16000 17877 16028
rect 17736 15988 17742 16000
rect 17865 15997 17877 16000
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 18012 16000 18061 16028
rect 18012 15988 18018 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 20809 16031 20867 16037
rect 20809 16028 20821 16031
rect 18049 15991 18107 15997
rect 18156 16000 20821 16028
rect 18156 15960 18184 16000
rect 20809 15997 20821 16000
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 16071 15932 16712 15960
rect 16776 15932 18184 15960
rect 18316 15963 18374 15969
rect 16071 15929 16083 15932
rect 16025 15923 16083 15929
rect 16684 15901 16712 15932
rect 18316 15929 18328 15963
rect 18362 15960 18374 15963
rect 19334 15960 19340 15972
rect 18362 15932 19340 15960
rect 18362 15929 18374 15932
rect 18316 15923 18374 15929
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 20162 15960 20168 15972
rect 20123 15932 20168 15960
rect 20162 15920 20168 15932
rect 20220 15920 20226 15972
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15960 20315 15963
rect 20898 15960 20904 15972
rect 20303 15932 20904 15960
rect 20303 15929 20315 15932
rect 20257 15923 20315 15929
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 16485 15895 16543 15901
rect 16485 15892 16497 15895
rect 15948 15864 16497 15892
rect 16485 15861 16497 15864
rect 16531 15861 16543 15895
rect 16485 15855 16543 15861
rect 16669 15895 16727 15901
rect 16669 15861 16681 15895
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 17681 15895 17739 15901
rect 17681 15861 17693 15895
rect 17727 15892 17739 15895
rect 17954 15892 17960 15904
rect 17727 15864 17960 15892
rect 17727 15861 17739 15864
rect 17681 15855 17739 15861
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 18782 15852 18788 15904
rect 18840 15892 18846 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 18840 15864 19441 15892
rect 18840 15852 18846 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 19794 15892 19800 15904
rect 19755 15864 19800 15892
rect 19429 15855 19487 15861
rect 19794 15852 19800 15864
rect 19852 15852 19858 15904
rect 20990 15892 20996 15904
rect 20951 15864 20996 15892
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 8772 15660 10333 15688
rect 6448 15623 6506 15629
rect 6448 15589 6460 15623
rect 6494 15620 6506 15623
rect 8772 15620 8800 15660
rect 10321 15657 10333 15660
rect 10367 15657 10379 15691
rect 10321 15651 10379 15657
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15657 10471 15691
rect 10413 15651 10471 15657
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 11330 15688 11336 15700
rect 10827 15660 11336 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 10428 15620 10456 15651
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 13170 15688 13176 15700
rect 13131 15660 13176 15688
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14093 15691 14151 15697
rect 14093 15688 14105 15691
rect 13964 15660 14105 15688
rect 13964 15648 13970 15660
rect 14093 15657 14105 15660
rect 14139 15657 14151 15691
rect 14093 15651 14151 15657
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 15252 15660 15301 15688
rect 15252 15648 15258 15660
rect 15289 15657 15301 15660
rect 15335 15657 15347 15691
rect 15654 15688 15660 15700
rect 15615 15660 15660 15688
rect 15289 15651 15347 15657
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 17310 15648 17316 15700
rect 17368 15688 17374 15700
rect 17773 15691 17831 15697
rect 17773 15688 17785 15691
rect 17368 15660 17785 15688
rect 17368 15648 17374 15660
rect 17773 15657 17785 15660
rect 17819 15657 17831 15691
rect 17773 15651 17831 15657
rect 18049 15691 18107 15697
rect 18049 15657 18061 15691
rect 18095 15688 18107 15691
rect 19426 15688 19432 15700
rect 18095 15660 19432 15688
rect 18095 15657 18107 15660
rect 18049 15651 18107 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 11882 15620 11888 15632
rect 6494 15592 8800 15620
rect 8864 15592 10456 15620
rect 11532 15592 11888 15620
rect 6494 15589 6506 15592
rect 6448 15583 6506 15589
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 6914 15552 6920 15564
rect 6227 15524 6920 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 8864 15561 8892 15592
rect 8849 15555 8907 15561
rect 8849 15521 8861 15555
rect 8895 15521 8907 15555
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 8849 15515 8907 15521
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 10134 15552 10140 15564
rect 9824 15524 10140 15552
rect 9824 15512 9830 15524
rect 10134 15512 10140 15524
rect 10192 15512 10198 15564
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 10778 15552 10784 15564
rect 10367 15524 10784 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10778 15512 10784 15524
rect 10836 15552 10842 15564
rect 11532 15561 11560 15592
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 14553 15623 14611 15629
rect 14553 15589 14565 15623
rect 14599 15620 14611 15623
rect 15838 15620 15844 15632
rect 14599 15592 15844 15620
rect 14599 15589 14611 15592
rect 14553 15583 14611 15589
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 17954 15620 17960 15632
rect 16408 15592 17960 15620
rect 11790 15561 11796 15564
rect 11517 15555 11575 15561
rect 10836 15524 11008 15552
rect 10836 15512 10842 15524
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9858 15484 9864 15496
rect 9171 15456 9864 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15453 10011 15487
rect 10870 15484 10876 15496
rect 10831 15456 10876 15484
rect 9953 15447 10011 15453
rect 7558 15348 7564 15360
rect 7519 15320 7564 15348
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 9968 15348 9996 15447
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 10980 15493 11008 15524
rect 11517 15521 11529 15555
rect 11563 15521 11575 15555
rect 11517 15515 11575 15521
rect 11784 15515 11796 15561
rect 11848 15552 11854 15564
rect 13541 15555 13599 15561
rect 11848 15524 11884 15552
rect 11790 15512 11796 15515
rect 11848 15512 11854 15524
rect 13541 15521 13553 15555
rect 13587 15552 13599 15555
rect 13587 15524 15240 15552
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15453 11023 15487
rect 13630 15484 13636 15496
rect 13591 15456 13636 15484
rect 10965 15447 11023 15453
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 13722 15444 13728 15496
rect 13780 15484 13786 15496
rect 14093 15487 14151 15493
rect 13780 15456 13825 15484
rect 13780 15444 13786 15456
rect 14093 15453 14105 15487
rect 14139 15484 14151 15487
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14139 15456 14657 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 15010 15484 15016 15496
rect 14875 15456 15016 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 15212 15484 15240 15524
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15436 15524 15884 15552
rect 15436 15512 15442 15524
rect 15654 15484 15660 15496
rect 15212 15456 15660 15484
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 15856 15493 15884 15524
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 15841 15487 15899 15493
rect 15841 15453 15853 15487
rect 15887 15453 15899 15487
rect 15841 15447 15899 15453
rect 14185 15419 14243 15425
rect 12728 15388 13032 15416
rect 12728 15348 12756 15388
rect 12894 15348 12900 15360
rect 9968 15320 12756 15348
rect 12855 15320 12900 15348
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13004 15348 13032 15388
rect 14185 15385 14197 15419
rect 14231 15416 14243 15419
rect 15764 15416 15792 15447
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 16408 15493 16436 15592
rect 17954 15580 17960 15592
rect 18012 15620 18018 15632
rect 18782 15629 18788 15632
rect 18776 15620 18788 15629
rect 18012 15592 18552 15620
rect 18743 15592 18788 15620
rect 18012 15580 18018 15592
rect 16660 15555 16718 15561
rect 16660 15521 16672 15555
rect 16706 15552 16718 15555
rect 17494 15552 17500 15564
rect 16706 15524 17500 15552
rect 16706 15521 16718 15524
rect 16660 15515 16718 15521
rect 17494 15512 17500 15524
rect 17552 15512 17558 15564
rect 18524 15561 18552 15592
rect 18776 15583 18788 15592
rect 18782 15580 18788 15583
rect 18840 15580 18846 15632
rect 18509 15555 18567 15561
rect 18509 15521 18521 15555
rect 18555 15521 18567 15555
rect 20254 15552 20260 15564
rect 18509 15515 18567 15521
rect 18616 15524 19840 15552
rect 20215 15524 20260 15552
rect 16393 15487 16451 15493
rect 16393 15484 16405 15487
rect 16172 15456 16405 15484
rect 16172 15444 16178 15456
rect 16393 15453 16405 15456
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 17770 15444 17776 15496
rect 17828 15484 17834 15496
rect 18616 15484 18644 15524
rect 17828 15456 18644 15484
rect 19812 15484 19840 15524
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 20898 15484 20904 15496
rect 19812 15456 20904 15484
rect 17828 15444 17834 15456
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 14231 15388 15792 15416
rect 14231 15385 14243 15388
rect 14185 15379 14243 15385
rect 17402 15348 17408 15360
rect 13004 15320 17408 15348
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 17586 15308 17592 15360
rect 17644 15348 17650 15360
rect 20162 15348 20168 15360
rect 17644 15320 20168 15348
rect 17644 15308 17650 15320
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 5767 15116 9812 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 8846 15036 8852 15088
rect 8904 15076 8910 15088
rect 9030 15076 9036 15088
rect 8904 15048 9036 15076
rect 8904 15036 8910 15048
rect 9030 15036 9036 15048
rect 9088 15036 9094 15088
rect 6178 15008 6184 15020
rect 6139 14980 6184 15008
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 7558 15008 7564 15020
rect 6411 14980 7564 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 9784 15017 9812 15116
rect 9858 15104 9864 15156
rect 9916 15104 9922 15156
rect 10321 15147 10379 15153
rect 10321 15113 10333 15147
rect 10367 15144 10379 15147
rect 10870 15144 10876 15156
rect 10367 15116 10876 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 10980 15116 16160 15144
rect 9876 15076 9904 15104
rect 10980 15076 11008 15116
rect 9876 15048 11008 15076
rect 12805 15079 12863 15085
rect 12805 15045 12817 15079
rect 12851 15076 12863 15079
rect 12851 15048 13952 15076
rect 12851 15045 12863 15048
rect 12805 15039 12863 15045
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 9858 14968 9864 15020
rect 9916 15008 9922 15020
rect 9916 14980 9961 15008
rect 9916 14968 9922 14980
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10744 14980 10793 15008
rect 10744 14968 10750 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10962 15008 10968 15020
rect 10923 14980 10968 15008
rect 10781 14971 10839 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 11885 15011 11943 15017
rect 11885 15008 11897 15011
rect 11848 14980 11897 15008
rect 11848 14968 11854 14980
rect 11885 14977 11897 14980
rect 11931 15008 11943 15011
rect 12342 15008 12348 15020
rect 11931 14980 12348 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12342 14968 12348 14980
rect 12400 15008 12406 15020
rect 13633 15011 13691 15017
rect 13633 15008 13645 15011
rect 12400 14980 13645 15008
rect 12400 14968 12406 14980
rect 13633 14977 13645 14980
rect 13679 14977 13691 15011
rect 13633 14971 13691 14977
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6086 14940 6092 14952
rect 5592 14912 6092 14940
rect 5592 14900 5598 14912
rect 6086 14900 6092 14912
rect 6144 14900 6150 14952
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 7920 14943 7978 14949
rect 7920 14909 7932 14943
rect 7966 14940 7978 14943
rect 9876 14940 9904 14968
rect 7966 14912 9904 14940
rect 7966 14909 7978 14912
rect 7920 14903 7978 14909
rect 6822 14832 6828 14884
rect 6880 14872 6886 14884
rect 7668 14872 7696 14903
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 12710 14940 12716 14952
rect 11572 14912 12716 14940
rect 11572 14900 11578 14912
rect 12710 14900 12716 14912
rect 12768 14940 12774 14952
rect 12989 14943 13047 14949
rect 12989 14940 13001 14943
rect 12768 14912 13001 14940
rect 12768 14900 12774 14912
rect 12989 14909 13001 14912
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 9766 14872 9772 14884
rect 6880 14844 9772 14872
rect 6880 14832 6886 14844
rect 9766 14832 9772 14844
rect 9824 14832 9830 14884
rect 10689 14875 10747 14881
rect 10689 14841 10701 14875
rect 10735 14872 10747 14875
rect 11054 14872 11060 14884
rect 10735 14844 11060 14872
rect 10735 14841 10747 14844
rect 10689 14835 10747 14841
rect 11054 14832 11060 14844
rect 11112 14832 11118 14884
rect 13722 14872 13728 14884
rect 11348 14844 13728 14872
rect 9306 14804 9312 14816
rect 9267 14776 9312 14804
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 9677 14807 9735 14813
rect 9677 14773 9689 14807
rect 9723 14804 9735 14807
rect 10226 14804 10232 14816
rect 9723 14776 10232 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 11348 14813 11376 14844
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 13924 14872 13952 15048
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 14056 14980 14289 15008
rect 14056 14968 14062 14980
rect 14277 14977 14289 14980
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 15470 15008 15476 15020
rect 15344 14980 15476 15008
rect 15344 14968 15350 14980
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 14544 14943 14602 14949
rect 14544 14909 14556 14943
rect 14590 14940 14602 14943
rect 15378 14940 15384 14952
rect 14590 14912 15384 14940
rect 14590 14909 14602 14912
rect 14544 14903 14602 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 16132 14949 16160 15116
rect 17862 15104 17868 15156
rect 17920 15144 17926 15156
rect 18509 15147 18567 15153
rect 18509 15144 18521 15147
rect 17920 15116 18521 15144
rect 17920 15104 17926 15116
rect 18509 15113 18521 15116
rect 18555 15113 18567 15147
rect 18509 15107 18567 15113
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 20070 15144 20076 15156
rect 19659 15116 20076 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 20806 15144 20812 15156
rect 20767 15116 20812 15144
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 17034 15036 17040 15088
rect 17092 15076 17098 15088
rect 19702 15076 19708 15088
rect 17092 15048 19708 15076
rect 17092 15036 17098 15048
rect 19702 15036 19708 15048
rect 19760 15036 19766 15088
rect 19886 15036 19892 15088
rect 19944 15076 19950 15088
rect 20346 15076 20352 15088
rect 19944 15048 20352 15076
rect 19944 15036 19950 15048
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 16390 14968 16396 15020
rect 16448 15008 16454 15020
rect 16850 15008 16856 15020
rect 16448 14980 16856 15008
rect 16448 14968 16454 14980
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 17218 15008 17224 15020
rect 17179 14980 17224 15008
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 18782 14968 18788 15020
rect 18840 15008 18846 15020
rect 19061 15011 19119 15017
rect 19061 15008 19073 15011
rect 18840 14980 19073 15008
rect 18840 14968 18846 14980
rect 19061 14977 19073 14980
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19852 14980 20085 15008
rect 19852 14968 19858 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 15008 20315 15011
rect 20438 15008 20444 15020
rect 20303 14980 20444 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14909 16175 14943
rect 16482 14940 16488 14952
rect 16117 14903 16175 14909
rect 16316 14912 16488 14940
rect 16316 14872 16344 14912
rect 16482 14900 16488 14912
rect 16540 14940 16546 14952
rect 17678 14940 17684 14952
rect 16540 14912 17684 14940
rect 16540 14900 16546 14912
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 18874 14940 18880 14952
rect 18835 14912 18880 14940
rect 18874 14900 18880 14912
rect 18932 14900 18938 14952
rect 20530 14900 20536 14952
rect 20588 14940 20594 14952
rect 20625 14943 20683 14949
rect 20625 14940 20637 14943
rect 20588 14912 20637 14940
rect 20588 14900 20594 14912
rect 20625 14909 20637 14912
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 13924 14844 16344 14872
rect 16390 14832 16396 14884
rect 16448 14872 16454 14884
rect 17037 14875 17095 14881
rect 17037 14872 17049 14875
rect 16448 14844 17049 14872
rect 16448 14832 16454 14844
rect 17037 14841 17049 14844
rect 17083 14841 17095 14875
rect 17037 14835 17095 14841
rect 18598 14832 18604 14884
rect 18656 14872 18662 14884
rect 18969 14875 19027 14881
rect 18969 14872 18981 14875
rect 18656 14844 18981 14872
rect 18656 14832 18662 14844
rect 18969 14841 18981 14844
rect 19015 14841 19027 14875
rect 18969 14835 19027 14841
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14773 11391 14807
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11333 14767 11391 14773
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 13078 14804 13084 14816
rect 11848 14776 11893 14804
rect 13039 14776 13084 14804
rect 11848 14764 11854 14776
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13446 14804 13452 14816
rect 13407 14776 13452 14804
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13541 14807 13599 14813
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 14550 14804 14556 14816
rect 13587 14776 14556 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15344 14776 15669 14804
rect 15344 14764 15350 14776
rect 15657 14773 15669 14776
rect 15703 14773 15715 14807
rect 16298 14804 16304 14816
rect 16259 14776 16304 14804
rect 15657 14767 15715 14773
rect 16298 14764 16304 14776
rect 16356 14764 16362 14816
rect 16666 14804 16672 14816
rect 16627 14776 16672 14804
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17126 14804 17132 14816
rect 17087 14776 17132 14804
rect 17126 14764 17132 14776
rect 17184 14764 17190 14816
rect 18874 14764 18880 14816
rect 18932 14804 18938 14816
rect 19610 14804 19616 14816
rect 18932 14776 19616 14804
rect 18932 14764 18938 14776
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 19978 14804 19984 14816
rect 19939 14776 19984 14804
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 8481 14603 8539 14609
rect 8481 14569 8493 14603
rect 8527 14569 8539 14603
rect 8481 14563 8539 14569
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9306 14600 9312 14612
rect 8987 14572 9312 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 7092 14535 7150 14541
rect 7092 14501 7104 14535
rect 7138 14532 7150 14535
rect 7558 14532 7564 14544
rect 7138 14504 7564 14532
rect 7138 14501 7150 14504
rect 7092 14495 7150 14501
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 8496 14532 8524 14563
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 11333 14603 11391 14609
rect 11333 14600 11345 14603
rect 9548 14572 11345 14600
rect 9548 14560 9554 14572
rect 11333 14569 11345 14572
rect 11379 14569 11391 14603
rect 11333 14563 11391 14569
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12400 14572 13001 14600
rect 12400 14560 12406 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 13136 14572 13645 14600
rect 13136 14560 13142 14572
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13633 14563 13691 14569
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 13780 14572 13825 14600
rect 13780 14560 13786 14572
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 16114 14600 16120 14612
rect 14056 14572 16120 14600
rect 14056 14560 14062 14572
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 17494 14600 17500 14612
rect 17455 14572 17500 14600
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 17586 14560 17592 14612
rect 17644 14600 17650 14612
rect 18506 14600 18512 14612
rect 17644 14572 18512 14600
rect 17644 14560 17650 14572
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 20438 14600 20444 14612
rect 20399 14572 20444 14600
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 9674 14532 9680 14544
rect 8496 14504 9680 14532
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 9944 14535 10002 14541
rect 9944 14501 9956 14535
rect 9990 14532 10002 14535
rect 13262 14532 13268 14544
rect 9990 14504 13268 14532
rect 9990 14501 10002 14504
rect 9944 14495 10002 14501
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 14553 14535 14611 14541
rect 14553 14532 14565 14535
rect 14424 14504 14565 14532
rect 14424 14492 14430 14504
rect 14553 14501 14565 14504
rect 14599 14501 14611 14535
rect 14553 14495 14611 14501
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 16384 14535 16442 14541
rect 15252 14504 15332 14532
rect 15252 14492 15258 14504
rect 6822 14464 6828 14476
rect 6783 14436 6828 14464
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 8849 14467 8907 14473
rect 8849 14464 8861 14467
rect 8536 14436 8861 14464
rect 8536 14424 8542 14436
rect 8849 14433 8861 14436
rect 8895 14433 8907 14467
rect 9766 14464 9772 14476
rect 9679 14436 9772 14464
rect 8849 14427 8907 14433
rect 9692 14408 9720 14436
rect 9766 14424 9772 14436
rect 9824 14464 9830 14476
rect 11514 14464 11520 14476
rect 9824 14436 10732 14464
rect 11475 14436 11520 14464
rect 9824 14424 9830 14436
rect 9030 14396 9036 14408
rect 8991 14368 9036 14396
rect 9030 14356 9036 14368
rect 9088 14356 9094 14408
rect 9674 14396 9680 14408
rect 9587 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 10704 14396 10732 14436
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 11882 14473 11888 14476
rect 11876 14427 11888 14473
rect 11940 14464 11946 14476
rect 15304 14473 15332 14504
rect 16384 14501 16396 14535
rect 16430 14532 16442 14535
rect 17218 14532 17224 14544
rect 16430 14504 17224 14532
rect 16430 14501 16442 14504
rect 16384 14495 16442 14501
rect 17218 14492 17224 14504
rect 17276 14532 17282 14544
rect 17276 14504 18276 14532
rect 17276 14492 17282 14504
rect 14277 14467 14335 14473
rect 11940 14436 11976 14464
rect 11882 14424 11888 14427
rect 11940 14424 11946 14436
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 15289 14467 15347 14473
rect 14323 14436 15240 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 15212 14408 15240 14436
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 16114 14464 16120 14476
rect 16075 14436 16120 14464
rect 15289 14427 15347 14433
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 17770 14464 17776 14476
rect 16816 14436 17776 14464
rect 16816 14424 16822 14436
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 18012 14436 18153 14464
rect 18012 14424 18018 14436
rect 18141 14433 18153 14436
rect 18187 14433 18199 14467
rect 18248 14464 18276 14504
rect 19518 14492 19524 14544
rect 19576 14532 19582 14544
rect 20162 14532 20168 14544
rect 19576 14504 20168 14532
rect 19576 14492 19582 14504
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 19061 14467 19119 14473
rect 18248 14436 18368 14464
rect 18141 14427 18199 14433
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 10704 14368 11621 14396
rect 11609 14365 11621 14368
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 12952 14368 13829 14396
rect 12952 14356 12958 14368
rect 13817 14365 13829 14368
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 15194 14356 15200 14408
rect 15252 14356 15258 14408
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14396 15623 14399
rect 15746 14396 15752 14408
rect 15611 14368 15752 14396
rect 15611 14365 15623 14368
rect 15565 14359 15623 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 18340 14405 18368 14436
rect 19061 14433 19073 14467
rect 19107 14464 19119 14467
rect 19150 14464 19156 14476
rect 19107 14436 19156 14464
rect 19107 14433 19119 14436
rect 19061 14427 19119 14433
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 19328 14467 19386 14473
rect 19328 14433 19340 14467
rect 19374 14464 19386 14467
rect 20346 14464 20352 14476
rect 19374 14436 20352 14464
rect 19374 14433 19386 14436
rect 19328 14427 19386 14433
rect 20346 14424 20352 14436
rect 20404 14424 20410 14476
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 17920 14368 18245 14396
rect 17920 14356 17926 14368
rect 18233 14365 18245 14368
rect 18279 14365 18291 14399
rect 18233 14359 18291 14365
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20220 14368 20913 14396
rect 20220 14356 20226 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 17402 14288 17408 14340
rect 17460 14328 17466 14340
rect 18506 14328 18512 14340
rect 17460 14300 18512 14328
rect 17460 14288 17466 14300
rect 18506 14288 18512 14300
rect 18564 14288 18570 14340
rect 8205 14263 8263 14269
rect 8205 14229 8217 14263
rect 8251 14260 8263 14263
rect 9858 14260 9864 14272
rect 8251 14232 9864 14260
rect 8251 14229 8263 14232
rect 8205 14223 8263 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 11054 14260 11060 14272
rect 11015 14232 11060 14260
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 13265 14263 13323 14269
rect 13265 14260 13277 14263
rect 13136 14232 13277 14260
rect 13136 14220 13142 14232
rect 13265 14229 13277 14232
rect 13311 14229 13323 14263
rect 17770 14260 17776 14272
rect 17731 14232 17776 14260
rect 13265 14223 13323 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 8478 14056 8484 14068
rect 8439 14028 8484 14056
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 11756 14028 12449 14056
rect 11756 14016 11762 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 12437 14019 12495 14025
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 13504 14028 13645 14056
rect 13504 14016 13510 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 14608 14028 14657 14056
rect 14608 14016 14614 14028
rect 14645 14025 14657 14028
rect 14691 14025 14703 14059
rect 15286 14056 15292 14068
rect 14645 14019 14703 14025
rect 14752 14028 15292 14056
rect 11333 13991 11391 13997
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 11790 13988 11796 14000
rect 11379 13960 11796 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 13096 13960 14320 13988
rect 8570 13880 8576 13932
rect 8628 13920 8634 13932
rect 9125 13923 9183 13929
rect 8628 13892 9076 13920
rect 8628 13880 8634 13892
rect 8938 13852 8944 13864
rect 8899 13824 8944 13852
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 9048 13852 9076 13892
rect 9125 13889 9137 13923
rect 9171 13920 9183 13923
rect 9858 13920 9864 13932
rect 9171 13892 9864 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 10870 13920 10876 13932
rect 10827 13892 10876 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 11882 13920 11888 13932
rect 11020 13892 11468 13920
rect 11843 13892 11888 13920
rect 11020 13880 11026 13892
rect 10597 13855 10655 13861
rect 9048 13824 10548 13852
rect 8849 13787 8907 13793
rect 8849 13753 8861 13787
rect 8895 13784 8907 13787
rect 9493 13787 9551 13793
rect 9493 13784 9505 13787
rect 8895 13756 9505 13784
rect 8895 13753 8907 13756
rect 8849 13747 8907 13753
rect 9493 13753 9505 13756
rect 9539 13753 9551 13787
rect 10520 13784 10548 13824
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 11330 13852 11336 13864
rect 10643 13824 11336 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 11440 13852 11468 13892
rect 11882 13880 11888 13892
rect 11940 13920 11946 13932
rect 13096 13929 13124 13960
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 11940 13892 13093 13920
rect 11940 13880 11946 13892
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13814 13880 13820 13932
rect 13872 13920 13878 13932
rect 14292 13929 14320 13960
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 13872 13892 14105 13920
rect 13872 13880 13878 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13920 14335 13923
rect 14752 13920 14780 14028
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 16114 14016 16120 14068
rect 16172 14056 16178 14068
rect 16574 14056 16580 14068
rect 16172 14028 16580 14056
rect 16172 14016 16178 14028
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17276 14028 17693 14056
rect 17276 14016 17282 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 17681 14019 17739 14025
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 18012 14028 18061 14056
rect 18012 14016 18018 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 19978 14056 19984 14068
rect 19843 14028 19984 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 20993 14059 21051 14065
rect 20993 14056 21005 14059
rect 20680 14028 21005 14056
rect 20680 14016 20686 14028
rect 20993 14025 21005 14028
rect 21039 14025 21051 14059
rect 20993 14019 21051 14025
rect 15654 13988 15660 14000
rect 15120 13960 15660 13988
rect 15120 13929 15148 13960
rect 15654 13948 15660 13960
rect 15712 13988 15718 14000
rect 16209 13991 16267 13997
rect 16209 13988 16221 13991
rect 15712 13960 16221 13988
rect 15712 13948 15718 13960
rect 16209 13957 16221 13960
rect 16255 13957 16267 13991
rect 16209 13951 16267 13957
rect 14323 13892 14780 13920
rect 15105 13923 15163 13929
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 15105 13889 15117 13923
rect 15151 13889 15163 13923
rect 15286 13920 15292 13932
rect 15247 13892 15292 13920
rect 15105 13883 15163 13889
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 18598 13920 18604 13932
rect 18559 13892 18604 13920
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 20346 13920 20352 13932
rect 20307 13892 20352 13920
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11440 13824 11805 13852
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12676 13824 12817 13852
rect 12676 13812 12682 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 15746 13852 15752 13864
rect 15707 13824 15752 13852
rect 12805 13815 12863 13821
rect 12820 13784 12848 13815
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 16298 13852 16304 13864
rect 16259 13824 16304 13852
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 16408 13824 18521 13852
rect 15013 13787 15071 13793
rect 10520 13756 11100 13784
rect 12820 13756 14596 13784
rect 9493 13747 9551 13753
rect 10134 13716 10140 13728
rect 10095 13688 10140 13716
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10686 13716 10692 13728
rect 10551 13688 10692 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 11072 13716 11100 13756
rect 11701 13719 11759 13725
rect 11701 13716 11713 13719
rect 11072 13688 11713 13716
rect 11701 13685 11713 13688
rect 11747 13716 11759 13719
rect 11790 13716 11796 13728
rect 11747 13688 11796 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 12434 13716 12440 13728
rect 12308 13688 12440 13716
rect 12308 13676 12314 13688
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 12894 13716 12900 13728
rect 12584 13688 12900 13716
rect 12584 13676 12590 13688
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 13998 13716 14004 13728
rect 13959 13688 14004 13716
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 14568 13716 14596 13756
rect 15013 13753 15025 13787
rect 15059 13784 15071 13787
rect 15654 13784 15660 13796
rect 15059 13756 15660 13784
rect 15059 13753 15071 13756
rect 15013 13747 15071 13753
rect 15654 13744 15660 13756
rect 15712 13744 15718 13796
rect 16408 13784 16436 13824
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 18509 13815 18567 13821
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18840 13824 19073 13852
rect 18840 13812 18846 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 20162 13852 20168 13864
rect 20123 13824 20168 13852
rect 19061 13815 19119 13821
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20806 13852 20812 13864
rect 20767 13824 20812 13852
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 15856 13756 16436 13784
rect 16568 13787 16626 13793
rect 15856 13716 15884 13756
rect 16568 13753 16580 13787
rect 16614 13784 16626 13787
rect 18598 13784 18604 13796
rect 16614 13756 18604 13784
rect 16614 13753 16626 13756
rect 16568 13747 16626 13753
rect 18598 13744 18604 13756
rect 18656 13744 18662 13796
rect 19334 13784 19340 13796
rect 19295 13756 19340 13784
rect 19334 13744 19340 13756
rect 19392 13744 19398 13796
rect 19794 13744 19800 13796
rect 19852 13784 19858 13796
rect 20070 13784 20076 13796
rect 19852 13756 20076 13784
rect 19852 13744 19858 13756
rect 20070 13744 20076 13756
rect 20128 13784 20134 13796
rect 20257 13787 20315 13793
rect 20257 13784 20269 13787
rect 20128 13756 20269 13784
rect 20128 13744 20134 13756
rect 20257 13753 20269 13756
rect 20303 13753 20315 13787
rect 20257 13747 20315 13753
rect 14568 13688 15884 13716
rect 15930 13676 15936 13728
rect 15988 13716 15994 13728
rect 16209 13719 16267 13725
rect 15988 13688 16033 13716
rect 15988 13676 15994 13688
rect 16209 13685 16221 13719
rect 16255 13716 16267 13719
rect 17678 13716 17684 13728
rect 16255 13688 17684 13716
rect 16255 13685 16267 13688
rect 16209 13679 16267 13685
rect 17678 13676 17684 13688
rect 17736 13716 17742 13728
rect 18417 13719 18475 13725
rect 18417 13716 18429 13719
rect 17736 13688 18429 13716
rect 17736 13676 17742 13688
rect 18417 13685 18429 13688
rect 18463 13685 18475 13719
rect 18417 13679 18475 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13512 9367 13515
rect 9674 13512 9680 13524
rect 9355 13484 9680 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 11330 13512 11336 13524
rect 11291 13484 11336 13512
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11701 13515 11759 13521
rect 11701 13481 11713 13515
rect 11747 13512 11759 13515
rect 12526 13512 12532 13524
rect 11747 13484 12532 13512
rect 11747 13481 11759 13484
rect 11701 13475 11759 13481
rect 10226 13404 10232 13456
rect 10284 13444 10290 13456
rect 11716 13444 11744 13475
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12710 13512 12716 13524
rect 12671 13484 12716 13512
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 13998 13512 14004 13524
rect 13959 13484 14004 13512
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 16114 13512 16120 13524
rect 14108 13484 16120 13512
rect 10284 13416 11744 13444
rect 11793 13447 11851 13453
rect 10284 13404 10290 13416
rect 11793 13413 11805 13447
rect 11839 13444 11851 13447
rect 12066 13444 12072 13456
rect 11839 13416 12072 13444
rect 11839 13413 11851 13416
rect 11793 13407 11851 13413
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 14108 13444 14136 13484
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13512 16359 13515
rect 16390 13512 16396 13524
rect 16347 13484 16396 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16666 13472 16672 13524
rect 16724 13512 16730 13524
rect 17129 13515 17187 13521
rect 17129 13512 17141 13515
rect 16724 13484 17141 13512
rect 16724 13472 16730 13484
rect 17129 13481 17141 13484
rect 17175 13481 17187 13515
rect 17129 13475 17187 13481
rect 17221 13515 17279 13521
rect 17221 13481 17233 13515
rect 17267 13512 17279 13515
rect 17770 13512 17776 13524
rect 17267 13484 17776 13512
rect 17267 13481 17279 13484
rect 17221 13475 17279 13481
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 18969 13515 19027 13521
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19058 13512 19064 13524
rect 19015 13484 19064 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 19797 13515 19855 13521
rect 19797 13481 19809 13515
rect 19843 13512 19855 13515
rect 19886 13512 19892 13524
rect 19843 13484 19892 13512
rect 19843 13481 19855 13484
rect 19797 13475 19855 13481
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 19334 13444 19340 13456
rect 12728 13416 14136 13444
rect 14660 13416 19340 13444
rect 12728 13388 12756 13416
rect 9490 13376 9496 13388
rect 9451 13348 9496 13376
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9674 13376 9680 13388
rect 9635 13348 9680 13376
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 9944 13379 10002 13385
rect 9944 13345 9956 13379
rect 9990 13376 10002 13379
rect 11054 13376 11060 13388
rect 9990 13348 11060 13376
rect 9990 13345 10002 13348
rect 9944 13339 10002 13345
rect 11054 13336 11060 13348
rect 11112 13376 11118 13388
rect 11112 13348 11928 13376
rect 11112 13336 11118 13348
rect 11900 13317 11928 13348
rect 12710 13336 12716 13388
rect 12768 13336 12774 13388
rect 12897 13379 12955 13385
rect 12897 13345 12909 13379
rect 12943 13345 12955 13379
rect 13078 13376 13084 13388
rect 13039 13348 13084 13376
rect 12897 13339 12955 13345
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 12912 13240 12940 13339
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 14660 13385 14688 13416
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 14645 13379 14703 13385
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 15470 13376 15476 13388
rect 14645 13339 14703 13345
rect 14844 13348 15476 13376
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13403 13280 14780 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 14274 13240 14280 13252
rect 12912 13212 14280 13240
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 10870 13132 10876 13184
rect 10928 13172 10934 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10928 13144 11069 13172
rect 10928 13132 10934 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 14642 13172 14648 13184
rect 12124 13144 14648 13172
rect 12124 13132 12130 13144
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 14752 13172 14780 13280
rect 14844 13249 14872 13348
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 18138 13376 18144 13388
rect 18099 13348 18144 13376
rect 18138 13336 18144 13348
rect 18196 13336 18202 13388
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 18785 13379 18843 13385
rect 18785 13376 18797 13379
rect 18564 13348 18797 13376
rect 18564 13336 18570 13348
rect 18785 13345 18797 13348
rect 18831 13345 18843 13379
rect 19702 13376 19708 13388
rect 19663 13348 19708 13376
rect 18785 13339 18843 13345
rect 19702 13336 19708 13348
rect 19760 13336 19766 13388
rect 15746 13308 15752 13320
rect 15707 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 15930 13308 15936 13320
rect 15891 13280 15936 13308
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13308 17463 13311
rect 17494 13308 17500 13320
rect 17451 13280 17500 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13308 18475 13311
rect 18598 13308 18604 13320
rect 18463 13280 18604 13308
rect 18463 13277 18475 13280
rect 18417 13271 18475 13277
rect 18598 13268 18604 13280
rect 18656 13308 18662 13320
rect 19058 13308 19064 13320
rect 18656 13280 19064 13308
rect 18656 13268 18662 13280
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19978 13308 19984 13320
rect 19939 13280 19984 13308
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 14829 13243 14887 13249
rect 14829 13209 14841 13243
rect 14875 13209 14887 13243
rect 14829 13203 14887 13209
rect 15194 13200 15200 13252
rect 15252 13240 15258 13252
rect 15289 13243 15347 13249
rect 15289 13240 15301 13243
rect 15252 13212 15301 13240
rect 15252 13200 15258 13212
rect 15289 13209 15301 13212
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 17773 13243 17831 13249
rect 17773 13209 17785 13243
rect 17819 13240 17831 13243
rect 17862 13240 17868 13252
rect 17819 13212 17868 13240
rect 17819 13209 17831 13212
rect 17773 13203 17831 13209
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 16574 13172 16580 13184
rect 14752 13144 16580 13172
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 16761 13175 16819 13181
rect 16761 13141 16773 13175
rect 16807 13172 16819 13175
rect 18782 13172 18788 13184
rect 16807 13144 18788 13172
rect 16807 13141 16819 13144
rect 16761 13135 16819 13141
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 19337 13175 19395 13181
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 20438 13172 20444 13184
rect 19383 13144 20444 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 10597 12971 10655 12977
rect 8996 12940 9904 12968
rect 8996 12928 9002 12940
rect 9876 12900 9904 12940
rect 10597 12937 10609 12971
rect 10643 12968 10655 12971
rect 11146 12968 11152 12980
rect 10643 12940 11152 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 12710 12968 12716 12980
rect 11256 12940 12716 12968
rect 11256 12900 11284 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16577 12971 16635 12977
rect 16577 12968 16589 12971
rect 15988 12940 16589 12968
rect 15988 12928 15994 12940
rect 16577 12937 16589 12940
rect 16623 12937 16635 12971
rect 16577 12931 16635 12937
rect 16853 12971 16911 12977
rect 16853 12937 16865 12971
rect 16899 12968 16911 12971
rect 17126 12968 17132 12980
rect 16899 12940 17132 12968
rect 16899 12937 16911 12940
rect 16853 12931 16911 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 18966 12968 18972 12980
rect 18616 12940 18972 12968
rect 9876 12872 11284 12900
rect 12437 12903 12495 12909
rect 12437 12869 12449 12903
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10192 12804 11069 12832
rect 10192 12792 10198 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12764 8999 12767
rect 9674 12764 9680 12776
rect 8987 12736 9680 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 11164 12764 11192 12795
rect 10336 12736 11192 12764
rect 11609 12767 11667 12773
rect 9208 12699 9266 12705
rect 9208 12665 9220 12699
rect 9254 12696 9266 12699
rect 10226 12696 10232 12708
rect 9254 12668 10232 12696
rect 9254 12665 9266 12668
rect 9208 12659 9266 12665
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 10336 12637 10364 12736
rect 11609 12733 11621 12767
rect 11655 12764 11667 12767
rect 12452 12764 12480 12863
rect 15194 12860 15200 12912
rect 15252 12860 15258 12912
rect 13078 12832 13084 12844
rect 13039 12804 13084 12832
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 15212 12832 15240 12860
rect 14700 12804 15240 12832
rect 17497 12835 17555 12841
rect 14700 12792 14706 12804
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 18325 12835 18383 12841
rect 17543 12804 18276 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 11655 12736 12480 12764
rect 11655 12733 11667 12736
rect 11609 12727 11667 12733
rect 12802 12724 12808 12776
rect 12860 12724 12866 12776
rect 12986 12724 12992 12776
rect 13044 12764 13050 12776
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 13044 12736 13553 12764
rect 13044 12724 13050 12736
rect 13541 12733 13553 12736
rect 13587 12764 13599 12767
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 13587 12736 15209 12764
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 15197 12733 15209 12736
rect 15243 12764 15255 12767
rect 16298 12764 16304 12776
rect 15243 12736 16304 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 18012 12736 18061 12764
rect 18012 12724 18018 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18248 12764 18276 12804
rect 18325 12801 18337 12835
rect 18371 12832 18383 12835
rect 18616 12832 18644 12940
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 19058 12928 19064 12980
rect 19116 12968 19122 12980
rect 20165 12971 20223 12977
rect 20165 12968 20177 12971
rect 19116 12940 20177 12968
rect 19116 12928 19122 12940
rect 20165 12937 20177 12940
rect 20211 12937 20223 12971
rect 20165 12931 20223 12937
rect 20714 12832 20720 12844
rect 18371 12804 18644 12832
rect 20675 12804 20720 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 18598 12764 18604 12776
rect 18248 12736 18604 12764
rect 18049 12727 18107 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12733 18843 12767
rect 20438 12764 20444 12776
rect 20399 12736 20444 12764
rect 18785 12727 18843 12733
rect 11885 12699 11943 12705
rect 11885 12665 11897 12699
rect 11931 12696 11943 12699
rect 12820 12696 12848 12724
rect 13814 12705 13820 12708
rect 13808 12696 13820 12705
rect 11931 12668 12848 12696
rect 13775 12668 13820 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 13808 12659 13820 12668
rect 13814 12656 13820 12659
rect 13872 12656 13878 12708
rect 15464 12699 15522 12705
rect 15464 12696 15476 12699
rect 14936 12668 15476 12696
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9640 12600 10333 12628
rect 9640 12588 9646 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10962 12628 10968 12640
rect 10923 12600 10968 12628
rect 10321 12591 10379 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12492 12600 12817 12628
rect 12492 12588 12498 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 12805 12591 12863 12597
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 12952 12600 12997 12628
rect 12952 12588 12958 12600
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14366 12628 14372 12640
rect 13964 12600 14372 12628
rect 13964 12588 13970 12600
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 14936 12637 14964 12668
rect 15464 12665 15476 12668
rect 15510 12696 15522 12699
rect 16022 12696 16028 12708
rect 15510 12668 16028 12696
rect 15510 12665 15522 12668
rect 15464 12659 15522 12665
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 17218 12696 17224 12708
rect 17179 12668 17224 12696
rect 17218 12656 17224 12668
rect 17276 12656 17282 12708
rect 14921 12631 14979 12637
rect 14921 12597 14933 12631
rect 14967 12597 14979 12631
rect 14921 12591 14979 12597
rect 15838 12588 15844 12640
rect 15896 12628 15902 12640
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 15896 12600 17325 12628
rect 15896 12588 15902 12600
rect 17313 12597 17325 12600
rect 17359 12628 17371 12631
rect 17402 12628 17408 12640
rect 17359 12600 17408 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 18800 12628 18828 12727
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 19052 12699 19110 12705
rect 19052 12665 19064 12699
rect 19098 12696 19110 12699
rect 19978 12696 19984 12708
rect 19098 12668 19984 12696
rect 19098 12665 19110 12668
rect 19052 12659 19110 12665
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 19150 12628 19156 12640
rect 18656 12600 19156 12628
rect 18656 12588 18662 12600
rect 19150 12588 19156 12600
rect 19208 12628 19214 12640
rect 19334 12628 19340 12640
rect 19208 12600 19340 12628
rect 19208 12588 19214 12600
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 10870 12424 10876 12436
rect 10284 12396 10876 12424
rect 10284 12384 10290 12396
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12393 12863 12427
rect 12805 12387 12863 12393
rect 8012 12359 8070 12365
rect 8012 12325 8024 12359
rect 8058 12356 8070 12359
rect 9582 12356 9588 12368
rect 8058 12328 9588 12356
rect 8058 12325 8070 12328
rect 8012 12319 8070 12325
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 12820 12356 12848 12387
rect 13078 12384 13084 12436
rect 13136 12384 13142 12436
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 19702 12424 19708 12436
rect 17635 12396 19708 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 13096 12356 13124 12384
rect 13326 12359 13384 12365
rect 13326 12356 13338 12359
rect 12820 12328 13338 12356
rect 13326 12325 13338 12328
rect 13372 12325 13384 12359
rect 13326 12319 13384 12325
rect 15930 12316 15936 12368
rect 15988 12356 15994 12368
rect 16178 12359 16236 12365
rect 16178 12356 16190 12359
rect 15988 12328 16190 12356
rect 15988 12316 15994 12328
rect 16178 12325 16190 12328
rect 16224 12325 16236 12359
rect 16178 12319 16236 12325
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 16850 12356 16856 12368
rect 16448 12328 16856 12356
rect 16448 12316 16454 12328
rect 16850 12316 16856 12328
rect 16908 12316 16914 12368
rect 17957 12359 18015 12365
rect 17957 12325 17969 12359
rect 18003 12356 18015 12359
rect 20901 12359 20959 12365
rect 20901 12356 20913 12359
rect 18003 12328 20913 12356
rect 18003 12325 18015 12328
rect 17957 12319 18015 12325
rect 20901 12325 20913 12328
rect 20947 12325 20959 12359
rect 20901 12319 20959 12325
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12288 7803 12291
rect 9674 12288 9680 12300
rect 7791 12260 9680 12288
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 10652 12260 10701 12288
rect 10652 12248 10658 12260
rect 10689 12257 10701 12260
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11054 12288 11060 12300
rect 10827 12260 11060 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11692 12291 11750 12297
rect 11692 12257 11704 12291
rect 11738 12288 11750 12291
rect 12066 12288 12072 12300
rect 11738 12260 12072 12288
rect 11738 12257 11750 12260
rect 11692 12251 11750 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 13044 12260 13093 12288
rect 13044 12248 13050 12260
rect 13081 12257 13093 12260
rect 13127 12257 13139 12291
rect 13081 12251 13139 12257
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 17862 12288 17868 12300
rect 14608 12260 17868 12288
rect 14608 12248 14614 12260
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 18874 12297 18880 12300
rect 18868 12288 18880 12297
rect 18248 12260 18880 12288
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 11425 12223 11483 12229
rect 10928 12192 10973 12220
rect 10928 12180 10934 12192
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15470 12220 15476 12232
rect 15335 12192 15476 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 10321 12155 10379 12161
rect 10321 12121 10333 12155
rect 10367 12152 10379 12155
rect 10962 12152 10968 12164
rect 10367 12124 10968 12152
rect 10367 12121 10379 12124
rect 10321 12115 10379 12121
rect 10962 12112 10968 12124
rect 11020 12112 11026 12164
rect 9122 12084 9128 12096
rect 9083 12056 9128 12084
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10870 12084 10876 12096
rect 9732 12056 10876 12084
rect 9732 12044 9738 12056
rect 10870 12044 10876 12056
rect 10928 12084 10934 12096
rect 11440 12084 11468 12183
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 14366 12112 14372 12164
rect 14424 12152 14430 12164
rect 14424 12124 15148 12152
rect 14424 12112 14430 12124
rect 10928 12056 11468 12084
rect 14461 12087 14519 12093
rect 10928 12044 10934 12056
rect 14461 12053 14473 12087
rect 14507 12084 14519 12087
rect 14642 12084 14648 12096
rect 14507 12056 14648 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 15120 12084 15148 12124
rect 15194 12084 15200 12096
rect 15120 12056 15200 12084
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 15948 12084 15976 12183
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 18248 12229 18276 12260
rect 18868 12251 18880 12260
rect 18874 12248 18880 12251
rect 18932 12248 18938 12300
rect 19150 12248 19156 12300
rect 19208 12288 19214 12300
rect 20257 12291 20315 12297
rect 20257 12288 20269 12291
rect 19208 12260 20269 12288
rect 19208 12248 19214 12260
rect 20257 12257 20269 12260
rect 20303 12257 20315 12291
rect 20257 12251 20315 12257
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 17460 12192 18061 12220
rect 17460 12180 17466 12192
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12189 18291 12223
rect 18598 12220 18604 12232
rect 18559 12192 18604 12220
rect 18233 12183 18291 12189
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 16298 12084 16304 12096
rect 15948 12056 16304 12084
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 17310 12084 17316 12096
rect 17271 12056 17316 12084
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 19300 12056 20453 12084
rect 19300 12044 19306 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 12434 11880 12440 11892
rect 11563 11852 12440 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12529 11883 12587 11889
rect 12529 11849 12541 11883
rect 12575 11880 12587 11883
rect 12894 11880 12900 11892
rect 12575 11852 12900 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 12995 11852 13584 11880
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 12995 11812 13023 11852
rect 10744 11784 13023 11812
rect 13449 11815 13507 11821
rect 10744 11772 10750 11784
rect 13449 11781 13461 11815
rect 13495 11781 13507 11815
rect 13556 11812 13584 11852
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13998 11880 14004 11892
rect 13780 11852 14004 11880
rect 13780 11840 13786 11852
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 15473 11883 15531 11889
rect 15473 11849 15485 11883
rect 15519 11880 15531 11883
rect 15746 11880 15752 11892
rect 15519 11852 15752 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 16485 11883 16543 11889
rect 16485 11880 16497 11883
rect 16356 11852 16497 11880
rect 16356 11840 16362 11852
rect 16485 11849 16497 11852
rect 16531 11880 16543 11883
rect 18598 11880 18604 11892
rect 16531 11852 18604 11880
rect 16531 11849 16543 11852
rect 16485 11843 16543 11849
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19337 11883 19395 11889
rect 19337 11849 19349 11883
rect 19383 11880 19395 11883
rect 19426 11880 19432 11892
rect 19383 11852 19432 11880
rect 19383 11849 19395 11852
rect 19337 11843 19395 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 19536 11852 21097 11880
rect 17586 11812 17592 11824
rect 13556 11784 17592 11812
rect 13449 11775 13507 11781
rect 10594 11744 10600 11756
rect 10555 11716 10600 11744
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 12066 11744 12072 11756
rect 12027 11716 12072 11744
rect 12066 11704 12072 11716
rect 12124 11744 12130 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 12124 11716 13093 11744
rect 12124 11704 12130 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 9398 11676 9404 11688
rect 9359 11648 9404 11676
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11676 11299 11679
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11287 11648 11897 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 13464 11676 13492 11775
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 18874 11772 18880 11824
rect 18932 11812 18938 11824
rect 19536 11812 19564 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 21085 11843 21143 11849
rect 18932 11784 19564 11812
rect 18932 11772 18938 11784
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13872 11716 14105 11744
rect 13872 11704 13878 11716
rect 14093 11713 14105 11716
rect 14139 11744 14151 11747
rect 14642 11744 14648 11756
rect 14139 11716 14648 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14642 11704 14648 11716
rect 14700 11744 14706 11756
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14700 11716 14933 11744
rect 14700 11704 14706 11716
rect 14921 11713 14933 11716
rect 14967 11744 14979 11747
rect 15838 11744 15844 11756
rect 14967 11716 15844 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16022 11744 16028 11756
rect 15983 11716 16028 11744
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 16632 11716 16804 11744
rect 16632 11704 16638 11716
rect 15933 11679 15991 11685
rect 15933 11676 15945 11679
rect 13464 11648 15945 11676
rect 11885 11639 11943 11645
rect 15933 11645 15945 11648
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16540 11648 16681 11676
rect 16540 11636 16546 11648
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16776 11676 16804 11716
rect 17310 11704 17316 11756
rect 17368 11744 17374 11756
rect 17497 11747 17555 11753
rect 17497 11744 17509 11747
rect 17368 11716 17509 11744
rect 17368 11704 17374 11716
rect 17497 11713 17509 11716
rect 17543 11744 17555 11747
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17543 11716 18613 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 19705 11747 19763 11753
rect 19705 11744 19717 11747
rect 19392 11716 19717 11744
rect 19392 11704 19398 11716
rect 19705 11713 19717 11716
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 16776 11648 19165 11676
rect 16669 11639 16727 11645
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 19153 11639 19211 11645
rect 9677 11611 9735 11617
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 13998 11608 14004 11620
rect 9723 11580 14004 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 15841 11611 15899 11617
rect 15841 11608 15853 11611
rect 14292 11580 15853 11608
rect 8941 11543 8999 11549
rect 8941 11509 8953 11543
rect 8987 11540 8999 11543
rect 10042 11540 10048 11552
rect 8987 11512 10048 11540
rect 8987 11509 8999 11512
rect 8941 11503 8999 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 11977 11543 12035 11549
rect 11977 11509 11989 11543
rect 12023 11540 12035 11543
rect 12434 11540 12440 11552
rect 12023 11512 12440 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13044 11512 13089 11540
rect 13044 11500 13050 11512
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13688 11512 13829 11540
rect 13688 11500 13694 11512
rect 13817 11509 13829 11512
rect 13863 11509 13875 11543
rect 13817 11503 13875 11509
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 14292 11549 14320 11580
rect 15841 11577 15853 11580
rect 15887 11577 15899 11611
rect 15841 11571 15899 11577
rect 16114 11568 16120 11620
rect 16172 11608 16178 11620
rect 17221 11611 17279 11617
rect 17221 11608 17233 11611
rect 16172 11580 17233 11608
rect 16172 11568 16178 11580
rect 17221 11577 17233 11580
rect 17267 11577 17279 11611
rect 17221 11571 17279 11577
rect 17313 11611 17371 11617
rect 17313 11577 17325 11611
rect 17359 11608 17371 11611
rect 17494 11608 17500 11620
rect 17359 11580 17500 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 14277 11543 14335 11549
rect 13964 11512 14009 11540
rect 13964 11500 13970 11512
rect 14277 11509 14289 11543
rect 14323 11509 14335 11543
rect 14277 11503 14335 11509
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 14608 11512 14657 11540
rect 14608 11500 14614 11512
rect 14645 11509 14657 11512
rect 14691 11509 14703 11543
rect 14645 11503 14703 11509
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15930 11540 15936 11552
rect 14783 11512 15936 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16850 11540 16856 11552
rect 16811 11512 16856 11540
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17328 11540 17356 11571
rect 17494 11568 17500 11580
rect 17552 11568 17558 11620
rect 18417 11611 18475 11617
rect 18417 11577 18429 11611
rect 18463 11608 18475 11611
rect 18598 11608 18604 11620
rect 18463 11580 18604 11608
rect 18463 11577 18475 11580
rect 18417 11571 18475 11577
rect 18598 11568 18604 11580
rect 18656 11568 18662 11620
rect 19972 11611 20030 11617
rect 19972 11577 19984 11611
rect 20018 11608 20030 11611
rect 20070 11608 20076 11620
rect 20018 11580 20076 11608
rect 20018 11577 20030 11580
rect 19972 11571 20030 11577
rect 20070 11568 20076 11580
rect 20128 11568 20134 11620
rect 17184 11512 17356 11540
rect 17184 11500 17190 11512
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17828 11512 18061 11540
rect 17828 11500 17834 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11540 18567 11543
rect 19058 11540 19064 11552
rect 18555 11512 19064 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 19058 11500 19064 11512
rect 19116 11500 19122 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9456 11308 9689 11336
rect 9456 11296 9462 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 9677 11299 9735 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 12124 11308 12265 11336
rect 12124 11296 12130 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 14274 11336 14280 11348
rect 14235 11308 14280 11336
rect 12253 11299 12311 11305
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 15746 11336 15752 11348
rect 15703 11308 15752 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 17034 11336 17040 11348
rect 16040 11308 17040 11336
rect 8196 11271 8254 11277
rect 8196 11237 8208 11271
rect 8242 11268 8254 11271
rect 9122 11268 9128 11280
rect 8242 11240 9128 11268
rect 8242 11237 8254 11240
rect 8196 11231 8254 11237
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 10686 11268 10692 11280
rect 10560 11240 10692 11268
rect 10560 11228 10566 11240
rect 10686 11228 10692 11240
rect 10744 11268 10750 11280
rect 13906 11268 13912 11280
rect 10744 11240 13912 11268
rect 10744 11228 10750 11240
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11200 7987 11203
rect 10870 11200 10876 11212
rect 7975 11172 10876 11200
rect 7975 11169 7987 11172
rect 7929 11163 7987 11169
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 11140 11203 11198 11209
rect 11140 11169 11152 11203
rect 11186 11200 11198 11203
rect 11882 11200 11888 11212
rect 11186 11172 11888 11200
rect 11186 11169 11198 11172
rect 11140 11163 11198 11169
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12342 11200 12348 11212
rect 12124 11172 12348 11200
rect 12124 11160 12130 11172
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 16040 11200 16068 11308
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17586 11296 17592 11348
rect 17644 11336 17650 11348
rect 20073 11339 20131 11345
rect 20073 11336 20085 11339
rect 17644 11308 20085 11336
rect 17644 11296 17650 11308
rect 20073 11305 20085 11308
rect 20119 11305 20131 11339
rect 20073 11299 20131 11305
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 16393 11271 16451 11277
rect 16393 11268 16405 11271
rect 16264 11240 16405 11268
rect 16264 11228 16270 11240
rect 16393 11237 16405 11240
rect 16439 11237 16451 11271
rect 16393 11231 16451 11237
rect 16936 11271 16994 11277
rect 16936 11237 16948 11271
rect 16982 11268 16994 11271
rect 17310 11268 17316 11280
rect 16982 11240 17316 11268
rect 16982 11237 16994 11240
rect 16936 11231 16994 11237
rect 17310 11228 17316 11240
rect 17368 11228 17374 11280
rect 18785 11271 18843 11277
rect 18785 11237 18797 11271
rect 18831 11268 18843 11271
rect 19794 11268 19800 11280
rect 18831 11240 19800 11268
rect 18831 11237 18843 11240
rect 18785 11231 18843 11237
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 13035 11172 16068 11200
rect 16117 11203 16175 11209
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 16758 11200 16764 11212
rect 16163 11172 16764 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16758 11160 16764 11172
rect 16816 11160 16822 11212
rect 18690 11200 18696 11212
rect 18651 11172 18696 11200
rect 18690 11160 18696 11172
rect 18748 11160 18754 11212
rect 19978 11200 19984 11212
rect 19939 11172 19984 11200
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9732 11104 10149 11132
rect 9732 11092 9738 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 9306 11064 9312 11076
rect 9267 11036 9312 11064
rect 9306 11024 9312 11036
rect 9364 11064 9370 11076
rect 10244 11064 10272 11095
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 15378 11132 15384 11144
rect 13412 11104 15384 11132
rect 13412 11092 13418 11104
rect 15378 11092 15384 11104
rect 15436 11132 15442 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15436 11104 15761 11132
rect 15436 11092 15442 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16669 11135 16727 11141
rect 15896 11104 15941 11132
rect 15896 11092 15902 11104
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 20165 11135 20223 11141
rect 20165 11101 20177 11135
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 9364 11036 10272 11064
rect 9364 11024 9370 11036
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 16114 11064 16120 11076
rect 13688 11036 16120 11064
rect 13688 11024 13694 11036
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 12986 10996 12992 11008
rect 11204 10968 12992 10996
rect 11204 10956 11210 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 15286 10996 15292 11008
rect 15247 10968 15292 10996
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 16684 10996 16712 11095
rect 17678 11024 17684 11076
rect 17736 11064 17742 11076
rect 18325 11067 18383 11073
rect 18325 11064 18337 11067
rect 17736 11036 18337 11064
rect 17736 11024 17742 11036
rect 18325 11033 18337 11036
rect 18371 11033 18383 11067
rect 18892 11064 18920 11095
rect 18325 11027 18383 11033
rect 18432 11036 18920 11064
rect 17034 10996 17040 11008
rect 16684 10968 17040 10996
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 17586 10956 17592 11008
rect 17644 10996 17650 11008
rect 18049 10999 18107 11005
rect 18049 10996 18061 10999
rect 17644 10968 18061 10996
rect 17644 10956 17650 10968
rect 18049 10965 18061 10968
rect 18095 10996 18107 10999
rect 18432 10996 18460 11036
rect 19242 11024 19248 11076
rect 19300 11064 19306 11076
rect 20180 11064 20208 11095
rect 19300 11036 20208 11064
rect 19300 11024 19306 11036
rect 18095 10968 18460 10996
rect 18095 10965 18107 10968
rect 18049 10959 18107 10965
rect 18506 10956 18512 11008
rect 18564 10996 18570 11008
rect 19613 10999 19671 11005
rect 19613 10996 19625 10999
rect 18564 10968 19625 10996
rect 18564 10956 18570 10968
rect 19613 10965 19625 10968
rect 19659 10965 19671 10999
rect 19613 10959 19671 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 8757 10795 8815 10801
rect 8757 10761 8769 10795
rect 8803 10792 8815 10795
rect 9674 10792 9680 10804
rect 8803 10764 9680 10792
rect 8803 10761 8815 10764
rect 8757 10755 8815 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 10060 10764 11468 10792
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 10060 10665 10088 10764
rect 11146 10684 11152 10736
rect 11204 10724 11210 10736
rect 11333 10727 11391 10733
rect 11333 10724 11345 10727
rect 11204 10696 11345 10724
rect 11204 10684 11210 10696
rect 11333 10693 11345 10696
rect 11379 10693 11391 10727
rect 11440 10724 11468 10764
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 12342 10792 12348 10804
rect 11664 10764 12348 10792
rect 11664 10752 11670 10764
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12492 10764 12537 10792
rect 12492 10752 12498 10764
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 12952 10764 13461 10792
rect 12952 10752 12958 10764
rect 13449 10761 13461 10764
rect 13495 10761 13507 10795
rect 13449 10755 13507 10761
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15654 10792 15660 10804
rect 15427 10764 15660 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 19150 10792 19156 10804
rect 16316 10764 19156 10792
rect 16316 10724 16344 10764
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 11440 10696 16344 10724
rect 11333 10687 11391 10693
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 9180 10628 9321 10656
rect 9180 10616 9186 10628
rect 9309 10625 9321 10628
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10625 10103 10659
rect 11882 10656 11888 10668
rect 11843 10628 11888 10656
rect 10045 10619 10103 10625
rect 11882 10616 11888 10628
rect 11940 10656 11946 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 11940 10628 13093 10656
rect 11940 10616 11946 10628
rect 13081 10625 13093 10628
rect 13127 10656 13139 10659
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13127 10628 14013 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 15102 10656 15108 10668
rect 15063 10628 15108 10656
rect 14001 10619 14059 10625
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15286 10616 15292 10668
rect 15344 10656 15350 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15344 10628 15853 10656
rect 15344 10616 15350 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 16022 10656 16028 10668
rect 15983 10628 16028 10656
rect 15841 10619 15899 10625
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18690 10656 18696 10668
rect 18095 10628 18696 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 19242 10656 19248 10668
rect 19203 10628 19248 10656
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 9766 10588 9772 10600
rect 9727 10560 9772 10588
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12584 10560 12817 10588
rect 12584 10548 12590 10560
rect 12805 10557 12817 10560
rect 12851 10588 12863 10591
rect 13170 10588 13176 10600
rect 12851 10560 13176 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 14366 10588 14372 10600
rect 13863 10560 14372 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14608 10560 15025 10588
rect 14608 10548 14614 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15470 10548 15476 10600
rect 15528 10588 15534 10600
rect 15749 10591 15807 10597
rect 15749 10588 15761 10591
rect 15528 10560 15761 10588
rect 15528 10548 15534 10560
rect 15749 10557 15761 10560
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 17034 10588 17040 10600
rect 16347 10560 17040 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 19061 10591 19119 10597
rect 19061 10588 19073 10591
rect 17920 10560 19073 10588
rect 17920 10548 17926 10560
rect 19061 10557 19073 10560
rect 19107 10557 19119 10591
rect 19061 10551 19119 10557
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 19392 10560 19625 10588
rect 19392 10548 19398 10560
rect 19613 10557 19625 10560
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 11793 10523 11851 10529
rect 11793 10520 11805 10523
rect 10744 10492 11805 10520
rect 10744 10480 10750 10492
rect 11793 10489 11805 10492
rect 11839 10489 11851 10523
rect 11793 10483 11851 10489
rect 14921 10523 14979 10529
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 15286 10520 15292 10532
rect 14967 10492 15292 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 16568 10523 16626 10529
rect 16568 10489 16580 10523
rect 16614 10520 16626 10523
rect 17494 10520 17500 10532
rect 16614 10492 17500 10520
rect 16614 10489 16626 10492
rect 16568 10483 16626 10489
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 18782 10480 18788 10532
rect 18840 10520 18846 10532
rect 19858 10523 19916 10529
rect 19858 10520 19870 10523
rect 18840 10492 19870 10520
rect 18840 10480 18846 10492
rect 19858 10489 19870 10492
rect 19904 10520 19916 10523
rect 20530 10520 20536 10532
rect 19904 10492 20536 10520
rect 19904 10489 19916 10492
rect 19858 10483 19916 10489
rect 20530 10480 20536 10492
rect 20588 10480 20594 10532
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 11606 10452 11612 10464
rect 9272 10424 11612 10452
rect 9272 10412 9278 10424
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10452 11759 10455
rect 12434 10452 12440 10464
rect 11747 10424 12440 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 12894 10452 12900 10464
rect 12855 10424 12900 10452
rect 12894 10412 12900 10424
rect 12952 10452 12958 10464
rect 13722 10452 13728 10464
rect 12952 10424 13728 10452
rect 12952 10412 12958 10424
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 13906 10452 13912 10464
rect 13867 10424 13912 10452
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 13998 10412 14004 10464
rect 14056 10452 14062 10464
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 14056 10424 14565 10452
rect 14056 10412 14062 10424
rect 14553 10421 14565 10424
rect 14599 10421 14611 10455
rect 14553 10415 14611 10421
rect 17586 10412 17592 10464
rect 17644 10452 17650 10464
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 17644 10424 17693 10452
rect 17644 10412 17650 10424
rect 17681 10421 17693 10424
rect 17727 10421 17739 10455
rect 18598 10452 18604 10464
rect 18559 10424 18604 10452
rect 17681 10415 17739 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 18966 10452 18972 10464
rect 18927 10424 18972 10452
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 20070 10452 20076 10464
rect 19116 10424 20076 10452
rect 19116 10412 19122 10424
rect 20070 10412 20076 10424
rect 20128 10452 20134 10464
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 20128 10424 21005 10452
rect 20128 10412 20134 10424
rect 20993 10421 21005 10424
rect 21039 10421 21051 10455
rect 20993 10415 21051 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 9088 10220 11836 10248
rect 9088 10208 9094 10220
rect 8196 10183 8254 10189
rect 8196 10149 8208 10183
rect 8242 10180 8254 10183
rect 9306 10180 9312 10192
rect 8242 10152 9312 10180
rect 8242 10149 8254 10152
rect 8196 10143 8254 10149
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 11698 10180 11704 10192
rect 10520 10152 11704 10180
rect 10520 10121 10548 10152
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10864 10115 10922 10121
rect 10864 10081 10876 10115
rect 10910 10112 10922 10115
rect 11146 10112 11152 10124
rect 10910 10084 11152 10112
rect 10910 10081 10922 10084
rect 10864 10075 10922 10081
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 7926 10044 7932 10056
rect 7887 10016 7932 10044
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10594 10044 10600 10056
rect 10336 10016 10600 10044
rect 10336 9985 10364 10016
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10321 9979 10379 9985
rect 10321 9945 10333 9979
rect 10367 9945 10379 9979
rect 11808 9976 11836 10220
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11940 10220 11989 10248
rect 11940 10208 11946 10220
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13446 10248 13452 10260
rect 12492 10220 13452 10248
rect 12492 10208 12498 10220
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 14185 10251 14243 10257
rect 14185 10248 14197 10251
rect 13679 10220 14197 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 14185 10217 14197 10220
rect 14231 10217 14243 10251
rect 14185 10211 14243 10217
rect 14550 10208 14556 10260
rect 14608 10248 14614 10260
rect 15010 10248 15016 10260
rect 14608 10220 15016 10248
rect 14608 10208 14614 10220
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 15102 10208 15108 10260
rect 15160 10248 15166 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 15160 10220 16681 10248
rect 15160 10208 15166 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 16945 10251 17003 10257
rect 16945 10248 16957 10251
rect 16816 10220 16957 10248
rect 16816 10208 16822 10220
rect 16945 10217 16957 10220
rect 16991 10217 17003 10251
rect 16945 10211 17003 10217
rect 17313 10251 17371 10257
rect 17313 10217 17325 10251
rect 17359 10248 17371 10251
rect 17678 10248 17684 10260
rect 17359 10220 17684 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 18012 10220 18153 10248
rect 18012 10208 18018 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18141 10211 18199 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 20530 10248 20536 10260
rect 20491 10220 20536 10248
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 13541 10183 13599 10189
rect 13541 10149 13553 10183
rect 13587 10180 13599 10183
rect 13998 10180 14004 10192
rect 13587 10152 14004 10180
rect 13587 10149 13599 10152
rect 13541 10143 13599 10149
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 14645 10183 14703 10189
rect 14645 10180 14657 10183
rect 14200 10152 14657 10180
rect 14200 10112 14228 10152
rect 14645 10149 14657 10152
rect 14691 10149 14703 10183
rect 14645 10143 14703 10149
rect 17402 10140 17408 10192
rect 17460 10180 17466 10192
rect 18506 10180 18512 10192
rect 17460 10152 17724 10180
rect 18467 10152 18512 10180
rect 17460 10140 17466 10152
rect 17696 10124 17724 10152
rect 18506 10140 18512 10152
rect 18564 10140 18570 10192
rect 19334 10180 19340 10192
rect 19168 10152 19340 10180
rect 14016 10084 14228 10112
rect 14553 10115 14611 10121
rect 14016 10056 14044 10084
rect 14553 10081 14565 10115
rect 14599 10112 14611 10115
rect 15378 10112 15384 10124
rect 14599 10084 15384 10112
rect 14599 10081 14611 10084
rect 14553 10075 14611 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15562 10121 15568 10124
rect 15556 10112 15568 10121
rect 15523 10084 15568 10112
rect 15556 10075 15568 10084
rect 15562 10072 15568 10075
rect 15620 10072 15626 10124
rect 17678 10072 17684 10124
rect 17736 10072 17742 10124
rect 19168 10121 19196 10152
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 19153 10115 19211 10121
rect 19153 10081 19165 10115
rect 19199 10081 19211 10115
rect 19153 10075 19211 10081
rect 19242 10072 19248 10124
rect 19300 10112 19306 10124
rect 19420 10115 19478 10121
rect 19420 10112 19432 10115
rect 19300 10084 19432 10112
rect 19300 10072 19306 10084
rect 19420 10081 19432 10084
rect 19466 10112 19478 10115
rect 19702 10112 19708 10124
rect 19466 10084 19708 10112
rect 19466 10081 19478 10084
rect 19420 10075 19478 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 13722 10044 13728 10056
rect 13683 10016 13728 10044
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 13998 10004 14004 10056
rect 14056 10004 14062 10056
rect 14734 10044 14740 10056
rect 14695 10016 14740 10044
rect 14734 10004 14740 10016
rect 14792 10044 14798 10056
rect 15102 10044 15108 10056
rect 14792 10016 15108 10044
rect 14792 10004 14798 10016
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 15252 10016 15301 10044
rect 15252 10004 15258 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 17402 10044 17408 10056
rect 17363 10016 17408 10044
rect 15289 10007 15347 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 17586 10044 17592 10056
rect 17547 10016 17592 10044
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 18782 10044 18788 10056
rect 18743 10016 18788 10044
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 11808 9948 13400 9976
rect 10321 9939 10379 9945
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 12618 9868 12624 9920
rect 12676 9908 12682 9920
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 12676 9880 13185 9908
rect 12676 9868 12682 9880
rect 13173 9877 13185 9880
rect 13219 9877 13231 9911
rect 13372 9908 13400 9948
rect 14366 9936 14372 9988
rect 14424 9976 14430 9988
rect 15010 9976 15016 9988
rect 14424 9948 15016 9976
rect 14424 9936 14430 9948
rect 15010 9936 15016 9948
rect 15068 9936 15074 9988
rect 18966 9908 18972 9920
rect 13372 9880 18972 9908
rect 13173 9871 13231 9877
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 14553 9707 14611 9713
rect 14553 9704 14565 9707
rect 14056 9676 14565 9704
rect 14056 9664 14062 9676
rect 14553 9673 14565 9676
rect 14599 9673 14611 9707
rect 14553 9667 14611 9673
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15565 9707 15623 9713
rect 15565 9704 15577 9707
rect 15436 9676 15577 9704
rect 15436 9664 15442 9676
rect 15565 9673 15577 9676
rect 15611 9673 15623 9707
rect 15565 9667 15623 9673
rect 16945 9707 17003 9713
rect 16945 9673 16957 9707
rect 16991 9704 17003 9707
rect 17402 9704 17408 9716
rect 16991 9676 17408 9704
rect 16991 9673 17003 9676
rect 16945 9667 17003 9673
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 11146 9596 11152 9648
rect 11204 9636 11210 9648
rect 11333 9639 11391 9645
rect 11333 9636 11345 9639
rect 11204 9608 11345 9636
rect 11204 9596 11210 9608
rect 11333 9605 11345 9608
rect 11379 9605 11391 9639
rect 11333 9599 11391 9605
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 11974 9568 11980 9580
rect 11931 9540 11980 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 15010 9568 15016 9580
rect 14240 9540 15016 9568
rect 14240 9528 14246 9540
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9568 15255 9571
rect 15562 9568 15568 9580
rect 15243 9540 15568 9568
rect 15243 9537 15255 9540
rect 15197 9531 15255 9537
rect 15562 9528 15568 9540
rect 15620 9568 15626 9580
rect 16206 9568 16212 9580
rect 15620 9540 16212 9568
rect 15620 9528 15626 9540
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 17494 9568 17500 9580
rect 17455 9540 17500 9568
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 7984 9472 8217 9500
rect 7984 9460 7990 9472
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 8472 9503 8530 9509
rect 8472 9469 8484 9503
rect 8518 9500 8530 9503
rect 8846 9500 8852 9512
rect 8518 9472 8852 9500
rect 8518 9469 8530 9472
rect 8472 9463 8530 9469
rect 8220 9432 8248 9463
rect 8846 9460 8852 9472
rect 8904 9500 8910 9512
rect 9306 9500 9312 9512
rect 8904 9472 9312 9500
rect 8904 9460 8910 9472
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9692 9472 9965 9500
rect 9692 9432 9720 9472
rect 9953 9469 9965 9472
rect 9999 9500 10011 9503
rect 10594 9500 10600 9512
rect 9999 9472 10600 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10594 9460 10600 9472
rect 10652 9500 10658 9512
rect 10652 9472 11100 9500
rect 10652 9460 10658 9472
rect 9858 9432 9864 9444
rect 8220 9404 9864 9432
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 10220 9435 10278 9441
rect 10220 9401 10232 9435
rect 10266 9432 10278 9435
rect 10962 9432 10968 9444
rect 10266 9404 10968 9432
rect 10266 9401 10278 9404
rect 10220 9395 10278 9401
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 11072 9432 11100 9472
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11480 9472 11621 9500
rect 11480 9460 11486 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12986 9500 12992 9512
rect 12483 9472 12992 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12452 9432 12480 9463
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 14274 9500 14280 9512
rect 14235 9472 14280 9500
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14642 9500 14648 9512
rect 14424 9472 14648 9500
rect 14424 9460 14430 9472
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9500 14979 9503
rect 16390 9500 16396 9512
rect 14967 9472 16396 9500
rect 14967 9469 14979 9472
rect 14921 9463 14979 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 16908 9472 17325 9500
rect 16908 9460 16914 9472
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 17405 9503 17463 9509
rect 17405 9469 17417 9503
rect 17451 9500 17463 9503
rect 17770 9500 17776 9512
rect 17451 9472 17776 9500
rect 17451 9469 17463 9472
rect 17405 9463 17463 9469
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 18046 9500 18052 9512
rect 17959 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 19334 9500 19340 9512
rect 18104 9472 19340 9500
rect 18104 9460 18110 9472
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 20530 9500 20536 9512
rect 20491 9472 20536 9500
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 11072 9404 12480 9432
rect 12704 9435 12762 9441
rect 12704 9401 12716 9435
rect 12750 9432 12762 9435
rect 14734 9432 14740 9444
rect 12750 9404 14740 9432
rect 12750 9401 12762 9404
rect 12704 9395 12762 9401
rect 14734 9392 14740 9404
rect 14792 9392 14798 9444
rect 17586 9392 17592 9444
rect 17644 9432 17650 9444
rect 18294 9435 18352 9441
rect 18294 9432 18306 9435
rect 17644 9404 18306 9432
rect 17644 9392 17650 9404
rect 18294 9401 18306 9404
rect 18340 9401 18352 9435
rect 18294 9395 18352 9401
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 9272 9336 9597 9364
rect 9272 9324 9278 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13780 9336 13829 9364
rect 13780 9324 13786 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 14090 9364 14096 9376
rect 14051 9336 14096 9364
rect 13817 9327 13875 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15930 9364 15936 9376
rect 15068 9336 15113 9364
rect 15891 9336 15936 9364
rect 15068 9324 15074 9336
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16025 9367 16083 9373
rect 16025 9333 16037 9367
rect 16071 9364 16083 9367
rect 16114 9364 16120 9376
rect 16071 9336 16120 9364
rect 16071 9333 16083 9336
rect 16025 9327 16083 9333
rect 16114 9324 16120 9336
rect 16172 9364 16178 9376
rect 17494 9364 17500 9376
rect 16172 9336 17500 9364
rect 16172 9324 16178 9336
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 20070 9364 20076 9376
rect 20031 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20438 9364 20444 9376
rect 20399 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 8941 9163 8999 9169
rect 8941 9129 8953 9163
rect 8987 9160 8999 9163
rect 9674 9160 9680 9172
rect 8987 9132 9680 9160
rect 8987 9129 8999 9132
rect 8941 9123 8999 9129
rect 8588 9092 8616 9123
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 11422 9160 11428 9172
rect 11383 9132 11428 9160
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12437 9163 12495 9169
rect 12437 9160 12449 9163
rect 11756 9132 12449 9160
rect 11756 9120 11762 9132
rect 12437 9129 12449 9132
rect 12483 9129 12495 9163
rect 14090 9160 14096 9172
rect 12437 9123 12495 9129
rect 12636 9132 14096 9160
rect 9766 9092 9772 9104
rect 8588 9064 9772 9092
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 11146 9052 11152 9104
rect 11204 9092 11210 9104
rect 11204 9064 11928 9092
rect 11204 9052 11210 9064
rect 9858 8984 9864 9036
rect 9916 8984 9922 9036
rect 10036 9027 10094 9033
rect 10036 8993 10048 9027
rect 10082 9024 10094 9027
rect 10594 9024 10600 9036
rect 10082 8996 10600 9024
rect 10082 8993 10094 8996
rect 10036 8987 10094 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 10928 8996 11805 9024
rect 10928 8984 10934 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11900 9024 11928 9064
rect 12636 9033 12664 9132
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 17129 9163 17187 9169
rect 17129 9160 17141 9163
rect 16264 9132 17141 9160
rect 16264 9120 16270 9132
rect 17129 9129 17141 9132
rect 17175 9129 17187 9163
rect 17129 9123 17187 9129
rect 17681 9163 17739 9169
rect 17681 9129 17693 9163
rect 17727 9160 17739 9163
rect 17862 9160 17868 9172
rect 17727 9132 17868 9160
rect 17727 9129 17739 9132
rect 17681 9123 17739 9129
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 18049 9163 18107 9169
rect 18049 9129 18061 9163
rect 18095 9160 18107 9163
rect 18095 9132 19932 9160
rect 18095 9129 18107 9132
rect 18049 9123 18107 9129
rect 13256 9095 13314 9101
rect 13256 9061 13268 9095
rect 13302 9092 13314 9095
rect 13722 9092 13728 9104
rect 13302 9064 13728 9092
rect 13302 9061 13314 9064
rect 13256 9055 13314 9061
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 15194 9052 15200 9104
rect 15252 9092 15258 9104
rect 17034 9092 17040 9104
rect 15252 9064 17040 9092
rect 15252 9052 15258 9064
rect 12621 9027 12679 9033
rect 11900 8996 12020 9024
rect 11793 8987 11851 8993
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8260 8928 9045 8956
rect 8260 8916 8266 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 9033 8919 9091 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 9876 8956 9904 8984
rect 11882 8956 11888 8968
rect 9815 8928 9904 8956
rect 11843 8928 11888 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 11992 8965 12020 8996
rect 12621 8993 12633 9027
rect 12667 8993 12679 9027
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12621 8987 12679 8993
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 15764 9033 15792 9064
rect 17034 9052 17040 9064
rect 17092 9052 17098 9104
rect 18960 9095 19018 9101
rect 18960 9092 18972 9095
rect 18616 9064 18972 9092
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 8993 15807 9027
rect 15749 8987 15807 8993
rect 16016 9027 16074 9033
rect 16016 8993 16028 9027
rect 16062 9024 16074 9027
rect 16390 9024 16396 9036
rect 16062 8996 16396 9024
rect 16062 8993 16074 8996
rect 16016 8987 16074 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 17586 9024 17592 9036
rect 17547 8996 17592 9024
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8956 18383 8959
rect 18616 8956 18644 9064
rect 18960 9061 18972 9064
rect 19006 9092 19018 9095
rect 19426 9092 19432 9104
rect 19006 9064 19432 9092
rect 19006 9061 19018 9064
rect 18960 9055 19018 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 19904 9092 19932 9132
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 20349 9163 20407 9169
rect 20349 9160 20361 9163
rect 20036 9132 20361 9160
rect 20036 9120 20042 9132
rect 20349 9129 20361 9132
rect 20395 9129 20407 9163
rect 20349 9123 20407 9129
rect 20530 9092 20536 9104
rect 19904 9064 20536 9092
rect 20530 9052 20536 9064
rect 20588 9052 20594 9104
rect 18693 9027 18751 9033
rect 18693 8993 18705 9027
rect 18739 9024 18751 9027
rect 19334 9024 19340 9036
rect 18739 8996 19340 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 18371 8928 18644 8956
rect 18371 8925 18383 8928
rect 18325 8919 18383 8925
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11149 8891 11207 8897
rect 11149 8888 11161 8891
rect 11020 8860 11161 8888
rect 11020 8848 11026 8860
rect 11149 8857 11161 8860
rect 11195 8857 11207 8891
rect 11149 8851 11207 8857
rect 17034 8848 17040 8900
rect 17092 8888 17098 8900
rect 17405 8891 17463 8897
rect 17405 8888 17417 8891
rect 17092 8860 17417 8888
rect 17092 8848 17098 8860
rect 17405 8857 17417 8860
rect 17451 8888 17463 8891
rect 18046 8888 18052 8900
rect 17451 8860 18052 8888
rect 17451 8857 17463 8860
rect 17405 8851 17463 8857
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 10778 8820 10784 8832
rect 8720 8792 10784 8820
rect 8720 8780 8726 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11606 8780 11612 8832
rect 11664 8820 11670 8832
rect 13630 8820 13636 8832
rect 11664 8792 13636 8820
rect 11664 8780 11670 8792
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 14366 8820 14372 8832
rect 14327 8792 14372 8820
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 18156 8820 18184 8919
rect 19702 8848 19708 8900
rect 19760 8888 19766 8900
rect 20073 8891 20131 8897
rect 20073 8888 20085 8891
rect 19760 8860 20085 8888
rect 19760 8848 19766 8860
rect 20073 8857 20085 8860
rect 20119 8857 20131 8891
rect 20073 8851 20131 8857
rect 19978 8820 19984 8832
rect 18156 8792 19984 8820
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 8202 8616 8208 8628
rect 8163 8588 8208 8616
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 10410 8616 10416 8628
rect 8772 8588 10416 8616
rect 8772 8548 8800 8588
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 16482 8616 16488 8628
rect 15243 8588 16488 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 16482 8576 16488 8588
rect 16540 8616 16546 8628
rect 17586 8616 17592 8628
rect 16540 8588 17592 8616
rect 16540 8576 16546 8588
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 8680 8520 8800 8548
rect 8680 8489 8708 8520
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 11664 8520 12449 8548
rect 11664 8508 11670 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 18601 8551 18659 8557
rect 12437 8511 12495 8517
rect 12636 8520 18184 8548
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8449 8723 8483
rect 8846 8480 8852 8492
rect 8807 8452 8852 8480
rect 8665 8443 8723 8449
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11425 8483 11483 8489
rect 11425 8480 11437 8483
rect 11020 8452 11437 8480
rect 11020 8440 11026 8452
rect 11425 8449 11437 8452
rect 11471 8449 11483 8483
rect 11425 8443 11483 8449
rect 3418 8372 3424 8424
rect 3476 8412 3482 8424
rect 9217 8415 9275 8421
rect 3476 8384 8708 8412
rect 3476 8372 3482 8384
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 8573 8347 8631 8353
rect 8573 8344 8585 8347
rect 6972 8316 8585 8344
rect 6972 8304 6978 8316
rect 8573 8313 8585 8316
rect 8619 8313 8631 8347
rect 8680 8344 8708 8384
rect 9217 8381 9229 8415
rect 9263 8412 9275 8415
rect 9858 8412 9864 8424
rect 9263 8384 9864 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 11333 8415 11391 8421
rect 11333 8412 11345 8415
rect 10152 8384 11345 8412
rect 10152 8356 10180 8384
rect 11333 8381 11345 8384
rect 11379 8412 11391 8415
rect 12066 8412 12072 8424
rect 11379 8384 12072 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 9484 8347 9542 8353
rect 8680 8316 9444 8344
rect 8573 8307 8631 8313
rect 9416 8276 9444 8316
rect 9484 8313 9496 8347
rect 9530 8344 9542 8347
rect 9766 8344 9772 8356
rect 9530 8316 9772 8344
rect 9530 8313 9542 8316
rect 9484 8307 9542 8313
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 10134 8304 10140 8356
rect 10192 8304 10198 8356
rect 11241 8347 11299 8353
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 11885 8347 11943 8353
rect 11885 8344 11897 8347
rect 11287 8316 11897 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 11885 8313 11897 8316
rect 11931 8313 11943 8347
rect 11885 8307 11943 8313
rect 12636 8276 12664 8520
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12768 8452 13001 8480
rect 12768 8440 12774 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 14366 8480 14372 8492
rect 14327 8452 14372 8480
rect 12989 8443 13047 8449
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 16390 8480 16396 8492
rect 16303 8452 16396 8480
rect 16390 8440 16396 8452
rect 16448 8480 16454 8492
rect 16850 8480 16856 8492
rect 16448 8452 16856 8480
rect 16448 8440 16454 8452
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 17184 8452 17233 8480
rect 17184 8440 17190 8452
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 17402 8480 17408 8492
rect 17363 8452 17408 8480
rect 17221 8443 17279 8449
rect 17402 8440 17408 8452
rect 17460 8440 17466 8492
rect 18156 8480 18184 8520
rect 18601 8517 18613 8551
rect 18647 8548 18659 8551
rect 19426 8548 19432 8560
rect 18647 8520 19432 8548
rect 18647 8517 18659 8520
rect 18601 8511 18659 8517
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 18156 8452 19165 8480
rect 19153 8449 19165 8452
rect 19199 8480 19211 8483
rect 20162 8480 20168 8492
rect 19199 8452 20168 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 20622 8480 20628 8492
rect 20303 8452 20628 8480
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 14148 8384 15393 8412
rect 14148 8372 14154 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 18969 8415 19027 8421
rect 18969 8381 18981 8415
rect 19015 8412 19027 8415
rect 20070 8412 20076 8424
rect 19015 8384 20076 8412
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 12802 8344 12808 8356
rect 12763 8316 12808 8344
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 14182 8344 14188 8356
rect 13504 8316 14044 8344
rect 14143 8316 14188 8344
rect 13504 8304 13510 8316
rect 12894 8276 12900 8288
rect 9416 8248 12664 8276
rect 12855 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 13814 8276 13820 8288
rect 13775 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 14016 8276 14044 8316
rect 14182 8304 14188 8316
rect 14240 8304 14246 8356
rect 15562 8304 15568 8356
rect 15620 8344 15626 8356
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 15620 8316 17141 8344
rect 15620 8304 15626 8316
rect 17129 8313 17141 8316
rect 17175 8313 17187 8347
rect 17129 8307 17187 8313
rect 17862 8304 17868 8356
rect 17920 8344 17926 8356
rect 17920 8316 20116 8344
rect 17920 8304 17926 8316
rect 14277 8279 14335 8285
rect 14277 8276 14289 8279
rect 14016 8248 14289 8276
rect 14277 8245 14289 8248
rect 14323 8276 14335 8279
rect 15378 8276 15384 8288
rect 14323 8248 15384 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 15470 8236 15476 8288
rect 15528 8276 15534 8288
rect 15749 8279 15807 8285
rect 15749 8276 15761 8279
rect 15528 8248 15761 8276
rect 15528 8236 15534 8248
rect 15749 8245 15761 8248
rect 15795 8245 15807 8279
rect 16114 8276 16120 8288
rect 16075 8248 16120 8276
rect 15749 8239 15807 8245
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 16264 8248 16309 8276
rect 16264 8236 16270 8248
rect 16390 8236 16396 8288
rect 16448 8276 16454 8288
rect 16761 8279 16819 8285
rect 16761 8276 16773 8279
rect 16448 8248 16773 8276
rect 16448 8236 16454 8248
rect 16761 8245 16773 8248
rect 16807 8245 16819 8279
rect 16761 8239 16819 8245
rect 19061 8279 19119 8285
rect 19061 8245 19073 8279
rect 19107 8276 19119 8279
rect 19613 8279 19671 8285
rect 19613 8276 19625 8279
rect 19107 8248 19625 8276
rect 19107 8245 19119 8248
rect 19061 8239 19119 8245
rect 19613 8245 19625 8248
rect 19659 8245 19671 8279
rect 19978 8276 19984 8288
rect 19939 8248 19984 8276
rect 19613 8239 19671 8245
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 20088 8285 20116 8316
rect 20073 8279 20131 8285
rect 20073 8245 20085 8279
rect 20119 8245 20131 8279
rect 20073 8239 20131 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 11882 8072 11888 8084
rect 9907 8044 11888 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12894 8072 12900 8084
rect 12575 8044 12900 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13814 8072 13820 8084
rect 13372 8044 13820 8072
rect 9125 8007 9183 8013
rect 9125 7973 9137 8007
rect 9171 8004 9183 8007
rect 9950 8004 9956 8016
rect 9171 7976 9956 8004
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 9950 7964 9956 7976
rect 10008 7964 10014 8016
rect 11790 7964 11796 8016
rect 11848 8004 11854 8016
rect 13170 8004 13176 8016
rect 11848 7976 13176 8004
rect 11848 7964 11854 7976
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 8849 7939 8907 7945
rect 8849 7905 8861 7939
rect 8895 7936 8907 7939
rect 9674 7936 9680 7948
rect 8895 7908 9680 7936
rect 8895 7905 8907 7908
rect 8849 7899 8907 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10226 7936 10232 7948
rect 10187 7908 10232 7936
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 10962 7936 10968 7948
rect 10520 7908 10968 7936
rect 10520 7877 10548 7908
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11140 7939 11198 7945
rect 11140 7905 11152 7939
rect 11186 7936 11198 7939
rect 12897 7939 12955 7945
rect 11186 7908 12848 7936
rect 11186 7905 11198 7908
rect 11140 7899 11198 7905
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10870 7868 10876 7880
rect 10831 7840 10876 7868
rect 10505 7831 10563 7837
rect 10336 7800 10364 7831
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 10778 7800 10784 7812
rect 10336 7772 10784 7800
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 12032 7704 12265 7732
rect 12032 7692 12038 7704
rect 12253 7701 12265 7704
rect 12299 7732 12311 7735
rect 12710 7732 12716 7744
rect 12299 7704 12716 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 12820 7732 12848 7908
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13372 7936 13400 8044
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 16114 8072 16120 8084
rect 15703 8044 16120 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 19334 8072 19340 8084
rect 18984 8044 19340 8072
rect 18984 8004 19012 8044
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 20220 8044 20269 8072
rect 20220 8032 20226 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 20257 8035 20315 8041
rect 20438 8032 20444 8084
rect 20496 8072 20502 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20496 8044 20913 8072
rect 20496 8032 20502 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 20901 8035 20959 8041
rect 16684 7976 19012 8004
rect 12943 7908 13400 7936
rect 13808 7939 13866 7945
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13808 7905 13820 7939
rect 13854 7936 13866 7939
rect 14366 7936 14372 7948
rect 13854 7908 14372 7936
rect 13854 7905 13866 7908
rect 13808 7899 13866 7905
rect 14366 7896 14372 7908
rect 14424 7936 14430 7948
rect 14734 7936 14740 7948
rect 14424 7908 14740 7936
rect 14424 7896 14430 7908
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 16022 7936 16028 7948
rect 15983 7908 16028 7936
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7936 16175 7939
rect 16390 7936 16396 7948
rect 16163 7908 16396 7936
rect 16163 7905 16175 7908
rect 16117 7899 16175 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 12986 7868 12992 7880
rect 12947 7840 12992 7868
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13188 7744 13216 7831
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13504 7840 13553 7868
rect 13504 7828 13510 7840
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 16684 7877 16712 7976
rect 16936 7939 16994 7945
rect 16936 7905 16948 7939
rect 16982 7936 16994 7939
rect 17402 7936 17408 7948
rect 16982 7908 17408 7936
rect 16982 7905 16994 7908
rect 16936 7899 16994 7905
rect 17402 7896 17408 7908
rect 17460 7936 17466 7948
rect 18598 7936 18604 7948
rect 17460 7908 18604 7936
rect 17460 7896 17466 7908
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7936 18935 7939
rect 18984 7936 19012 7976
rect 19144 8007 19202 8013
rect 19144 7973 19156 8007
rect 19190 8004 19202 8007
rect 20622 8004 20628 8016
rect 19190 7976 20628 8004
rect 19190 7973 19202 7976
rect 19144 7967 19202 7973
rect 20622 7964 20628 7976
rect 20680 7964 20686 8016
rect 18923 7908 19012 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 15804 7840 16313 7868
rect 15804 7828 15810 7840
rect 16301 7837 16313 7840
rect 16347 7868 16359 7871
rect 16669 7871 16727 7877
rect 16347 7840 16620 7868
rect 16347 7837 16359 7840
rect 16301 7831 16359 7837
rect 13170 7732 13176 7744
rect 12820 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7732 13234 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 13228 7704 14933 7732
rect 13228 7692 13234 7704
rect 14921 7701 14933 7704
rect 14967 7701 14979 7735
rect 16592 7732 16620 7840
rect 16669 7837 16681 7871
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 17586 7732 17592 7744
rect 16592 7704 17592 7732
rect 14921 7695 14979 7701
rect 17586 7692 17592 7704
rect 17644 7732 17650 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 17644 7704 18061 7732
rect 17644 7692 17650 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18049 7695 18107 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10284 7500 10333 7528
rect 10284 7488 10290 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 10778 7488 10784 7540
rect 10836 7528 10842 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 10836 7500 11345 7528
rect 10836 7488 10842 7500
rect 11333 7497 11345 7500
rect 11379 7497 11391 7531
rect 12802 7528 12808 7540
rect 12763 7500 12808 7528
rect 11333 7491 11391 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 12986 7488 12992 7540
rect 13044 7528 13050 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 13044 7500 13829 7528
rect 13044 7488 13050 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 16666 7528 16672 7540
rect 13817 7491 13875 7497
rect 15488 7500 16672 7528
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12342 7460 12348 7472
rect 12124 7432 12348 7460
rect 12124 7420 12130 7432
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 13446 7420 13452 7472
rect 13504 7460 13510 7472
rect 15488 7460 15516 7500
rect 16666 7488 16672 7500
rect 16724 7488 16730 7540
rect 16850 7528 16856 7540
rect 16811 7500 16856 7528
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 13504 7432 15516 7460
rect 13504 7420 13510 7432
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10652 7364 10885 7392
rect 10652 7352 10658 7364
rect 10873 7361 10885 7364
rect 10919 7392 10931 7395
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 10919 7364 11897 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13228 7364 13369 7392
rect 13228 7352 13234 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13780 7364 14289 7392
rect 13780 7352 13786 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14734 7392 14740 7404
rect 14507 7364 14740 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 15488 7401 15516 7432
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 15473 7355 15531 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 20438 7392 20444 7404
rect 20399 7364 20444 7392
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 8386 7324 8392 7336
rect 8347 7296 8392 7324
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7324 11759 7327
rect 13265 7327 13323 7333
rect 11747 7296 13124 7324
rect 11747 7293 11759 7296
rect 11701 7287 11759 7293
rect 8656 7259 8714 7265
rect 8656 7225 8668 7259
rect 8702 7256 8714 7259
rect 9858 7256 9864 7268
rect 8702 7228 9864 7256
rect 8702 7225 8714 7228
rect 8656 7219 8714 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10781 7259 10839 7265
rect 10781 7225 10793 7259
rect 10827 7256 10839 7259
rect 12802 7256 12808 7268
rect 10827 7228 12808 7256
rect 10827 7225 10839 7228
rect 10781 7219 10839 7225
rect 12802 7216 12808 7228
rect 12860 7216 12866 7268
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10686 7188 10692 7200
rect 10008 7160 10692 7188
rect 10008 7148 10014 7160
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 12250 7188 12256 7200
rect 11839 7160 12256 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 13096 7188 13124 7296
rect 13265 7293 13277 7327
rect 13311 7324 13323 7327
rect 13814 7324 13820 7336
rect 13311 7296 13820 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7324 14243 7327
rect 14918 7324 14924 7336
rect 14231 7296 14924 7324
rect 14231 7293 14243 7296
rect 14185 7287 14243 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 15746 7333 15752 7336
rect 15740 7324 15752 7333
rect 15707 7296 15752 7324
rect 15740 7287 15752 7296
rect 15746 7284 15752 7287
rect 15804 7284 15810 7336
rect 16022 7284 16028 7336
rect 16080 7324 16086 7336
rect 17129 7327 17187 7333
rect 17129 7324 17141 7327
rect 16080 7296 17141 7324
rect 16080 7284 16086 7296
rect 17129 7293 17141 7296
rect 17175 7293 17187 7327
rect 17129 7287 17187 7293
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18782 7324 18788 7336
rect 18463 7296 18788 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 20346 7324 20352 7336
rect 20307 7296 20352 7324
rect 20346 7284 20352 7296
rect 20404 7284 20410 7336
rect 13173 7259 13231 7265
rect 13173 7225 13185 7259
rect 13219 7256 13231 7259
rect 14829 7259 14887 7265
rect 14829 7256 14841 7259
rect 13219 7228 14841 7256
rect 13219 7225 13231 7228
rect 13173 7219 13231 7225
rect 14829 7225 14841 7228
rect 14875 7225 14887 7259
rect 14829 7219 14887 7225
rect 15102 7216 15108 7268
rect 15160 7256 15166 7268
rect 18690 7256 18696 7268
rect 15160 7228 18696 7256
rect 15160 7216 15166 7228
rect 18690 7216 18696 7228
rect 18748 7216 18754 7268
rect 15120 7188 15148 7216
rect 18046 7188 18052 7200
rect 13096 7160 15148 7188
rect 18007 7160 18052 7188
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 18782 7188 18788 7200
rect 18555 7160 18788 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 18782 7148 18788 7160
rect 18840 7188 18846 7200
rect 19058 7188 19064 7200
rect 18840 7160 19064 7188
rect 18840 7148 18846 7160
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 19889 7191 19947 7197
rect 19889 7188 19901 7191
rect 19208 7160 19901 7188
rect 19208 7148 19214 7160
rect 19889 7157 19901 7160
rect 19935 7157 19947 7191
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 19889 7151 19947 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 11057 6987 11115 6993
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 12710 6984 12716 6996
rect 11103 6956 12716 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13262 6984 13268 6996
rect 12860 6956 13268 6984
rect 12860 6944 12866 6956
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13814 6984 13820 6996
rect 13775 6956 13820 6984
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 14277 6987 14335 6993
rect 14277 6953 14289 6987
rect 14323 6984 14335 6987
rect 15194 6984 15200 6996
rect 14323 6956 15200 6984
rect 14323 6953 14335 6956
rect 14277 6947 14335 6953
rect 15194 6944 15200 6956
rect 15252 6944 15258 6996
rect 16206 6944 16212 6996
rect 16264 6984 16270 6996
rect 16853 6987 16911 6993
rect 16853 6984 16865 6987
rect 16264 6956 16865 6984
rect 16264 6944 16270 6956
rect 16853 6953 16865 6956
rect 16899 6953 16911 6987
rect 16853 6947 16911 6953
rect 17221 6987 17279 6993
rect 17221 6953 17233 6987
rect 17267 6984 17279 6987
rect 18046 6984 18052 6996
rect 17267 6956 18052 6984
rect 17267 6953 17279 6956
rect 17221 6947 17279 6953
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18230 6984 18236 6996
rect 18191 6956 18236 6984
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 20533 6987 20591 6993
rect 20533 6953 20545 6987
rect 20579 6984 20591 6987
rect 20622 6984 20628 6996
rect 20579 6956 20628 6984
rect 20579 6953 20591 6956
rect 20533 6947 20591 6953
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9824 6888 10180 6916
rect 9824 6876 9830 6888
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10152 6848 10180 6888
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 13906 6916 13912 6928
rect 10744 6888 13912 6916
rect 10744 6876 10750 6888
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 14090 6876 14096 6928
rect 14148 6916 14154 6928
rect 15657 6919 15715 6925
rect 15657 6916 15669 6919
rect 14148 6888 15669 6916
rect 14148 6876 14154 6888
rect 15657 6885 15669 6888
rect 15703 6916 15715 6919
rect 18506 6916 18512 6928
rect 15703 6888 18512 6916
rect 15703 6885 15715 6888
rect 15657 6879 15715 6885
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 11149 6851 11207 6857
rect 10152 6820 10272 6848
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9674 6780 9680 6792
rect 9171 6752 9680 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 10244 6789 10272 6820
rect 11149 6817 11161 6851
rect 11195 6848 11207 6851
rect 11330 6848 11336 6860
rect 11195 6820 11336 6848
rect 11195 6817 11207 6820
rect 11149 6811 11207 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11965 6857 11971 6860
rect 11957 6851 11971 6857
rect 11957 6848 11969 6851
rect 11926 6820 11969 6848
rect 11957 6817 11969 6820
rect 11957 6811 11971 6817
rect 11965 6808 11971 6811
rect 12023 6808 12029 6860
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 13504 6820 14197 6848
rect 13504 6808 13510 6820
rect 14185 6817 14197 6820
rect 14231 6848 14243 6851
rect 15562 6848 15568 6860
rect 14231 6820 15568 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 16022 6848 16028 6860
rect 15795 6820 16028 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16482 6848 16488 6860
rect 16443 6820 16488 6848
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 17218 6808 17224 6860
rect 17276 6848 17282 6860
rect 18325 6851 18383 6857
rect 18325 6848 18337 6851
rect 17276 6820 18337 6848
rect 17276 6808 17282 6820
rect 18325 6817 18337 6820
rect 18371 6817 18383 6851
rect 18325 6811 18383 6817
rect 19420 6851 19478 6857
rect 19420 6817 19432 6851
rect 19466 6848 19478 6851
rect 19794 6848 19800 6860
rect 19466 6820 19800 6848
rect 19466 6817 19478 6820
rect 19420 6811 19478 6817
rect 19794 6808 19800 6820
rect 19852 6848 19858 6860
rect 20622 6848 20628 6860
rect 19852 6820 20628 6848
rect 19852 6808 19858 6820
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9824 6752 10149 6780
rect 9824 6740 9830 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 11020 6752 11253 6780
rect 11020 6740 11026 6752
rect 11241 6749 11253 6752
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6749 11759 6783
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 11701 6743 11759 6749
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 11716 6712 11744 6743
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 15838 6780 15844 6792
rect 15799 6752 15844 6780
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 17236 6780 17264 6808
rect 16264 6752 17264 6780
rect 17313 6783 17371 6789
rect 16264 6740 16270 6752
rect 17313 6749 17325 6783
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17586 6780 17592 6792
rect 17543 6752 17592 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 14568 6712 14596 6740
rect 10928 6684 11744 6712
rect 13004 6684 14596 6712
rect 10928 6672 10934 6684
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10192 6616 10701 6644
rect 10192 6604 10198 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 13004 6644 13032 6684
rect 15378 6672 15384 6724
rect 15436 6712 15442 6724
rect 15562 6712 15568 6724
rect 15436 6684 15568 6712
rect 15436 6672 15442 6684
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 17328 6712 17356 6743
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18598 6780 18604 6792
rect 18555 6752 18604 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19153 6783 19211 6789
rect 19153 6780 19165 6783
rect 19116 6752 19165 6780
rect 19116 6740 19122 6752
rect 19153 6749 19165 6752
rect 19199 6749 19211 6783
rect 19153 6743 19211 6749
rect 17865 6715 17923 6721
rect 17865 6712 17877 6715
rect 17328 6684 17877 6712
rect 17865 6681 17877 6684
rect 17911 6681 17923 6715
rect 17865 6675 17923 6681
rect 11940 6616 13032 6644
rect 13081 6647 13139 6653
rect 11940 6604 11946 6616
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 13170 6644 13176 6656
rect 13127 6616 13176 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 15289 6647 15347 6653
rect 15289 6644 15301 6647
rect 14608 6616 15301 6644
rect 14608 6604 14614 6616
rect 15289 6613 15301 6616
rect 15335 6613 15347 6647
rect 15289 6607 15347 6613
rect 16301 6647 16359 6653
rect 16301 6613 16313 6647
rect 16347 6644 16359 6647
rect 16666 6644 16672 6656
rect 16347 6616 16672 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 9858 6440 9864 6452
rect 9819 6412 9864 6440
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 10100 6412 10149 6440
rect 10100 6400 10106 6412
rect 10137 6409 10149 6412
rect 10183 6409 10195 6443
rect 10137 6403 10195 6409
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 13538 6440 13544 6452
rect 11848 6412 13544 6440
rect 11848 6400 11854 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 18233 6443 18291 6449
rect 18233 6409 18245 6443
rect 18279 6440 18291 6443
rect 19610 6440 19616 6452
rect 18279 6412 19616 6440
rect 18279 6409 18291 6412
rect 18233 6403 18291 6409
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 20622 6440 20628 6452
rect 20583 6412 20628 6440
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 9876 6304 9904 6400
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 15286 6372 15292 6384
rect 12308 6344 15292 6372
rect 12308 6332 12314 6344
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 10318 6304 10324 6316
rect 9876 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6304 10382 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10376 6276 10701 6304
rect 10376 6264 10382 6276
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11020 6276 11713 6304
rect 11020 6264 11026 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 13078 6304 13084 6316
rect 13039 6276 13084 6304
rect 11701 6267 11759 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13228 6276 14105 6304
rect 13228 6264 13234 6276
rect 14093 6273 14105 6276
rect 14139 6304 14151 6307
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14139 6276 15025 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 17126 6304 17132 6316
rect 16347 6276 17132 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 18877 6307 18935 6313
rect 17276 6276 17321 6304
rect 17276 6264 17282 6276
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 18966 6304 18972 6316
rect 18923 6276 18972 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 8386 6236 8392 6248
rect 6871 6208 8392 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 8386 6196 8392 6208
rect 8444 6236 8450 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8444 6208 8493 6236
rect 8444 6196 8450 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9732 6208 10517 6236
rect 9732 6196 9738 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10652 6208 11100 6236
rect 10652 6196 10658 6208
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 7070 6171 7128 6177
rect 7070 6168 7082 6171
rect 4120 6140 7082 6168
rect 4120 6128 4126 6140
rect 7070 6137 7082 6140
rect 7116 6137 7128 6171
rect 8726 6171 8784 6177
rect 8726 6168 8738 6171
rect 7070 6131 7128 6137
rect 8220 6140 8738 6168
rect 8220 6109 8248 6140
rect 8726 6137 8738 6140
rect 8772 6168 8784 6171
rect 10962 6168 10968 6180
rect 8772 6140 10968 6168
rect 8772 6137 8784 6140
rect 8726 6131 8784 6137
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 11072 6168 11100 6208
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11204 6208 11621 6236
rect 11204 6196 11210 6208
rect 11609 6205 11621 6208
rect 11655 6236 11667 6239
rect 11882 6236 11888 6248
rect 11655 6208 11888 6236
rect 11655 6205 11667 6208
rect 11609 6199 11667 6205
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6236 13967 6239
rect 13998 6236 14004 6248
rect 13955 6208 14004 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 14240 6208 16129 6236
rect 14240 6196 14246 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 19058 6236 19064 6248
rect 18564 6208 19064 6236
rect 18564 6196 18570 6208
rect 19058 6196 19064 6208
rect 19116 6236 19122 6248
rect 19245 6239 19303 6245
rect 19245 6236 19257 6239
rect 19116 6208 19257 6236
rect 19116 6196 19122 6208
rect 19245 6205 19257 6208
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 19512 6239 19570 6245
rect 19512 6205 19524 6239
rect 19558 6236 19570 6239
rect 19886 6236 19892 6248
rect 19558 6208 19892 6236
rect 19558 6205 19570 6208
rect 19512 6199 19570 6205
rect 19886 6196 19892 6208
rect 19944 6236 19950 6248
rect 20438 6236 20444 6248
rect 19944 6208 20444 6236
rect 19944 6196 19950 6208
rect 20438 6196 20444 6208
rect 20496 6196 20502 6248
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 11072 6140 11529 6168
rect 11517 6137 11529 6140
rect 11563 6168 11575 6171
rect 11790 6168 11796 6180
rect 11563 6140 11796 6168
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 12805 6171 12863 6177
rect 12805 6137 12817 6171
rect 12851 6168 12863 6171
rect 14829 6171 14887 6177
rect 12851 6140 14504 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6069 8263 6103
rect 8205 6063 8263 6069
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 10643 6072 11161 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12897 6103 12955 6109
rect 12492 6072 12537 6100
rect 12492 6060 12498 6072
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 12943 6072 13461 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13449 6069 13461 6072
rect 13495 6069 13507 6103
rect 13449 6063 13507 6069
rect 13817 6103 13875 6109
rect 13817 6069 13829 6103
rect 13863 6100 13875 6103
rect 13906 6100 13912 6112
rect 13863 6072 13912 6100
rect 13863 6069 13875 6072
rect 13817 6063 13875 6069
rect 13906 6060 13912 6072
rect 13964 6100 13970 6112
rect 14274 6100 14280 6112
rect 13964 6072 14280 6100
rect 13964 6060 13970 6072
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 14476 6109 14504 6140
rect 14829 6137 14841 6171
rect 14875 6168 14887 6171
rect 15102 6168 15108 6180
rect 14875 6140 15108 6168
rect 14875 6137 14887 6140
rect 14829 6131 14887 6137
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 16071 6140 16712 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 15286 6100 15292 6112
rect 14967 6072 15292 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 15746 6100 15752 6112
rect 15703 6072 15752 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16684 6109 16712 6140
rect 16850 6128 16856 6180
rect 16908 6168 16914 6180
rect 17129 6171 17187 6177
rect 17129 6168 17141 6171
rect 16908 6140 17141 6168
rect 16908 6128 16914 6140
rect 17129 6137 17141 6140
rect 17175 6168 17187 6171
rect 17954 6168 17960 6180
rect 17175 6140 17960 6168
rect 17175 6137 17187 6140
rect 17129 6131 17187 6137
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 18601 6171 18659 6177
rect 18601 6137 18613 6171
rect 18647 6168 18659 6171
rect 18647 6140 19288 6168
rect 18647 6137 18659 6140
rect 18601 6131 18659 6137
rect 19260 6112 19288 6140
rect 16669 6103 16727 6109
rect 16669 6069 16681 6103
rect 16715 6069 16727 6103
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 16669 6063 16727 6069
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 18748 6072 18793 6100
rect 18748 6060 18754 6072
rect 19242 6060 19248 6112
rect 19300 6060 19306 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 9766 5896 9772 5908
rect 9727 5868 9772 5896
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10134 5896 10140 5908
rect 10095 5868 10140 5896
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 12492 5868 13093 5896
rect 12492 5856 12498 5868
rect 13081 5865 13093 5868
rect 13127 5865 13139 5899
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 13081 5859 13139 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14550 5896 14556 5908
rect 14511 5868 14556 5896
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15013 5899 15071 5905
rect 15013 5865 15025 5899
rect 15059 5896 15071 5899
rect 16482 5896 16488 5908
rect 15059 5868 16488 5896
rect 15059 5865 15071 5868
rect 15013 5859 15071 5865
rect 16482 5856 16488 5868
rect 16540 5896 16546 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 16540 5868 16681 5896
rect 16540 5856 16546 5868
rect 16669 5865 16681 5868
rect 16715 5896 16727 5899
rect 17218 5896 17224 5908
rect 16715 5868 17224 5896
rect 16715 5865 16727 5868
rect 16669 5859 16727 5865
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 18598 5896 18604 5908
rect 18559 5868 18604 5896
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 18966 5856 18972 5908
rect 19024 5896 19030 5908
rect 19518 5896 19524 5908
rect 19024 5868 19524 5896
rect 19024 5856 19030 5868
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20312 5868 20913 5896
rect 20312 5856 20318 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 11232 5831 11290 5837
rect 11232 5797 11244 5831
rect 11278 5828 11290 5831
rect 13170 5828 13176 5840
rect 11278 5800 13176 5828
rect 11278 5797 11290 5800
rect 11232 5791 11290 5797
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 15378 5828 15384 5840
rect 14056 5800 15384 5828
rect 14056 5788 14062 5800
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 15556 5831 15614 5837
rect 15556 5797 15568 5831
rect 15602 5828 15614 5831
rect 15838 5828 15844 5840
rect 15602 5800 15844 5828
rect 15602 5797 15614 5800
rect 15556 5791 15614 5797
rect 15838 5788 15844 5800
rect 15896 5788 15902 5840
rect 17126 5788 17132 5840
rect 17184 5828 17190 5840
rect 19122 5831 19180 5837
rect 19122 5828 19134 5831
rect 17184 5800 19134 5828
rect 17184 5788 17190 5800
rect 19122 5797 19134 5800
rect 19168 5797 19180 5831
rect 19122 5791 19180 5797
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 10870 5760 10876 5772
rect 8444 5732 10876 5760
rect 8444 5720 8450 5732
rect 10870 5720 10876 5732
rect 10928 5760 10934 5772
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10928 5732 10977 5760
rect 10928 5720 10934 5732
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 12986 5760 12992 5772
rect 12947 5732 12992 5760
rect 10965 5723 11023 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15194 5760 15200 5772
rect 14691 5732 15200 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 17488 5763 17546 5769
rect 15335 5732 16712 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 10226 5692 10232 5704
rect 10187 5664 10232 5692
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 13262 5692 13268 5704
rect 10376 5664 10421 5692
rect 13223 5664 13268 5692
rect 10376 5652 10382 5664
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13630 5692 13636 5704
rect 13591 5664 13636 5692
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 14875 5664 15025 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15304 5692 15332 5723
rect 16684 5704 16712 5732
rect 17488 5729 17500 5763
rect 17534 5760 17546 5763
rect 17954 5760 17960 5772
rect 17534 5732 17960 5760
rect 17534 5729 17546 5732
rect 17488 5723 17546 5729
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 15160 5664 15332 5692
rect 15160 5652 15166 5664
rect 16666 5652 16672 5704
rect 16724 5692 16730 5704
rect 17218 5692 17224 5704
rect 16724 5664 17224 5692
rect 16724 5652 16730 5664
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 18506 5652 18512 5704
rect 18564 5692 18570 5704
rect 18877 5695 18935 5701
rect 18877 5692 18889 5695
rect 18564 5664 18889 5692
rect 18564 5652 18570 5664
rect 18877 5661 18889 5664
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 12345 5627 12403 5633
rect 12345 5593 12357 5627
rect 12391 5624 12403 5627
rect 13078 5624 13084 5636
rect 12391 5596 13084 5624
rect 12391 5593 12403 5596
rect 12345 5587 12403 5593
rect 13078 5584 13084 5596
rect 13136 5584 13142 5636
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 16574 5624 16580 5636
rect 16356 5596 16580 5624
rect 16356 5584 16362 5596
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 12621 5559 12679 5565
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 13538 5556 13544 5568
rect 12667 5528 13544 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 19978 5556 19984 5568
rect 13964 5528 19984 5556
rect 13964 5516 13970 5528
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 10226 5312 10232 5364
rect 10284 5352 10290 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10284 5324 10425 5352
rect 10284 5312 10290 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 10928 5324 11345 5352
rect 10928 5312 10934 5324
rect 11333 5321 11345 5324
rect 11379 5352 11391 5355
rect 11425 5355 11483 5361
rect 11425 5352 11437 5355
rect 11379 5324 11437 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11425 5321 11437 5324
rect 11471 5321 11483 5355
rect 11425 5315 11483 5321
rect 12529 5355 12587 5361
rect 12529 5321 12541 5355
rect 12575 5352 12587 5355
rect 12986 5352 12992 5364
rect 12575 5324 12992 5352
rect 12575 5321 12587 5324
rect 12529 5315 12587 5321
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 15105 5355 15163 5361
rect 15105 5321 15117 5355
rect 15151 5352 15163 5355
rect 15838 5352 15844 5364
rect 15151 5324 15844 5352
rect 15151 5321 15163 5324
rect 15105 5315 15163 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17313 5355 17371 5361
rect 17313 5352 17325 5355
rect 17184 5324 17325 5352
rect 17184 5312 17190 5324
rect 17313 5321 17325 5324
rect 17359 5321 17371 5355
rect 19886 5352 19892 5364
rect 19847 5324 19892 5352
rect 17313 5315 17371 5321
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 20165 5287 20223 5293
rect 20165 5253 20177 5287
rect 20211 5284 20223 5287
rect 20438 5284 20444 5296
rect 20211 5256 20444 5284
rect 20211 5253 20223 5256
rect 20165 5247 20223 5253
rect 20438 5244 20444 5256
rect 20496 5244 20502 5296
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 13078 5216 13084 5228
rect 13039 5188 13084 5216
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 15562 5216 15568 5228
rect 15120 5188 15568 5216
rect 10796 5148 10824 5176
rect 15120 5160 15148 5188
rect 15562 5176 15568 5188
rect 15620 5216 15626 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15620 5188 15945 5216
rect 15620 5176 15626 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 17862 5216 17868 5228
rect 17276 5188 17868 5216
rect 17276 5176 17282 5188
rect 17862 5176 17868 5188
rect 17920 5216 17926 5228
rect 18506 5216 18512 5228
rect 17920 5188 18512 5216
rect 17920 5176 17926 5188
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 20272 5188 20729 5216
rect 20272 5160 20300 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10796 5120 10885 5148
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5148 11667 5151
rect 11698 5148 11704 5160
rect 11655 5120 11704 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13630 5148 13636 5160
rect 12943 5120 13636 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 15102 5148 15108 5160
rect 13771 5120 15108 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 15102 5108 15108 5120
rect 15160 5108 15166 5160
rect 15378 5148 15384 5160
rect 15339 5120 15384 5148
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 16200 5151 16258 5157
rect 16200 5117 16212 5151
rect 16246 5148 16258 5151
rect 16482 5148 16488 5160
rect 16246 5120 16488 5148
rect 16246 5117 16258 5120
rect 16200 5111 16258 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 18776 5151 18834 5157
rect 18776 5117 18788 5151
rect 18822 5148 18834 5151
rect 20254 5148 20260 5160
rect 18822 5120 20260 5148
rect 18822 5117 18834 5120
rect 18776 5111 18834 5117
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 10781 5083 10839 5089
rect 10781 5049 10793 5083
rect 10827 5080 10839 5083
rect 10827 5052 13216 5080
rect 10827 5049 10839 5052
rect 10781 5043 10839 5049
rect 11333 5015 11391 5021
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 11698 5012 11704 5024
rect 11379 4984 11704 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 13188 5012 13216 5052
rect 13262 5040 13268 5092
rect 13320 5080 13326 5092
rect 13970 5083 14028 5089
rect 13970 5080 13982 5083
rect 13320 5052 13982 5080
rect 13320 5040 13326 5052
rect 13970 5049 13982 5052
rect 14016 5049 14028 5083
rect 16022 5080 16028 5092
rect 13970 5043 14028 5049
rect 14292 5052 16028 5080
rect 14292 5012 14320 5052
rect 16022 5040 16028 5052
rect 16080 5080 16086 5092
rect 18598 5080 18604 5092
rect 16080 5052 18604 5080
rect 16080 5040 16086 5052
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 20070 5040 20076 5092
rect 20128 5080 20134 5092
rect 20533 5083 20591 5089
rect 20533 5080 20545 5083
rect 20128 5052 20545 5080
rect 20128 5040 20134 5052
rect 20533 5049 20545 5052
rect 20579 5080 20591 5083
rect 20714 5080 20720 5092
rect 20579 5052 20720 5080
rect 20579 5049 20591 5052
rect 20533 5043 20591 5049
rect 20714 5040 20720 5052
rect 20772 5040 20778 5092
rect 13044 4984 13089 5012
rect 13188 4984 14320 5012
rect 15565 5015 15623 5021
rect 13044 4972 13050 4984
rect 15565 4981 15577 5015
rect 15611 5012 15623 5015
rect 15838 5012 15844 5024
rect 15611 4984 15844 5012
rect 15611 4981 15623 4984
rect 15565 4975 15623 4981
rect 15838 4972 15844 4984
rect 15896 4972 15902 5024
rect 17770 4972 17776 5024
rect 17828 5012 17834 5024
rect 20625 5015 20683 5021
rect 20625 5012 20637 5015
rect 17828 4984 20637 5012
rect 17828 4972 17834 4984
rect 20625 4981 20637 4984
rect 20671 4981 20683 5015
rect 20625 4975 20683 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6144 4780 13216 4808
rect 6144 4768 6150 4780
rect 12520 4743 12578 4749
rect 12520 4709 12532 4743
rect 12566 4740 12578 4743
rect 13078 4740 13084 4752
rect 12566 4712 13084 4740
rect 12566 4709 12578 4712
rect 12520 4703 12578 4709
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 13188 4740 13216 4780
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13320 4780 13645 4808
rect 13320 4768 13326 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 15252 4780 15301 4808
rect 15252 4768 15258 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 15657 4811 15715 4817
rect 15657 4777 15669 4811
rect 15703 4808 15715 4811
rect 16301 4811 16359 4817
rect 15703 4780 16252 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 16224 4740 16252 4780
rect 16301 4777 16313 4811
rect 16347 4808 16359 4811
rect 17034 4808 17040 4820
rect 16347 4780 17040 4808
rect 16347 4777 16359 4780
rect 16301 4771 16359 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 18782 4808 18788 4820
rect 17819 4780 18788 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 19150 4808 19156 4820
rect 19111 4780 19156 4808
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 19242 4768 19248 4820
rect 19300 4808 19306 4820
rect 20165 4811 20223 4817
rect 20165 4808 20177 4811
rect 19300 4780 20177 4808
rect 19300 4768 19306 4780
rect 20165 4777 20177 4780
rect 20211 4777 20223 4811
rect 20165 4771 20223 4777
rect 16758 4740 16764 4752
rect 13188 4712 15792 4740
rect 16224 4712 16764 4740
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 11756 4644 12265 4672
rect 11756 4632 11762 4644
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 12253 4635 12311 4641
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 13909 4675 13967 4681
rect 13909 4672 13921 4675
rect 13872 4644 13921 4672
rect 13872 4632 13878 4644
rect 13909 4641 13921 4644
rect 13955 4641 13967 4675
rect 13909 4635 13967 4641
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 15764 4681 15792 4712
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 17954 4700 17960 4752
rect 18012 4740 18018 4752
rect 18012 4712 18368 4740
rect 18012 4700 18018 4712
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 14056 4644 14565 4672
rect 14056 4632 14062 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 15749 4675 15807 4681
rect 15749 4641 15761 4675
rect 15795 4672 15807 4675
rect 16574 4672 16580 4684
rect 15795 4644 16580 4672
rect 15795 4641 15807 4644
rect 15749 4635 15807 4641
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 15930 4604 15936 4616
rect 15891 4576 15936 4604
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 16776 4604 16804 4700
rect 17313 4675 17371 4681
rect 17313 4641 17325 4675
rect 17359 4672 17371 4675
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 17359 4644 18153 4672
rect 17359 4641 17371 4644
rect 17313 4635 17371 4641
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 16776 4576 17908 4604
rect 17770 4536 17776 4548
rect 14016 4508 17776 4536
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 14016 4468 14044 4508
rect 17770 4496 17776 4508
rect 17828 4496 17834 4548
rect 17880 4536 17908 4576
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18340 4613 18368 4712
rect 18690 4700 18696 4752
rect 18748 4740 18754 4752
rect 18748 4712 20300 4740
rect 18748 4700 18754 4712
rect 19245 4675 19303 4681
rect 19245 4641 19257 4675
rect 19291 4672 19303 4675
rect 19702 4672 19708 4684
rect 19291 4644 19708 4672
rect 19291 4641 19303 4644
rect 19245 4635 19303 4641
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 20272 4616 20300 4712
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 18012 4576 18245 4604
rect 18012 4564 18018 4576
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 19150 4604 19156 4616
rect 18371 4576 19156 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 19794 4604 19800 4616
rect 19475 4576 19800 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 20254 4604 20260 4616
rect 20215 4576 20260 4604
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 20346 4564 20352 4616
rect 20404 4604 20410 4616
rect 20404 4576 20449 4604
rect 20404 4564 20410 4576
rect 20530 4536 20536 4548
rect 17880 4508 20536 4536
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 7524 4440 14044 4468
rect 14093 4471 14151 4477
rect 7524 4428 7530 4440
rect 14093 4437 14105 4471
rect 14139 4468 14151 4471
rect 14182 4468 14188 4480
rect 14139 4440 14188 4468
rect 14139 4437 14151 4440
rect 14093 4431 14151 4437
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 14737 4471 14795 4477
rect 14737 4437 14749 4471
rect 14783 4468 14795 4471
rect 15286 4468 15292 4480
rect 14783 4440 15292 4468
rect 14783 4437 14795 4440
rect 14737 4431 14795 4437
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 18785 4471 18843 4477
rect 18785 4437 18797 4471
rect 18831 4468 18843 4471
rect 19058 4468 19064 4480
rect 18831 4440 19064 4468
rect 18831 4437 18843 4440
rect 18785 4431 18843 4437
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 12805 4267 12863 4273
rect 12805 4233 12817 4267
rect 12851 4264 12863 4267
rect 12986 4264 12992 4276
rect 12851 4236 12992 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 12986 4224 12992 4236
rect 13044 4224 13050 4276
rect 19702 4264 19708 4276
rect 19663 4236 19708 4264
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 11296 4168 11560 4196
rect 11296 4156 11302 4168
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 8938 4128 8944 4140
rect 5316 4100 8944 4128
rect 5316 4088 5322 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 11146 4128 11152 4140
rect 10192 4100 11152 4128
rect 10192 4088 10198 4100
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 11422 4128 11428 4140
rect 11383 4100 11428 4128
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 11532 4128 11560 4168
rect 13170 4156 13176 4208
rect 13228 4196 13234 4208
rect 14001 4199 14059 4205
rect 13228 4168 13400 4196
rect 13228 4156 13234 4168
rect 12894 4128 12900 4140
rect 11532 4100 12900 4128
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13372 4137 13400 4168
rect 14001 4165 14013 4199
rect 14047 4165 14059 4199
rect 14001 4159 14059 4165
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4097 13415 4131
rect 14016 4128 14044 4159
rect 19886 4156 19892 4208
rect 19944 4196 19950 4208
rect 19944 4168 20300 4196
rect 19944 4156 19950 4168
rect 14366 4128 14372 4140
rect 14016 4100 14372 4128
rect 13357 4091 13415 4097
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 17310 4088 17316 4140
rect 17368 4128 17374 4140
rect 20272 4137 20300 4168
rect 20257 4131 20315 4137
rect 17368 4100 18184 4128
rect 17368 4088 17374 4100
rect 842 4020 848 4072
rect 900 4060 906 4072
rect 7558 4060 7564 4072
rect 900 4032 7564 4060
rect 900 4020 906 4032
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8444 4032 9137 4060
rect 8444 4020 8450 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 9381 4063 9439 4069
rect 9381 4060 9393 4063
rect 9272 4032 9393 4060
rect 9272 4020 9278 4032
rect 9381 4029 9393 4032
rect 9427 4029 9439 4063
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 9381 4023 9439 4029
rect 10244 4032 13185 4060
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 7466 3992 7472 4004
rect 2556 3964 7472 3992
rect 2556 3952 2562 3964
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 10042 3992 10048 4004
rect 8260 3964 10048 3992
rect 8260 3952 8266 3964
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 290 3884 296 3936
rect 348 3924 354 3936
rect 10244 3924 10272 4032
rect 13173 4029 13185 4032
rect 13219 4060 13231 4063
rect 13446 4060 13452 4072
rect 13219 4032 13452 4060
rect 13219 4029 13231 4032
rect 13173 4023 13231 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 15010 4060 15016 4072
rect 14971 4032 15016 4060
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15746 4060 15752 4072
rect 15707 4032 15752 4060
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4060 16083 4063
rect 16485 4063 16543 4069
rect 16485 4060 16497 4063
rect 16071 4032 16497 4060
rect 16071 4029 16083 4032
rect 16025 4023 16083 4029
rect 16485 4029 16497 4032
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17678 4060 17684 4072
rect 17451 4032 17684 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 17678 4020 17684 4032
rect 17736 4020 17742 4072
rect 17862 4020 17868 4072
rect 17920 4060 17926 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17920 4032 18061 4060
rect 17920 4020 17926 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18156 4060 18184 4100
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 18690 4060 18696 4072
rect 18156 4032 18696 4060
rect 18049 4023 18107 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19794 4020 19800 4072
rect 19852 4060 19858 4072
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 19852 4032 20085 4060
rect 19852 4020 19858 4032
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4060 20223 4063
rect 20438 4060 20444 4072
rect 20211 4032 20444 4060
rect 20211 4029 20223 4032
rect 20165 4023 20223 4029
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 20714 4060 20720 4072
rect 20675 4032 20720 4060
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 11149 3995 11207 4001
rect 10468 3964 10824 3992
rect 10468 3952 10474 3964
rect 348 3896 10272 3924
rect 348 3884 354 3896
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10796 3933 10824 3964
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 11793 3995 11851 4001
rect 11793 3992 11805 3995
rect 11195 3964 11805 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 11793 3961 11805 3964
rect 11839 3961 11851 3995
rect 11793 3955 11851 3961
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 13265 3995 13323 4001
rect 13265 3992 13277 3995
rect 12860 3964 13277 3992
rect 12860 3952 12866 3964
rect 13265 3961 13277 3964
rect 13311 3961 13323 3995
rect 13265 3955 13323 3961
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 13412 3964 14473 3992
rect 13412 3952 13418 3964
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 14461 3955 14519 3961
rect 17218 3952 17224 4004
rect 17276 3992 17282 4004
rect 17880 3992 17908 4020
rect 17276 3964 17908 3992
rect 18316 3995 18374 4001
rect 17276 3952 17282 3964
rect 18316 3961 18328 3995
rect 18362 3992 18374 3995
rect 18598 3992 18604 4004
rect 18362 3964 18604 3992
rect 18362 3961 18374 3964
rect 18316 3955 18374 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10376 3896 10517 3924
rect 10376 3884 10382 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 10781 3927 10839 3933
rect 10781 3893 10793 3927
rect 10827 3893 10839 3927
rect 10781 3887 10839 3893
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10928 3896 11253 3924
rect 10928 3884 10934 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 14366 3924 14372 3936
rect 14327 3896 14372 3924
rect 11241 3887 11299 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 15068 3896 15209 3924
rect 15068 3884 15074 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 16448 3896 16681 3924
rect 16448 3884 16454 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 17862 3924 17868 3936
rect 17635 3896 17868 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 19208 3896 19441 3924
rect 19208 3884 19214 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19429 3887 19487 3893
rect 20901 3927 20959 3933
rect 20901 3893 20913 3927
rect 20947 3924 20959 3927
rect 22462 3924 22468 3936
rect 20947 3896 22468 3924
rect 20947 3893 20959 3896
rect 20901 3887 20959 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 11238 3720 11244 3732
rect 3660 3692 11244 3720
rect 3660 3680 3666 3692
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 11756 3692 13400 3720
rect 11756 3680 11762 3692
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 11440 3652 11468 3680
rect 11946 3655 12004 3661
rect 11946 3652 11958 3655
rect 7616 3624 10456 3652
rect 11440 3624 11958 3652
rect 7616 3612 7622 3624
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 10134 3584 10140 3596
rect 2004 3556 10140 3584
rect 2004 3544 2010 3556
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10318 3593 10324 3596
rect 10312 3584 10324 3593
rect 10279 3556 10324 3584
rect 10312 3547 10324 3556
rect 10318 3544 10324 3547
rect 10376 3544 10382 3596
rect 10428 3584 10456 3624
rect 11946 3621 11958 3624
rect 11992 3621 12004 3655
rect 11946 3615 12004 3621
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 13262 3652 13268 3664
rect 12492 3624 13268 3652
rect 12492 3612 12498 3624
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 13372 3593 13400 3692
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 14608 3692 14749 3720
rect 14608 3680 14614 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 16114 3720 16120 3732
rect 14737 3683 14795 3689
rect 15488 3692 16120 3720
rect 13446 3612 13452 3664
rect 13504 3652 13510 3664
rect 15488 3652 15516 3692
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16945 3723 17003 3729
rect 16945 3689 16957 3723
rect 16991 3689 17003 3723
rect 18598 3720 18604 3732
rect 18559 3692 18604 3720
rect 16945 3683 17003 3689
rect 13504 3624 15516 3652
rect 16960 3652 16988 3683
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 17126 3652 17132 3664
rect 16960 3624 17132 3652
rect 13504 3612 13510 3624
rect 17126 3612 17132 3624
rect 17184 3652 17190 3664
rect 17466 3655 17524 3661
rect 17466 3652 17478 3655
rect 17184 3624 17478 3652
rect 17184 3612 17190 3624
rect 17466 3621 17478 3624
rect 17512 3621 17524 3655
rect 17466 3615 17524 3621
rect 13357 3587 13415 3593
rect 10428 3556 13032 3584
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 8444 3488 10057 3516
rect 8444 3476 8450 3488
rect 10045 3485 10057 3488
rect 10091 3485 10103 3519
rect 11698 3516 11704 3528
rect 11659 3488 11704 3516
rect 10045 3479 10103 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 3050 3408 3056 3460
rect 3108 3448 3114 3460
rect 9950 3448 9956 3460
rect 3108 3420 9956 3448
rect 3108 3408 3114 3420
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 12342 3380 12348 3392
rect 4212 3352 12348 3380
rect 4212 3340 4218 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 13004 3380 13032 3556
rect 13357 3553 13369 3587
rect 13403 3553 13415 3587
rect 13613 3587 13671 3593
rect 13613 3584 13625 3587
rect 13357 3547 13415 3553
rect 13464 3556 13625 3584
rect 13464 3516 13492 3556
rect 13613 3553 13625 3556
rect 13659 3584 13671 3587
rect 13906 3584 13912 3596
rect 13659 3556 13912 3584
rect 13659 3553 13671 3556
rect 13613 3547 13671 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 15562 3584 15568 3596
rect 14516 3556 15568 3584
rect 14516 3544 14522 3556
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 15832 3587 15890 3593
rect 15832 3553 15844 3587
rect 15878 3584 15890 3587
rect 16114 3584 16120 3596
rect 15878 3556 16120 3584
rect 15878 3553 15890 3556
rect 15832 3547 15890 3553
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 17218 3584 17224 3596
rect 17179 3556 17224 3584
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 19058 3584 19064 3596
rect 19019 3556 19064 3584
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 19797 3587 19855 3593
rect 19797 3584 19809 3587
rect 19484 3556 19809 3584
rect 19484 3544 19490 3556
rect 19797 3553 19809 3556
rect 19843 3553 19855 3587
rect 19797 3547 19855 3553
rect 13096 3488 13492 3516
rect 19337 3519 19395 3525
rect 13096 3457 13124 3488
rect 19337 3485 19349 3519
rect 19383 3516 19395 3519
rect 19518 3516 19524 3528
rect 19383 3488 19524 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20346 3516 20352 3528
rect 20119 3488 20352 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 13081 3451 13139 3457
rect 13081 3417 13093 3451
rect 13127 3417 13139 3451
rect 13081 3411 13139 3417
rect 17586 3380 17592 3392
rect 13004 3352 17592 3380
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 9030 3176 9036 3188
rect 5868 3148 9036 3176
rect 5868 3136 5874 3148
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 10413 3179 10471 3185
rect 10413 3145 10425 3179
rect 10459 3176 10471 3179
rect 10870 3176 10876 3188
rect 10459 3148 10876 3176
rect 10459 3145 10471 3148
rect 10413 3139 10471 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 13170 3176 13176 3188
rect 11020 3148 13176 3176
rect 11020 3136 11026 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 13354 3176 13360 3188
rect 13315 3148 13360 3176
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14424 3148 15424 3176
rect 14424 3136 14430 3148
rect 7466 3068 7472 3120
rect 7524 3108 7530 3120
rect 10226 3108 10232 3120
rect 7524 3080 10232 3108
rect 7524 3068 7530 3080
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 10704 3080 10916 3108
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10704 3040 10732 3080
rect 10376 3012 10732 3040
rect 10888 3040 10916 3080
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10888 3012 10977 3040
rect 10376 3000 10382 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 10965 3003 11023 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14366 3040 14372 3052
rect 14327 3012 14372 3040
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 15396 3040 15424 3148
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 16206 3176 16212 3188
rect 15620 3148 16212 3176
rect 15620 3136 15626 3148
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 16485 3179 16543 3185
rect 16485 3145 16497 3179
rect 16531 3176 16543 3179
rect 16942 3176 16948 3188
rect 16531 3148 16948 3176
rect 16531 3145 16543 3148
rect 16485 3139 16543 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 18012 3148 18061 3176
rect 18012 3136 18018 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 15749 3111 15807 3117
rect 15749 3077 15761 3111
rect 15795 3108 15807 3111
rect 16114 3108 16120 3120
rect 15795 3080 16120 3108
rect 15795 3077 15807 3080
rect 15749 3071 15807 3077
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 20254 3108 20260 3120
rect 19659 3080 20260 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 20254 3068 20260 3080
rect 20312 3068 20318 3120
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 15396 3012 16037 3040
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 16025 3003 16083 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 10594 2972 10600 2984
rect 7524 2944 10600 2972
rect 7524 2932 7530 2944
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10870 2972 10876 2984
rect 10831 2944 10876 2972
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 11606 2972 11612 2984
rect 11567 2944 11612 2972
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12483 2944 12940 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 8570 2864 8576 2916
rect 8628 2904 8634 2916
rect 8628 2876 10916 2904
rect 8628 2864 8634 2876
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 10781 2839 10839 2845
rect 10781 2836 10793 2839
rect 4764 2808 10793 2836
rect 4764 2796 4770 2808
rect 10781 2805 10793 2808
rect 10827 2805 10839 2839
rect 10888 2836 10916 2876
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 11388 2876 11897 2904
rect 11388 2864 11394 2876
rect 11885 2873 11897 2876
rect 11931 2873 11943 2907
rect 11885 2867 11943 2873
rect 11974 2864 11980 2916
rect 12032 2904 12038 2916
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 12032 2876 12725 2904
rect 12032 2864 12038 2876
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 12912 2904 12940 2944
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13044 2944 13737 2972
rect 13044 2932 13050 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 15470 2972 15476 2984
rect 13725 2935 13783 2941
rect 13823 2944 15476 2972
rect 13823 2904 13851 2944
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17644 2944 18429 2972
rect 17644 2932 17650 2944
rect 18417 2941 18429 2944
rect 18463 2972 18475 2975
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 18463 2944 18889 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 19610 2972 19616 2984
rect 19475 2944 19616 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20530 2972 20536 2984
rect 20491 2944 20536 2972
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 12912 2876 13851 2904
rect 12713 2867 12771 2873
rect 14550 2864 14556 2916
rect 14608 2913 14614 2916
rect 14608 2907 14672 2913
rect 14608 2873 14626 2907
rect 14660 2873 14672 2907
rect 14608 2867 14672 2873
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 17497 2907 17555 2913
rect 17497 2904 17509 2907
rect 16899 2876 17509 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 17497 2873 17509 2876
rect 17543 2873 17555 2907
rect 17497 2867 17555 2873
rect 18509 2907 18567 2913
rect 18509 2873 18521 2907
rect 18555 2904 18567 2907
rect 18690 2904 18696 2916
rect 18555 2876 18696 2904
rect 18555 2873 18567 2876
rect 18509 2867 18567 2873
rect 14608 2864 14614 2867
rect 18690 2864 18696 2876
rect 18748 2864 18754 2916
rect 21358 2904 21364 2916
rect 20180 2876 21364 2904
rect 12526 2836 12532 2848
rect 10888 2808 12532 2836
rect 10781 2799 10839 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 13817 2839 13875 2845
rect 13817 2805 13829 2839
rect 13863 2836 13875 2839
rect 16758 2836 16764 2848
rect 13863 2808 16764 2836
rect 13863 2805 13875 2808
rect 13817 2799 13875 2805
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 20180 2845 20208 2876
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 20165 2839 20223 2845
rect 17000 2808 17045 2836
rect 17000 2796 17006 2808
rect 20165 2805 20177 2839
rect 20211 2805 20223 2839
rect 20165 2799 20223 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 21910 2836 21916 2848
rect 20763 2808 21916 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 12526 2592 12532 2644
rect 12584 2632 12590 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 12584 2604 14473 2632
rect 12584 2592 12590 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 15565 2635 15623 2641
rect 15565 2601 15577 2635
rect 15611 2632 15623 2635
rect 16942 2632 16948 2644
rect 15611 2604 16948 2632
rect 15611 2601 15623 2604
rect 15565 2595 15623 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 13814 2564 13820 2576
rect 12912 2536 13656 2564
rect 13775 2536 13820 2564
rect 11330 2496 11336 2508
rect 11291 2468 11336 2496
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 11885 2499 11943 2505
rect 11885 2465 11897 2499
rect 11931 2496 11943 2499
rect 11974 2496 11980 2508
rect 11931 2468 11980 2496
rect 11931 2465 11943 2468
rect 11885 2459 11943 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 12805 2499 12863 2505
rect 12805 2496 12817 2499
rect 12676 2468 12817 2496
rect 12676 2456 12682 2468
rect 12805 2465 12817 2468
rect 12851 2465 12863 2499
rect 12805 2459 12863 2465
rect 1394 2388 1400 2440
rect 1452 2428 1458 2440
rect 12912 2428 12940 2536
rect 13446 2456 13452 2508
rect 13504 2496 13510 2508
rect 13541 2499 13599 2505
rect 13541 2496 13553 2499
rect 13504 2468 13553 2496
rect 13504 2456 13510 2468
rect 13541 2465 13553 2468
rect 13587 2465 13599 2499
rect 13628 2496 13656 2536
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 13924 2536 15945 2564
rect 13924 2496 13952 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 16758 2524 16764 2576
rect 16816 2564 16822 2576
rect 17494 2564 17500 2576
rect 16816 2536 17500 2564
rect 16816 2524 16822 2536
rect 17494 2524 17500 2536
rect 17552 2564 17558 2576
rect 18598 2564 18604 2576
rect 17552 2536 18604 2564
rect 17552 2524 17558 2536
rect 18598 2524 18604 2536
rect 18656 2524 18662 2576
rect 13628 2468 13952 2496
rect 14277 2499 14335 2505
rect 13541 2459 13599 2465
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 15562 2496 15568 2508
rect 14875 2468 15568 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 1452 2400 12940 2428
rect 13081 2431 13139 2437
rect 1452 2388 1458 2400
rect 13081 2397 13093 2431
rect 13127 2428 13139 2431
rect 14292 2428 14320 2459
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 16574 2496 16580 2508
rect 16535 2468 16580 2496
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 17313 2499 17371 2505
rect 17313 2465 17325 2499
rect 17359 2496 17371 2499
rect 17770 2496 17776 2508
rect 17359 2468 17776 2496
rect 17359 2465 17371 2468
rect 17313 2459 17371 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 18414 2496 18420 2508
rect 18375 2468 18420 2496
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 18969 2499 19027 2505
rect 18969 2465 18981 2499
rect 19015 2465 19027 2499
rect 19518 2496 19524 2508
rect 19479 2468 19524 2496
rect 18969 2459 19027 2465
rect 13127 2400 14320 2428
rect 13127 2397 13139 2400
rect 13081 2391 13139 2397
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15712 2400 16037 2428
rect 15712 2388 15718 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16172 2400 16217 2428
rect 16172 2388 16178 2400
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 18984 2428 19012 2459
rect 19518 2456 19524 2468
rect 19576 2456 19582 2508
rect 20346 2496 20352 2508
rect 20307 2468 20352 2496
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 16356 2400 19012 2428
rect 16356 2388 16362 2400
rect 11517 2363 11575 2369
rect 11517 2329 11529 2363
rect 11563 2360 11575 2363
rect 11563 2332 13124 2360
rect 11563 2329 11575 2332
rect 11517 2323 11575 2329
rect 13096 2304 13124 2332
rect 13630 2320 13636 2372
rect 13688 2360 13694 2372
rect 15013 2363 15071 2369
rect 15013 2360 15025 2363
rect 13688 2332 15025 2360
rect 13688 2320 13694 2332
rect 15013 2329 15025 2332
rect 15059 2329 15071 2363
rect 15013 2323 15071 2329
rect 18690 2320 18696 2372
rect 18748 2360 18754 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 18748 2332 19717 2360
rect 18748 2320 18754 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12069 2295 12127 2301
rect 12069 2292 12081 2295
rect 12032 2264 12081 2292
rect 12032 2252 12038 2264
rect 12069 2261 12081 2264
rect 12115 2261 12127 2295
rect 12069 2255 12127 2261
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 16761 2295 16819 2301
rect 16761 2261 16773 2295
rect 16807 2292 16819 2295
rect 16942 2292 16948 2304
rect 16807 2264 16948 2292
rect 16807 2261 16819 2264
rect 16761 2255 16819 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17494 2292 17500 2304
rect 17455 2264 17500 2292
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 19058 2292 19064 2304
rect 18647 2264 19064 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 19153 2295 19211 2301
rect 19153 2261 19165 2295
rect 19199 2292 19211 2295
rect 19610 2292 19616 2304
rect 19199 2264 19616 2292
rect 19199 2261 19211 2264
rect 19153 2255 19211 2261
rect 19610 2252 19616 2264
rect 19668 2252 19674 2304
rect 20533 2295 20591 2301
rect 20533 2261 20545 2295
rect 20579 2292 20591 2295
rect 20806 2292 20812 2304
rect 20579 2264 20812 2292
rect 20579 2261 20591 2264
rect 20533 2255 20591 2261
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 9674 1368 9680 1420
rect 9732 1408 9738 1420
rect 10962 1408 10968 1420
rect 9732 1380 10968 1408
rect 9732 1368 9738 1380
rect 10962 1368 10968 1380
rect 11020 1368 11026 1420
rect 10226 1096 10232 1148
rect 10284 1136 10290 1148
rect 12066 1136 12072 1148
rect 10284 1108 12072 1136
rect 10284 1096 10290 1108
rect 12066 1096 12072 1108
rect 12124 1096 12130 1148
<< via1 >>
rect 7472 20272 7524 20324
rect 11888 20272 11940 20324
rect 8760 20204 8812 20256
rect 22468 20204 22520 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 10600 20000 10652 20052
rect 11336 20000 11388 20052
rect 13084 20000 13136 20052
rect 14188 20000 14240 20052
rect 15844 20000 15896 20052
rect 16580 20000 16632 20052
rect 17500 20000 17552 20052
rect 18512 20043 18564 20052
rect 18512 20009 18521 20043
rect 18521 20009 18555 20043
rect 18555 20009 18564 20043
rect 18512 20000 18564 20009
rect 18604 20000 18656 20052
rect 19340 20000 19392 20052
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20628 20000 20680 20052
rect 17316 19932 17368 19984
rect 10232 19864 10284 19916
rect 11888 19864 11940 19916
rect 12808 19907 12860 19916
rect 12808 19873 12817 19907
rect 12817 19873 12851 19907
rect 12851 19873 12860 19907
rect 12808 19864 12860 19873
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 14372 19907 14424 19916
rect 14372 19873 14381 19907
rect 14381 19873 14415 19907
rect 14415 19873 14424 19907
rect 14372 19864 14424 19873
rect 15568 19907 15620 19916
rect 15568 19873 15577 19907
rect 15577 19873 15611 19907
rect 15611 19873 15620 19907
rect 15568 19864 15620 19873
rect 15752 19864 15804 19916
rect 16396 19864 16448 19916
rect 16764 19864 16816 19916
rect 18604 19864 18656 19916
rect 18880 19907 18932 19916
rect 18880 19873 18889 19907
rect 18889 19873 18923 19907
rect 18923 19873 18932 19907
rect 18880 19864 18932 19873
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 19984 19907 20036 19916
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 20168 19864 20220 19916
rect 10508 19796 10560 19848
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 19248 19796 19300 19848
rect 21364 19796 21416 19848
rect 9772 19728 9824 19780
rect 15292 19728 15344 19780
rect 18144 19728 18196 19780
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 12256 19660 12308 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 7748 19252 7800 19304
rect 10232 19456 10284 19508
rect 15936 19456 15988 19508
rect 1952 19184 2004 19236
rect 2964 19184 3016 19236
rect 3056 19184 3108 19236
rect 10140 19252 10192 19304
rect 16672 19320 16724 19372
rect 10324 19252 10376 19304
rect 12164 19252 12216 19304
rect 12532 19252 12584 19304
rect 14188 19252 14240 19304
rect 14280 19252 14332 19304
rect 9220 19184 9272 19236
rect 10416 19184 10468 19236
rect 10692 19184 10744 19236
rect 10876 19184 10928 19236
rect 1400 19116 1452 19168
rect 8484 19116 8536 19168
rect 8576 19116 8628 19168
rect 10784 19116 10836 19168
rect 11612 19159 11664 19168
rect 11612 19125 11621 19159
rect 11621 19125 11655 19159
rect 11655 19125 11664 19159
rect 11612 19116 11664 19125
rect 11980 19184 12032 19236
rect 13636 19184 13688 19236
rect 14464 19252 14516 19304
rect 15568 19252 15620 19304
rect 16856 19252 16908 19304
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 18420 19252 18472 19304
rect 12072 19116 12124 19168
rect 12348 19116 12400 19168
rect 12532 19116 12584 19168
rect 12992 19116 13044 19168
rect 13544 19116 13596 19168
rect 17224 19184 17276 19236
rect 18604 19184 18656 19236
rect 18972 19184 19024 19236
rect 19800 19184 19852 19236
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 19064 19116 19116 19168
rect 19340 19116 19392 19168
rect 21916 19116 21968 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 2964 18912 3016 18964
rect 9220 18955 9272 18964
rect 9220 18921 9229 18955
rect 9229 18921 9263 18955
rect 9263 18921 9272 18955
rect 9220 18912 9272 18921
rect 11796 18912 11848 18964
rect 11980 18955 12032 18964
rect 11980 18921 11989 18955
rect 11989 18921 12023 18955
rect 12023 18921 12032 18955
rect 11980 18912 12032 18921
rect 12164 18912 12216 18964
rect 14280 18912 14332 18964
rect 14556 18912 14608 18964
rect 15936 18912 15988 18964
rect 16488 18912 16540 18964
rect 16672 18955 16724 18964
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 16948 18912 17000 18964
rect 17960 18912 18012 18964
rect 20904 18912 20956 18964
rect 9772 18844 9824 18896
rect 10692 18844 10744 18896
rect 11612 18844 11664 18896
rect 12992 18887 13044 18896
rect 12992 18853 13026 18887
rect 13026 18853 13044 18887
rect 12992 18844 13044 18853
rect 13084 18844 13136 18896
rect 19984 18887 20036 18896
rect 7748 18776 7800 18828
rect 8852 18776 8904 18828
rect 9956 18776 10008 18828
rect 12532 18776 12584 18828
rect 14280 18776 14332 18828
rect 15384 18776 15436 18828
rect 15844 18776 15896 18828
rect 10508 18708 10560 18760
rect 13912 18708 13964 18760
rect 15108 18708 15160 18760
rect 16580 18776 16632 18828
rect 17316 18776 17368 18828
rect 19708 18819 19760 18828
rect 18788 18751 18840 18760
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 18788 18708 18840 18717
rect 19708 18785 19717 18819
rect 19717 18785 19751 18819
rect 19751 18785 19760 18819
rect 19708 18776 19760 18785
rect 19984 18853 19993 18887
rect 19993 18853 20027 18887
rect 20027 18853 20036 18887
rect 19984 18844 20036 18853
rect 20260 18776 20312 18828
rect 20720 18708 20772 18760
rect 296 18640 348 18692
rect 7656 18640 7708 18692
rect 8208 18572 8260 18624
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 14188 18572 14240 18624
rect 15016 18572 15068 18624
rect 16304 18640 16356 18692
rect 19616 18640 19668 18692
rect 16028 18572 16080 18624
rect 16856 18572 16908 18624
rect 17776 18572 17828 18624
rect 18512 18572 18564 18624
rect 19248 18572 19300 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 2504 18368 2556 18420
rect 10508 18368 10560 18420
rect 12440 18368 12492 18420
rect 13084 18368 13136 18420
rect 13176 18368 13228 18420
rect 15384 18411 15436 18420
rect 4160 18300 4212 18352
rect 4712 18232 4764 18284
rect 6184 18232 6236 18284
rect 3608 18164 3660 18216
rect 8576 18232 8628 18284
rect 10140 18300 10192 18352
rect 10232 18300 10284 18352
rect 14004 18300 14056 18352
rect 15384 18377 15393 18411
rect 15393 18377 15427 18411
rect 15427 18377 15436 18411
rect 15384 18368 15436 18377
rect 16304 18368 16356 18420
rect 18788 18368 18840 18420
rect 19156 18368 19208 18420
rect 15844 18300 15896 18352
rect 9036 18232 9088 18284
rect 9220 18232 9272 18284
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 10784 18232 10836 18284
rect 6368 18164 6420 18216
rect 8668 18164 8720 18216
rect 10048 18164 10100 18216
rect 11060 18207 11112 18216
rect 11060 18173 11069 18207
rect 11069 18173 11103 18207
rect 11103 18173 11112 18207
rect 11060 18164 11112 18173
rect 11980 18164 12032 18216
rect 13176 18232 13228 18284
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 15108 18232 15160 18284
rect 18604 18275 18656 18284
rect 9128 18096 9180 18148
rect 9680 18096 9732 18148
rect 13912 18164 13964 18216
rect 14096 18164 14148 18216
rect 15660 18164 15712 18216
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 16856 18164 16908 18216
rect 18512 18164 18564 18216
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 5816 18028 5868 18080
rect 7472 18028 7524 18080
rect 7656 18028 7708 18080
rect 9864 18028 9916 18080
rect 10324 18028 10376 18080
rect 13084 18028 13136 18080
rect 13268 18028 13320 18080
rect 14188 18028 14240 18080
rect 16672 18096 16724 18148
rect 20076 18164 20128 18216
rect 20536 18096 20588 18148
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 7748 17824 7800 17876
rect 8852 17867 8904 17876
rect 8852 17833 8861 17867
rect 8861 17833 8895 17867
rect 8895 17833 8904 17867
rect 8852 17824 8904 17833
rect 9496 17824 9548 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10140 17824 10192 17833
rect 9128 17756 9180 17808
rect 13268 17824 13320 17876
rect 13636 17824 13688 17876
rect 15476 17824 15528 17876
rect 16120 17824 16172 17876
rect 18512 17824 18564 17876
rect 18972 17824 19024 17876
rect 20904 17867 20956 17876
rect 20904 17833 20913 17867
rect 20913 17833 20947 17867
rect 20947 17833 20956 17867
rect 20904 17824 20956 17833
rect 13176 17756 13228 17808
rect 8300 17688 8352 17740
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 10324 17688 10376 17740
rect 12624 17688 12676 17740
rect 14004 17731 14056 17740
rect 10416 17620 10468 17672
rect 12072 17663 12124 17672
rect 12072 17629 12081 17663
rect 12081 17629 12115 17663
rect 12115 17629 12124 17663
rect 12072 17620 12124 17629
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 12900 17620 12952 17672
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 14004 17697 14013 17731
rect 14013 17697 14047 17731
rect 14047 17697 14056 17731
rect 14004 17688 14056 17697
rect 16948 17756 17000 17808
rect 17224 17756 17276 17808
rect 16856 17688 16908 17740
rect 18788 17688 18840 17740
rect 19156 17731 19208 17740
rect 19156 17697 19165 17731
rect 19165 17697 19199 17731
rect 19199 17697 19208 17731
rect 19156 17688 19208 17697
rect 13544 17620 13596 17629
rect 15476 17620 15528 17672
rect 15660 17620 15712 17672
rect 16304 17620 16356 17672
rect 15200 17552 15252 17604
rect 18604 17552 18656 17604
rect 18788 17552 18840 17604
rect 848 17484 900 17536
rect 8484 17484 8536 17536
rect 11152 17484 11204 17536
rect 11704 17484 11756 17536
rect 12348 17484 12400 17536
rect 16764 17484 16816 17536
rect 16856 17484 16908 17536
rect 17132 17484 17184 17536
rect 17408 17484 17460 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 8300 17280 8352 17332
rect 9036 17280 9088 17332
rect 8484 17212 8536 17264
rect 8760 17144 8812 17196
rect 9496 17144 9548 17196
rect 7748 17076 7800 17128
rect 8208 17076 8260 17128
rect 7656 17008 7708 17060
rect 13452 17280 13504 17332
rect 10508 17144 10560 17196
rect 11704 17144 11756 17196
rect 11612 17076 11664 17128
rect 12900 17212 12952 17264
rect 12992 17212 13044 17264
rect 15660 17280 15712 17332
rect 16212 17280 16264 17332
rect 16948 17280 17000 17332
rect 19340 17280 19392 17332
rect 12256 17144 12308 17196
rect 13544 17144 13596 17196
rect 15292 17212 15344 17264
rect 16764 17212 16816 17264
rect 18052 17212 18104 17264
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 16488 17144 16540 17196
rect 12716 17076 12768 17128
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 15476 17076 15528 17128
rect 17132 17008 17184 17060
rect 19616 17144 19668 17196
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 17868 17076 17920 17128
rect 18604 17076 18656 17128
rect 19892 17076 19944 17128
rect 19524 17008 19576 17060
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9680 16983 9732 16992
rect 9128 16940 9180 16949
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 9864 16940 9916 16992
rect 10508 16940 10560 16992
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 13268 16940 13320 16992
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 14188 16940 14240 16992
rect 15476 16940 15528 16992
rect 16304 16940 16356 16992
rect 17960 16940 18012 16992
rect 19340 16940 19392 16992
rect 19984 16983 20036 16992
rect 19984 16949 19993 16983
rect 19993 16949 20027 16983
rect 20027 16949 20036 16983
rect 19984 16940 20036 16949
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 6920 16736 6972 16788
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 8208 16779 8260 16788
rect 7472 16736 7524 16745
rect 8208 16745 8217 16779
rect 8217 16745 8251 16779
rect 8251 16745 8260 16779
rect 8208 16736 8260 16745
rect 9036 16736 9088 16788
rect 10876 16736 10928 16788
rect 10968 16736 11020 16788
rect 12072 16736 12124 16788
rect 13268 16736 13320 16788
rect 14096 16736 14148 16788
rect 16948 16736 17000 16788
rect 17132 16779 17184 16788
rect 17132 16745 17141 16779
rect 17141 16745 17175 16779
rect 17175 16745 17184 16779
rect 17132 16736 17184 16745
rect 18880 16736 18932 16788
rect 19892 16736 19944 16788
rect 9220 16600 9272 16652
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 12440 16668 12492 16720
rect 20260 16668 20312 16720
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 8208 16532 8260 16584
rect 8760 16575 8812 16584
rect 8760 16541 8769 16575
rect 8769 16541 8803 16575
rect 8803 16541 8812 16575
rect 8760 16532 8812 16541
rect 11704 16600 11756 16652
rect 11888 16643 11940 16652
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 12900 16600 12952 16652
rect 13636 16600 13688 16652
rect 15292 16600 15344 16652
rect 15568 16600 15620 16652
rect 7748 16464 7800 16516
rect 9404 16464 9456 16516
rect 13268 16439 13320 16448
rect 13268 16405 13277 16439
rect 13277 16405 13311 16439
rect 13311 16405 13320 16439
rect 13268 16396 13320 16405
rect 13360 16396 13412 16448
rect 15200 16532 15252 16584
rect 15752 16532 15804 16584
rect 16028 16600 16080 16652
rect 17592 16600 17644 16652
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 18512 16600 18564 16652
rect 19432 16600 19484 16652
rect 16212 16575 16264 16584
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 17316 16575 17368 16584
rect 15292 16464 15344 16516
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 17684 16532 17736 16584
rect 19340 16532 19392 16584
rect 16488 16464 16540 16516
rect 15016 16396 15068 16448
rect 15752 16439 15804 16448
rect 15752 16405 15761 16439
rect 15761 16405 15795 16439
rect 15795 16405 15804 16439
rect 15752 16396 15804 16405
rect 15844 16396 15896 16448
rect 18604 16439 18656 16448
rect 18604 16405 18613 16439
rect 18613 16405 18647 16439
rect 18647 16405 18656 16439
rect 18604 16396 18656 16405
rect 20720 16396 20772 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 8208 16235 8260 16244
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 6920 15988 6972 16040
rect 7656 15988 7708 16040
rect 9680 16192 9732 16244
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 10876 16056 10928 16108
rect 12256 16192 12308 16244
rect 12624 16192 12676 16244
rect 14280 16192 14332 16244
rect 12164 16124 12216 16176
rect 12716 16124 12768 16176
rect 13636 16124 13688 16176
rect 15016 16124 15068 16176
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 13268 16056 13320 16108
rect 13728 16056 13780 16108
rect 14004 16099 14056 16108
rect 14004 16065 14013 16099
rect 14013 16065 14047 16099
rect 14047 16065 14056 16099
rect 14004 16056 14056 16065
rect 15752 16056 15804 16108
rect 20720 16192 20772 16244
rect 17316 16099 17368 16108
rect 17316 16065 17325 16099
rect 17325 16065 17359 16099
rect 17359 16065 17368 16099
rect 17316 16056 17368 16065
rect 19892 16056 19944 16108
rect 8852 15920 8904 15972
rect 10968 15920 11020 15972
rect 12164 15920 12216 15972
rect 12532 15988 12584 16040
rect 13360 15988 13412 16040
rect 15016 15920 15068 15972
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 12256 15852 12308 15904
rect 12992 15852 13044 15904
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 16948 15988 17000 16040
rect 17684 15988 17736 16040
rect 17960 15988 18012 16040
rect 19340 15920 19392 15972
rect 20168 15963 20220 15972
rect 20168 15929 20177 15963
rect 20177 15929 20211 15963
rect 20211 15929 20220 15963
rect 20168 15920 20220 15929
rect 20904 15920 20956 15972
rect 17960 15852 18012 15904
rect 18788 15852 18840 15904
rect 19800 15895 19852 15904
rect 19800 15861 19809 15895
rect 19809 15861 19843 15895
rect 19843 15861 19852 15895
rect 19800 15852 19852 15861
rect 20996 15895 21048 15904
rect 20996 15861 21005 15895
rect 21005 15861 21039 15895
rect 21039 15861 21048 15895
rect 20996 15852 21048 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 11336 15648 11388 15700
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 13912 15648 13964 15700
rect 15200 15648 15252 15700
rect 15660 15691 15712 15700
rect 15660 15657 15669 15691
rect 15669 15657 15703 15691
rect 15703 15657 15712 15691
rect 15660 15648 15712 15657
rect 17316 15648 17368 15700
rect 19432 15648 19484 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 6920 15512 6972 15564
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 9772 15512 9824 15564
rect 10140 15512 10192 15564
rect 10784 15512 10836 15564
rect 11888 15580 11940 15632
rect 15844 15580 15896 15632
rect 9864 15444 9916 15496
rect 10876 15487 10928 15496
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 11796 15555 11848 15564
rect 11796 15521 11830 15555
rect 11830 15521 11848 15555
rect 11796 15512 11848 15521
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 15016 15444 15068 15496
rect 15384 15512 15436 15564
rect 15660 15444 15712 15496
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 16120 15444 16172 15496
rect 17960 15580 18012 15632
rect 18788 15623 18840 15632
rect 17500 15512 17552 15564
rect 18788 15589 18822 15623
rect 18822 15589 18840 15623
rect 18788 15580 18840 15589
rect 20260 15555 20312 15564
rect 17776 15444 17828 15496
rect 20260 15521 20269 15555
rect 20269 15521 20303 15555
rect 20303 15521 20312 15555
rect 20260 15512 20312 15521
rect 20904 15444 20956 15496
rect 17408 15308 17460 15360
rect 17592 15308 17644 15360
rect 20168 15308 20220 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 8852 15036 8904 15088
rect 9036 15079 9088 15088
rect 9036 15045 9045 15079
rect 9045 15045 9079 15079
rect 9079 15045 9088 15079
rect 9036 15036 9088 15045
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 7564 14968 7616 15020
rect 9864 15104 9916 15156
rect 10876 15104 10928 15156
rect 9864 15011 9916 15020
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 10692 14968 10744 15020
rect 10968 15011 11020 15020
rect 10968 14977 10977 15011
rect 10977 14977 11011 15011
rect 11011 14977 11020 15011
rect 10968 14968 11020 14977
rect 11796 14968 11848 15020
rect 12348 14968 12400 15020
rect 5540 14900 5592 14952
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6092 14900 6144 14909
rect 6828 14832 6880 14884
rect 11520 14900 11572 14952
rect 12716 14900 12768 14952
rect 9772 14832 9824 14884
rect 11060 14832 11112 14884
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 10232 14764 10284 14816
rect 13728 14832 13780 14884
rect 14004 14968 14056 15020
rect 15292 14968 15344 15020
rect 15476 14968 15528 15020
rect 15384 14900 15436 14952
rect 17868 15104 17920 15156
rect 20076 15104 20128 15156
rect 20812 15147 20864 15156
rect 20812 15113 20821 15147
rect 20821 15113 20855 15147
rect 20855 15113 20864 15147
rect 20812 15104 20864 15113
rect 17040 15036 17092 15088
rect 19708 15036 19760 15088
rect 19892 15036 19944 15088
rect 20352 15036 20404 15088
rect 16396 14968 16448 15020
rect 16856 14968 16908 15020
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 18788 14968 18840 15020
rect 19800 14968 19852 15020
rect 20444 14968 20496 15020
rect 16488 14900 16540 14952
rect 17684 14900 17736 14952
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 20536 14900 20588 14952
rect 16396 14832 16448 14884
rect 18604 14832 18656 14884
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 13084 14807 13136 14816
rect 11796 14764 11848 14773
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 14556 14764 14608 14816
rect 15292 14764 15344 14816
rect 16304 14807 16356 14816
rect 16304 14773 16313 14807
rect 16313 14773 16347 14807
rect 16347 14773 16356 14807
rect 16304 14764 16356 14773
rect 16672 14807 16724 14816
rect 16672 14773 16681 14807
rect 16681 14773 16715 14807
rect 16715 14773 16724 14807
rect 16672 14764 16724 14773
rect 17132 14807 17184 14816
rect 17132 14773 17141 14807
rect 17141 14773 17175 14807
rect 17175 14773 17184 14807
rect 17132 14764 17184 14773
rect 18880 14764 18932 14816
rect 19616 14764 19668 14816
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 7564 14492 7616 14544
rect 9312 14560 9364 14612
rect 9496 14560 9548 14612
rect 12348 14560 12400 14612
rect 13084 14560 13136 14612
rect 13728 14603 13780 14612
rect 13728 14569 13737 14603
rect 13737 14569 13771 14603
rect 13771 14569 13780 14603
rect 13728 14560 13780 14569
rect 14004 14560 14056 14612
rect 16120 14560 16172 14612
rect 17500 14603 17552 14612
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 17592 14560 17644 14612
rect 18512 14560 18564 14612
rect 20444 14603 20496 14612
rect 20444 14569 20453 14603
rect 20453 14569 20487 14603
rect 20487 14569 20496 14603
rect 20444 14560 20496 14569
rect 9680 14492 9732 14544
rect 13268 14492 13320 14544
rect 14372 14492 14424 14544
rect 15200 14492 15252 14544
rect 6828 14467 6880 14476
rect 6828 14433 6837 14467
rect 6837 14433 6871 14467
rect 6871 14433 6880 14467
rect 6828 14424 6880 14433
rect 8484 14424 8536 14476
rect 9772 14424 9824 14476
rect 11520 14467 11572 14476
rect 9036 14399 9088 14408
rect 9036 14365 9045 14399
rect 9045 14365 9079 14399
rect 9079 14365 9088 14399
rect 9036 14356 9088 14365
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 11888 14467 11940 14476
rect 11888 14433 11922 14467
rect 11922 14433 11940 14467
rect 17224 14492 17276 14544
rect 11888 14424 11940 14433
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 16764 14424 16816 14476
rect 17776 14424 17828 14476
rect 17960 14424 18012 14476
rect 19524 14492 19576 14544
rect 20168 14492 20220 14544
rect 12900 14356 12952 14408
rect 15200 14356 15252 14408
rect 15752 14356 15804 14408
rect 17868 14356 17920 14408
rect 19156 14424 19208 14476
rect 20352 14424 20404 14476
rect 20168 14356 20220 14408
rect 17408 14288 17460 14340
rect 18512 14288 18564 14340
rect 9864 14220 9916 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 13084 14220 13136 14272
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 11704 14016 11756 14068
rect 13452 14016 13504 14068
rect 14556 14016 14608 14068
rect 11796 13948 11848 14000
rect 8576 13880 8628 13932
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 9864 13880 9916 13932
rect 10876 13880 10928 13932
rect 10968 13880 11020 13932
rect 11888 13923 11940 13932
rect 11336 13812 11388 13864
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 13820 13880 13872 13932
rect 15292 14016 15344 14068
rect 16120 14016 16172 14068
rect 16580 14016 16632 14068
rect 17224 14016 17276 14068
rect 17960 14016 18012 14068
rect 19984 14016 20036 14068
rect 20628 14016 20680 14068
rect 15660 13948 15712 14000
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 12624 13812 12676 13864
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 16304 13855 16356 13864
rect 16304 13821 16313 13855
rect 16313 13821 16347 13855
rect 16347 13821 16356 13855
rect 16304 13812 16356 13821
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 10692 13676 10744 13728
rect 11796 13676 11848 13728
rect 12256 13676 12308 13728
rect 12440 13676 12492 13728
rect 12532 13676 12584 13728
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 14004 13719 14056 13728
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 15660 13744 15712 13796
rect 18788 13812 18840 13864
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 18604 13744 18656 13796
rect 19340 13787 19392 13796
rect 19340 13753 19349 13787
rect 19349 13753 19383 13787
rect 19383 13753 19392 13787
rect 19340 13744 19392 13753
rect 19800 13744 19852 13796
rect 20076 13744 20128 13796
rect 15936 13719 15988 13728
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 17684 13676 17736 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 9680 13472 9732 13524
rect 11336 13515 11388 13524
rect 11336 13481 11345 13515
rect 11345 13481 11379 13515
rect 11379 13481 11388 13515
rect 11336 13472 11388 13481
rect 10232 13404 10284 13456
rect 12532 13472 12584 13524
rect 12716 13515 12768 13524
rect 12716 13481 12725 13515
rect 12725 13481 12759 13515
rect 12759 13481 12768 13515
rect 12716 13472 12768 13481
rect 14004 13515 14056 13524
rect 14004 13481 14013 13515
rect 14013 13481 14047 13515
rect 14047 13481 14056 13515
rect 14004 13472 14056 13481
rect 12072 13404 12124 13456
rect 16120 13472 16172 13524
rect 16396 13472 16448 13524
rect 16672 13472 16724 13524
rect 17776 13472 17828 13524
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 19064 13472 19116 13524
rect 19892 13472 19944 13524
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 11060 13336 11112 13388
rect 12716 13336 12768 13388
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 19340 13404 19392 13456
rect 14280 13200 14332 13252
rect 10876 13132 10928 13184
rect 12072 13132 12124 13184
rect 14648 13132 14700 13184
rect 15476 13336 15528 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 18144 13379 18196 13388
rect 18144 13345 18153 13379
rect 18153 13345 18187 13379
rect 18187 13345 18196 13379
rect 18144 13336 18196 13345
rect 18512 13336 18564 13388
rect 19708 13379 19760 13388
rect 19708 13345 19717 13379
rect 19717 13345 19751 13379
rect 19751 13345 19760 13379
rect 19708 13336 19760 13345
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 17500 13268 17552 13320
rect 18604 13268 18656 13320
rect 19064 13268 19116 13320
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 15200 13200 15252 13252
rect 17868 13200 17920 13252
rect 16580 13132 16632 13184
rect 18788 13132 18840 13184
rect 20444 13132 20496 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 8944 12928 8996 12980
rect 11152 12928 11204 12980
rect 12716 12928 12768 12980
rect 15936 12928 15988 12980
rect 17132 12928 17184 12980
rect 10140 12792 10192 12844
rect 9680 12724 9732 12776
rect 10232 12656 10284 12708
rect 9588 12588 9640 12640
rect 15200 12860 15252 12912
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 14648 12792 14700 12844
rect 12808 12724 12860 12776
rect 12992 12724 13044 12776
rect 16304 12724 16356 12776
rect 17960 12724 18012 12776
rect 18972 12928 19024 12980
rect 19064 12928 19116 12980
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 18604 12724 18656 12776
rect 20444 12767 20496 12776
rect 13820 12699 13872 12708
rect 13820 12665 13854 12699
rect 13854 12665 13872 12699
rect 13820 12656 13872 12665
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 12440 12588 12492 12640
rect 12900 12631 12952 12640
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 13912 12588 13964 12640
rect 14372 12588 14424 12640
rect 16028 12656 16080 12708
rect 17224 12699 17276 12708
rect 17224 12665 17233 12699
rect 17233 12665 17267 12699
rect 17267 12665 17276 12699
rect 17224 12656 17276 12665
rect 15844 12588 15896 12640
rect 17408 12588 17460 12640
rect 18604 12588 18656 12640
rect 20444 12733 20453 12767
rect 20453 12733 20487 12767
rect 20487 12733 20496 12767
rect 20444 12724 20496 12733
rect 19984 12656 20036 12708
rect 19156 12588 19208 12640
rect 19340 12588 19392 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 10232 12384 10284 12436
rect 10876 12384 10928 12436
rect 9588 12316 9640 12368
rect 13084 12384 13136 12436
rect 19708 12384 19760 12436
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 15936 12316 15988 12368
rect 16396 12316 16448 12368
rect 16856 12316 16908 12368
rect 9680 12248 9732 12300
rect 10600 12248 10652 12300
rect 11060 12248 11112 12300
rect 12072 12248 12124 12300
rect 12992 12248 13044 12300
rect 14556 12248 14608 12300
rect 17868 12248 17920 12300
rect 18880 12291 18932 12300
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 10968 12112 11020 12164
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9680 12044 9732 12096
rect 10876 12044 10928 12096
rect 15476 12180 15528 12232
rect 14372 12112 14424 12164
rect 14648 12044 14700 12096
rect 15200 12044 15252 12096
rect 17408 12180 17460 12232
rect 18880 12257 18914 12291
rect 18914 12257 18932 12291
rect 18880 12248 18932 12257
rect 19156 12248 19208 12300
rect 18604 12223 18656 12232
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 18604 12180 18656 12189
rect 16304 12044 16356 12096
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 19248 12044 19300 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 12440 11840 12492 11892
rect 12900 11840 12952 11892
rect 10692 11772 10744 11824
rect 13728 11840 13780 11892
rect 14004 11840 14056 11892
rect 15752 11840 15804 11892
rect 16304 11840 16356 11892
rect 18604 11840 18656 11892
rect 19432 11840 19484 11892
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 17592 11772 17644 11824
rect 18880 11772 18932 11824
rect 13820 11704 13872 11756
rect 14648 11704 14700 11756
rect 15844 11704 15896 11756
rect 16028 11747 16080 11756
rect 16028 11713 16037 11747
rect 16037 11713 16071 11747
rect 16071 11713 16080 11747
rect 16028 11704 16080 11713
rect 16580 11704 16632 11756
rect 16488 11636 16540 11688
rect 17316 11704 17368 11756
rect 19340 11704 19392 11756
rect 14004 11568 14056 11620
rect 10048 11500 10100 11552
rect 12440 11500 12492 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 13636 11500 13688 11552
rect 13912 11543 13964 11552
rect 13912 11509 13921 11543
rect 13921 11509 13955 11543
rect 13955 11509 13964 11543
rect 16120 11568 16172 11620
rect 13912 11500 13964 11509
rect 14556 11500 14608 11552
rect 15936 11500 15988 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 17132 11500 17184 11552
rect 17500 11568 17552 11620
rect 18604 11568 18656 11620
rect 20076 11568 20128 11620
rect 17776 11500 17828 11552
rect 19064 11500 19116 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 9404 11296 9456 11348
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 12072 11296 12124 11348
rect 14280 11339 14332 11348
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 15752 11296 15804 11348
rect 9128 11228 9180 11280
rect 10508 11228 10560 11280
rect 10692 11228 10744 11280
rect 13912 11228 13964 11280
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 11888 11160 11940 11212
rect 12072 11160 12124 11212
rect 12348 11160 12400 11212
rect 17040 11296 17092 11348
rect 17592 11296 17644 11348
rect 16212 11228 16264 11280
rect 17316 11228 17368 11280
rect 19800 11228 19852 11280
rect 16764 11160 16816 11212
rect 18696 11203 18748 11212
rect 18696 11169 18705 11203
rect 18705 11169 18739 11203
rect 18739 11169 18748 11203
rect 18696 11160 18748 11169
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 9680 11092 9732 11144
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 13360 11092 13412 11144
rect 15384 11092 15436 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 9312 11024 9364 11033
rect 13636 11024 13688 11076
rect 16120 11024 16172 11076
rect 11152 10956 11204 11008
rect 12992 10956 13044 11008
rect 15292 10999 15344 11008
rect 15292 10965 15301 10999
rect 15301 10965 15335 10999
rect 15335 10965 15344 10999
rect 15292 10956 15344 10965
rect 17684 11024 17736 11076
rect 17040 10956 17092 11008
rect 17592 10956 17644 11008
rect 19248 11024 19300 11076
rect 18512 10956 18564 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 9680 10752 9732 10804
rect 9128 10616 9180 10668
rect 11152 10684 11204 10736
rect 11612 10752 11664 10804
rect 12348 10752 12400 10804
rect 12440 10795 12492 10804
rect 12440 10761 12449 10795
rect 12449 10761 12483 10795
rect 12483 10761 12492 10795
rect 12440 10752 12492 10761
rect 12900 10752 12952 10804
rect 15660 10752 15712 10804
rect 19156 10752 19208 10804
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15292 10616 15344 10668
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 18696 10616 18748 10668
rect 19248 10659 19300 10668
rect 19248 10625 19257 10659
rect 19257 10625 19291 10659
rect 19291 10625 19300 10659
rect 19248 10616 19300 10625
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 12532 10548 12584 10600
rect 13176 10548 13228 10600
rect 14372 10548 14424 10600
rect 14556 10548 14608 10600
rect 15476 10548 15528 10600
rect 17040 10548 17092 10600
rect 17868 10548 17920 10600
rect 19340 10548 19392 10600
rect 10692 10480 10744 10532
rect 15292 10480 15344 10532
rect 17500 10480 17552 10532
rect 18788 10480 18840 10532
rect 20536 10480 20588 10532
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 11612 10412 11664 10464
rect 12440 10412 12492 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13728 10412 13780 10464
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 14004 10412 14056 10464
rect 17592 10412 17644 10464
rect 18604 10455 18656 10464
rect 18604 10421 18613 10455
rect 18613 10421 18647 10455
rect 18647 10421 18656 10455
rect 18604 10412 18656 10421
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 19064 10412 19116 10464
rect 20076 10412 20128 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 9036 10208 9088 10260
rect 9312 10140 9364 10192
rect 11704 10140 11756 10192
rect 11152 10072 11204 10124
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 11888 10208 11940 10260
rect 12440 10208 12492 10260
rect 13452 10208 13504 10260
rect 14556 10208 14608 10260
rect 15016 10208 15068 10260
rect 15108 10208 15160 10260
rect 16764 10208 16816 10260
rect 17684 10208 17736 10260
rect 17960 10208 18012 10260
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 14004 10140 14056 10192
rect 17408 10140 17460 10192
rect 18512 10183 18564 10192
rect 18512 10149 18521 10183
rect 18521 10149 18555 10183
rect 18555 10149 18564 10183
rect 18512 10140 18564 10149
rect 15384 10072 15436 10124
rect 15568 10115 15620 10124
rect 15568 10081 15602 10115
rect 15602 10081 15620 10115
rect 15568 10072 15620 10081
rect 17684 10072 17736 10124
rect 19340 10140 19392 10192
rect 19248 10072 19300 10124
rect 19708 10072 19760 10124
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 14004 10004 14056 10056
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 15108 10004 15160 10056
rect 15200 10004 15252 10056
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 18788 10047 18840 10056
rect 18788 10013 18797 10047
rect 18797 10013 18831 10047
rect 18831 10013 18840 10047
rect 18788 10004 18840 10013
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 12624 9868 12676 9920
rect 14372 9936 14424 9988
rect 15016 9936 15068 9988
rect 18972 9868 19024 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 14004 9664 14056 9716
rect 15384 9664 15436 9716
rect 17408 9664 17460 9716
rect 11152 9596 11204 9648
rect 11980 9528 12032 9580
rect 14188 9528 14240 9580
rect 15016 9528 15068 9580
rect 15568 9528 15620 9580
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 7932 9460 7984 9512
rect 8852 9460 8904 9512
rect 9312 9460 9364 9512
rect 10600 9460 10652 9512
rect 9864 9392 9916 9444
rect 10968 9392 11020 9444
rect 11428 9460 11480 9512
rect 12992 9460 13044 9512
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 14372 9460 14424 9512
rect 14648 9460 14700 9512
rect 16396 9460 16448 9512
rect 16856 9460 16908 9512
rect 17776 9460 17828 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 19340 9460 19392 9512
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 14740 9392 14792 9444
rect 17592 9392 17644 9444
rect 9220 9324 9272 9376
rect 13728 9324 13780 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15936 9367 15988 9376
rect 15016 9324 15068 9333
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 16120 9324 16172 9376
rect 17500 9324 17552 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 20076 9367 20128 9376
rect 20076 9333 20085 9367
rect 20085 9333 20119 9367
rect 20119 9333 20128 9367
rect 20076 9324 20128 9333
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 9680 9120 9732 9172
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 11704 9120 11756 9172
rect 9772 9052 9824 9104
rect 11152 9052 11204 9104
rect 9864 8984 9916 9036
rect 10600 8984 10652 9036
rect 10876 8984 10928 9036
rect 14096 9120 14148 9172
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 16212 9120 16264 9172
rect 17868 9120 17920 9172
rect 13728 9052 13780 9104
rect 15200 9052 15252 9104
rect 8208 8916 8260 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 17040 9052 17092 9104
rect 16396 8984 16448 9036
rect 17592 9027 17644 9036
rect 17592 8993 17601 9027
rect 17601 8993 17635 9027
rect 17635 8993 17644 9027
rect 17592 8984 17644 8993
rect 19432 9052 19484 9104
rect 19984 9120 20036 9172
rect 20536 9052 20588 9104
rect 19340 8984 19392 9036
rect 10968 8848 11020 8900
rect 17040 8848 17092 8900
rect 18052 8848 18104 8900
rect 8668 8780 8720 8832
rect 10784 8780 10836 8832
rect 11612 8780 11664 8832
rect 13636 8780 13688 8832
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 19708 8848 19760 8900
rect 19984 8780 20036 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 10416 8576 10468 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 16488 8576 16540 8628
rect 17592 8576 17644 8628
rect 11612 8508 11664 8560
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 10968 8440 11020 8492
rect 3424 8372 3476 8424
rect 6920 8304 6972 8356
rect 9864 8372 9916 8424
rect 12072 8372 12124 8424
rect 9772 8304 9824 8356
rect 10140 8304 10192 8356
rect 12716 8440 12768 8492
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 16396 8483 16448 8492
rect 16396 8449 16405 8483
rect 16405 8449 16439 8483
rect 16439 8449 16448 8483
rect 16396 8440 16448 8449
rect 16856 8440 16908 8492
rect 17132 8440 17184 8492
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 19432 8508 19484 8560
rect 20168 8440 20220 8492
rect 20628 8440 20680 8492
rect 14096 8372 14148 8424
rect 20076 8372 20128 8424
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 13452 8304 13504 8356
rect 14188 8347 14240 8356
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 13820 8279 13872 8288
rect 13820 8245 13829 8279
rect 13829 8245 13863 8279
rect 13863 8245 13872 8279
rect 13820 8236 13872 8245
rect 14188 8313 14197 8347
rect 14197 8313 14231 8347
rect 14231 8313 14240 8347
rect 14188 8304 14240 8313
rect 15568 8304 15620 8356
rect 17868 8304 17920 8356
rect 15384 8236 15436 8288
rect 15476 8236 15528 8288
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 16396 8236 16448 8288
rect 19984 8279 20036 8288
rect 19984 8245 19993 8279
rect 19993 8245 20027 8279
rect 20027 8245 20036 8279
rect 19984 8236 20036 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 11888 8032 11940 8084
rect 12900 8032 12952 8084
rect 9956 7964 10008 8016
rect 11796 7964 11848 8016
rect 13176 7964 13228 8016
rect 9680 7896 9732 7948
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 10968 7896 11020 7948
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 10784 7760 10836 7812
rect 11980 7692 12032 7744
rect 12716 7692 12768 7744
rect 13820 8032 13872 8084
rect 16120 8032 16172 8084
rect 19340 8032 19392 8084
rect 20168 8032 20220 8084
rect 20444 8032 20496 8084
rect 14372 7896 14424 7948
rect 14740 7896 14792 7948
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 16396 7896 16448 7948
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13452 7828 13504 7880
rect 15752 7828 15804 7880
rect 17408 7896 17460 7948
rect 18604 7896 18656 7948
rect 20628 7964 20680 8016
rect 13176 7692 13228 7744
rect 17592 7692 17644 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10232 7488 10284 7540
rect 10784 7488 10836 7540
rect 12808 7531 12860 7540
rect 12808 7497 12817 7531
rect 12817 7497 12851 7531
rect 12851 7497 12860 7531
rect 12808 7488 12860 7497
rect 12992 7488 13044 7540
rect 12072 7420 12124 7472
rect 12348 7420 12400 7472
rect 13452 7420 13504 7472
rect 16672 7488 16724 7540
rect 16856 7531 16908 7540
rect 16856 7497 16865 7531
rect 16865 7497 16899 7531
rect 16899 7497 16908 7531
rect 16856 7488 16908 7497
rect 10600 7352 10652 7404
rect 13176 7352 13228 7404
rect 13728 7352 13780 7404
rect 14740 7352 14792 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9864 7216 9916 7268
rect 12808 7216 12860 7268
rect 9956 7148 10008 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 12256 7148 12308 7200
rect 13820 7284 13872 7336
rect 14924 7284 14976 7336
rect 15752 7327 15804 7336
rect 15752 7293 15786 7327
rect 15786 7293 15804 7327
rect 15752 7284 15804 7293
rect 16028 7284 16080 7336
rect 18788 7284 18840 7336
rect 20352 7327 20404 7336
rect 20352 7293 20361 7327
rect 20361 7293 20395 7327
rect 20395 7293 20404 7327
rect 20352 7284 20404 7293
rect 15108 7216 15160 7268
rect 18696 7216 18748 7268
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 18788 7148 18840 7200
rect 19064 7148 19116 7200
rect 19156 7148 19208 7200
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 12716 6944 12768 6996
rect 12808 6944 12860 6996
rect 13268 6944 13320 6996
rect 13820 6987 13872 6996
rect 13820 6953 13829 6987
rect 13829 6953 13863 6987
rect 13863 6953 13872 6987
rect 13820 6944 13872 6953
rect 15200 6944 15252 6996
rect 16212 6944 16264 6996
rect 18052 6944 18104 6996
rect 18236 6987 18288 6996
rect 18236 6953 18245 6987
rect 18245 6953 18279 6987
rect 18279 6953 18288 6987
rect 18236 6944 18288 6953
rect 20628 6944 20680 6996
rect 9772 6876 9824 6928
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10692 6876 10744 6928
rect 13912 6876 13964 6928
rect 14096 6876 14148 6928
rect 18512 6876 18564 6928
rect 9680 6740 9732 6792
rect 9772 6740 9824 6792
rect 11336 6808 11388 6860
rect 11971 6851 12023 6860
rect 11971 6817 12003 6851
rect 12003 6817 12023 6851
rect 11971 6808 12023 6817
rect 13452 6808 13504 6860
rect 15568 6808 15620 6860
rect 16028 6808 16080 6860
rect 16488 6851 16540 6860
rect 16488 6817 16497 6851
rect 16497 6817 16531 6851
rect 16531 6817 16540 6851
rect 16488 6808 16540 6817
rect 17224 6808 17276 6860
rect 19800 6808 19852 6860
rect 20628 6808 20680 6860
rect 10968 6740 11020 6792
rect 14372 6783 14424 6792
rect 10876 6672 10928 6724
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 14556 6740 14608 6792
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 16212 6740 16264 6792
rect 10140 6604 10192 6656
rect 11888 6604 11940 6656
rect 15384 6672 15436 6724
rect 15568 6672 15620 6724
rect 17592 6740 17644 6792
rect 18604 6740 18656 6792
rect 19064 6740 19116 6792
rect 13176 6604 13228 6656
rect 14556 6604 14608 6656
rect 16672 6604 16724 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 10048 6400 10100 6452
rect 11796 6400 11848 6452
rect 13544 6400 13596 6452
rect 19616 6400 19668 6452
rect 20628 6443 20680 6452
rect 20628 6409 20637 6443
rect 20637 6409 20671 6443
rect 20671 6409 20680 6443
rect 20628 6400 20680 6409
rect 12256 6332 12308 6384
rect 15292 6332 15344 6384
rect 10324 6264 10376 6316
rect 10968 6264 11020 6316
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 13176 6264 13228 6316
rect 17132 6264 17184 6316
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 18972 6264 19024 6316
rect 8392 6196 8444 6248
rect 9680 6196 9732 6248
rect 10600 6196 10652 6248
rect 4068 6128 4120 6180
rect 10968 6128 11020 6180
rect 11152 6196 11204 6248
rect 11888 6196 11940 6248
rect 14004 6196 14056 6248
rect 14188 6196 14240 6248
rect 18512 6196 18564 6248
rect 19064 6196 19116 6248
rect 19892 6196 19944 6248
rect 20444 6196 20496 6248
rect 11796 6128 11848 6180
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 13912 6060 13964 6112
rect 14280 6060 14332 6112
rect 15108 6128 15160 6180
rect 15292 6060 15344 6112
rect 15752 6060 15804 6112
rect 16856 6128 16908 6180
rect 17960 6128 18012 6180
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 18696 6103 18748 6112
rect 18696 6069 18705 6103
rect 18705 6069 18739 6103
rect 18739 6069 18748 6103
rect 18696 6060 18748 6069
rect 19248 6060 19300 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 9772 5899 9824 5908
rect 9772 5865 9781 5899
rect 9781 5865 9815 5899
rect 9815 5865 9824 5899
rect 9772 5856 9824 5865
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 12440 5856 12492 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 16488 5856 16540 5908
rect 17224 5856 17276 5908
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 18972 5856 19024 5908
rect 19524 5856 19576 5908
rect 20260 5856 20312 5908
rect 13176 5788 13228 5840
rect 14004 5788 14056 5840
rect 15384 5788 15436 5840
rect 15844 5788 15896 5840
rect 17132 5788 17184 5840
rect 8392 5720 8444 5772
rect 10876 5720 10928 5772
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 15200 5720 15252 5772
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 13268 5695 13320 5704
rect 10324 5652 10376 5661
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 13636 5695 13688 5704
rect 13636 5661 13645 5695
rect 13645 5661 13679 5695
rect 13679 5661 13688 5695
rect 13636 5652 13688 5661
rect 15108 5652 15160 5704
rect 17960 5720 18012 5772
rect 16672 5652 16724 5704
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 18512 5652 18564 5704
rect 13084 5584 13136 5636
rect 16304 5584 16356 5636
rect 16580 5584 16632 5636
rect 13544 5516 13596 5568
rect 13912 5516 13964 5568
rect 19984 5516 20036 5568
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 10232 5312 10284 5364
rect 10876 5312 10928 5364
rect 12992 5312 13044 5364
rect 15844 5312 15896 5364
rect 17132 5312 17184 5364
rect 19892 5355 19944 5364
rect 19892 5321 19901 5355
rect 19901 5321 19935 5355
rect 19935 5321 19944 5355
rect 19892 5312 19944 5321
rect 20444 5244 20496 5296
rect 10784 5176 10836 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 15568 5176 15620 5228
rect 17224 5176 17276 5228
rect 17868 5176 17920 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 11704 5108 11756 5160
rect 13636 5108 13688 5160
rect 15108 5108 15160 5160
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 16488 5108 16540 5160
rect 20260 5108 20312 5160
rect 11704 4972 11756 5024
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 13268 5040 13320 5092
rect 16028 5040 16080 5092
rect 18604 5040 18656 5092
rect 20076 5040 20128 5092
rect 20720 5040 20772 5092
rect 12992 4972 13044 4981
rect 15844 4972 15896 5024
rect 17776 4972 17828 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 6092 4768 6144 4820
rect 13084 4700 13136 4752
rect 13268 4768 13320 4820
rect 15200 4768 15252 4820
rect 17040 4768 17092 4820
rect 18788 4768 18840 4820
rect 19156 4811 19208 4820
rect 19156 4777 19165 4811
rect 19165 4777 19199 4811
rect 19199 4777 19208 4811
rect 19156 4768 19208 4777
rect 19248 4768 19300 4820
rect 11704 4632 11756 4684
rect 13820 4632 13872 4684
rect 14004 4632 14056 4684
rect 16764 4700 16816 4752
rect 17960 4700 18012 4752
rect 16580 4632 16632 4684
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 7472 4428 7524 4480
rect 17776 4496 17828 4548
rect 17960 4564 18012 4616
rect 18696 4700 18748 4752
rect 19708 4632 19760 4684
rect 19156 4564 19208 4616
rect 19800 4564 19852 4616
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 20536 4496 20588 4548
rect 14188 4428 14240 4480
rect 15292 4428 15344 4480
rect 19064 4428 19116 4480
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 12992 4224 13044 4276
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 11244 4156 11296 4208
rect 5264 4088 5316 4140
rect 8944 4088 8996 4140
rect 10140 4088 10192 4140
rect 11152 4088 11204 4140
rect 11428 4131 11480 4140
rect 11428 4097 11437 4131
rect 11437 4097 11471 4131
rect 11471 4097 11480 4131
rect 11428 4088 11480 4097
rect 13176 4156 13228 4208
rect 12900 4088 12952 4140
rect 19892 4156 19944 4208
rect 14372 4088 14424 4140
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 17316 4088 17368 4140
rect 848 4020 900 4072
rect 7564 4020 7616 4072
rect 8392 4020 8444 4072
rect 9220 4020 9272 4072
rect 2504 3952 2556 4004
rect 7472 3952 7524 4004
rect 8208 3952 8260 4004
rect 10048 3952 10100 4004
rect 296 3884 348 3936
rect 13452 4020 13504 4072
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 15752 4063 15804 4072
rect 15752 4029 15761 4063
rect 15761 4029 15795 4063
rect 15795 4029 15804 4063
rect 15752 4020 15804 4029
rect 17684 4020 17736 4072
rect 17868 4020 17920 4072
rect 18696 4020 18748 4072
rect 19800 4020 19852 4072
rect 20444 4020 20496 4072
rect 20720 4063 20772 4072
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 10416 3952 10468 4004
rect 10324 3884 10376 3936
rect 12808 3952 12860 4004
rect 13360 3952 13412 4004
rect 17224 3952 17276 4004
rect 18604 3952 18656 4004
rect 10876 3884 10928 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 15016 3884 15068 3936
rect 16396 3884 16448 3936
rect 17868 3884 17920 3936
rect 19156 3884 19208 3936
rect 22468 3884 22520 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3608 3680 3660 3732
rect 11244 3680 11296 3732
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 11704 3680 11756 3732
rect 7564 3612 7616 3664
rect 1952 3544 2004 3596
rect 10140 3544 10192 3596
rect 10324 3587 10376 3596
rect 10324 3553 10358 3587
rect 10358 3553 10376 3587
rect 10324 3544 10376 3553
rect 12440 3612 12492 3664
rect 13268 3612 13320 3664
rect 14556 3680 14608 3732
rect 13452 3612 13504 3664
rect 16120 3680 16172 3732
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 17132 3612 17184 3664
rect 8392 3476 8444 3528
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 3056 3408 3108 3460
rect 9956 3408 10008 3460
rect 4160 3340 4212 3392
rect 12348 3340 12400 3392
rect 13912 3544 13964 3596
rect 14464 3544 14516 3596
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 16120 3544 16172 3596
rect 17224 3587 17276 3596
rect 17224 3553 17233 3587
rect 17233 3553 17267 3587
rect 17267 3553 17276 3587
rect 17224 3544 17276 3553
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 19432 3544 19484 3596
rect 19524 3476 19576 3528
rect 20352 3476 20404 3528
rect 17592 3340 17644 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 5816 3136 5868 3188
rect 9036 3136 9088 3188
rect 10876 3136 10928 3188
rect 10968 3136 11020 3188
rect 13176 3136 13228 3188
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 14372 3136 14424 3188
rect 7472 3068 7524 3120
rect 10232 3068 10284 3120
rect 10324 3000 10376 3052
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 15568 3136 15620 3188
rect 16212 3136 16264 3188
rect 16948 3136 17000 3188
rect 17960 3136 18012 3188
rect 16120 3068 16172 3120
rect 20260 3068 20312 3120
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 7472 2932 7524 2984
rect 10600 2932 10652 2984
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 10876 2932 10928 2941
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 8576 2864 8628 2916
rect 4712 2796 4764 2848
rect 11336 2864 11388 2916
rect 11980 2864 12032 2916
rect 12992 2932 13044 2984
rect 15476 2932 15528 2984
rect 17592 2932 17644 2984
rect 19616 2932 19668 2984
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 14556 2864 14608 2916
rect 18696 2864 18748 2916
rect 12532 2796 12584 2848
rect 16764 2796 16816 2848
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 21364 2864 21416 2916
rect 16948 2796 17000 2805
rect 21916 2796 21968 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 12532 2592 12584 2644
rect 16948 2592 17000 2644
rect 13820 2567 13872 2576
rect 11336 2499 11388 2508
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 11980 2456 12032 2508
rect 12624 2456 12676 2508
rect 1400 2388 1452 2440
rect 13452 2456 13504 2508
rect 13820 2533 13829 2567
rect 13829 2533 13863 2567
rect 13863 2533 13872 2567
rect 13820 2524 13872 2533
rect 16764 2524 16816 2576
rect 17500 2524 17552 2576
rect 18604 2524 18656 2576
rect 15568 2456 15620 2508
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 16580 2456 16632 2465
rect 17776 2456 17828 2508
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 19524 2499 19576 2508
rect 15660 2388 15712 2440
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 16304 2388 16356 2440
rect 19524 2465 19533 2499
rect 19533 2465 19567 2499
rect 19567 2465 19576 2499
rect 19524 2456 19576 2465
rect 20352 2499 20404 2508
rect 20352 2465 20361 2499
rect 20361 2465 20395 2499
rect 20395 2465 20404 2499
rect 20352 2456 20404 2465
rect 13636 2320 13688 2372
rect 18696 2320 18748 2372
rect 11980 2252 12032 2304
rect 13084 2252 13136 2304
rect 16948 2252 17000 2304
rect 17500 2295 17552 2304
rect 17500 2261 17509 2295
rect 17509 2261 17543 2295
rect 17543 2261 17552 2295
rect 17500 2252 17552 2261
rect 19064 2252 19116 2304
rect 19616 2252 19668 2304
rect 20812 2252 20864 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 9680 1368 9732 1420
rect 10968 1368 11020 1420
rect 10232 1096 10284 1148
rect 12072 1096 12124 1148
<< metal2 >>
rect 294 22320 350 22800
rect 846 22320 902 22800
rect 1398 22320 1454 22800
rect 1950 22320 2006 22800
rect 2502 22320 2558 22800
rect 3054 22320 3110 22800
rect 3606 22320 3662 22800
rect 4158 22320 4214 22800
rect 4710 22320 4766 22800
rect 5262 22320 5318 22800
rect 5814 22320 5870 22800
rect 6366 22320 6422 22800
rect 6918 22320 6974 22800
rect 7470 22320 7526 22800
rect 8022 22320 8078 22800
rect 8574 22320 8630 22800
rect 9126 22320 9182 22800
rect 9678 22320 9734 22800
rect 10230 22320 10286 22800
rect 10782 22320 10838 22800
rect 11334 22320 11390 22800
rect 11978 22320 12034 22800
rect 12530 22320 12586 22800
rect 13082 22320 13138 22800
rect 13634 22320 13690 22800
rect 14186 22320 14242 22800
rect 14738 22320 14794 22800
rect 15290 22320 15346 22800
rect 15842 22320 15898 22800
rect 16394 22320 16450 22800
rect 16946 22320 17002 22800
rect 17498 22320 17554 22800
rect 18050 22320 18106 22800
rect 18602 22320 18658 22800
rect 18970 22536 19026 22545
rect 18970 22471 19026 22480
rect 308 18698 336 22320
rect 296 18692 348 18698
rect 296 18634 348 18640
rect 860 17542 888 22320
rect 1412 19174 1440 22320
rect 1964 19242 1992 22320
rect 1952 19236 2004 19242
rect 1952 19178 2004 19184
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 2516 18426 2544 22320
rect 3068 19242 3096 22320
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 2976 18970 3004 19178
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 3620 18222 3648 22320
rect 4172 18358 4200 22320
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4724 18290 4752 22320
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 5276 18034 5304 22320
rect 5828 18086 5856 22320
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 5816 18080 5868 18086
rect 5276 18006 5580 18034
rect 5816 18022 5868 18028
rect 848 17536 900 17542
rect 848 17478 900 17484
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 3422 17232 3478 17241
rect 3422 17167 3478 17176
rect 3436 8430 3464 17167
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 5552 14958 5580 18006
rect 6196 15026 6224 18226
rect 6380 18222 6408 22320
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6932 16794 6960 22320
rect 7484 20330 7512 22320
rect 8036 20346 8064 22320
rect 7472 20324 7524 20330
rect 8036 20318 8248 20346
rect 7472 20266 7524 20272
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7760 18834 7788 19246
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7668 18086 7696 18634
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7484 16794 7512 18022
rect 7760 17882 7788 18770
rect 8220 18630 8248 20318
rect 8588 19174 8616 22320
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8772 20058 8800 20198
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8484 19168 8536 19174
rect 8482 19136 8484 19145
rect 8576 19168 8628 19174
rect 8536 19136 8538 19145
rect 8576 19110 8628 19116
rect 8482 19071 8538 19080
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7760 17134 7788 17818
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8312 17338 8340 17682
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8496 17270 8524 17478
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6932 15570 6960 15982
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5817 4108 6122
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 6104 4826 6132 14894
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6840 14482 6868 14826
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 848 4072 900 4078
rect 848 4014 900 4020
rect 296 3936 348 3942
rect 296 3878 348 3884
rect 308 480 336 3878
rect 860 480 888 4014
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 480 1440 2382
rect 1964 480 1992 3538
rect 2516 480 2544 3946
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3068 480 3096 3402
rect 3620 480 3648 3674
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 480 4200 3334
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 480 4752 2790
rect 5276 480 5304 4082
rect 6366 3496 6422 3505
rect 6366 3431 6422 3440
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5828 480 5856 3130
rect 6380 480 6408 3431
rect 6932 480 6960 8298
rect 7484 4486 7512 16730
rect 7668 16590 7696 17002
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7760 16522 7788 17070
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8220 16794 8248 17070
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7656 16040 7708 16046
rect 7760 16028 7788 16458
rect 8220 16250 8248 16526
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 7708 16000 7788 16028
rect 7656 15982 7708 15988
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 15026 7604 15302
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7576 14550 7604 14962
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8496 14074 8524 14418
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8588 13938 8616 18226
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9518 7972 9998
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8634 8248 8910
rect 8680 8838 8708 18158
rect 8864 17882 8892 18770
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 9048 17338 9076 18226
rect 9140 18154 9168 22320
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9232 18970 9260 19178
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9232 18290 9260 18906
rect 9692 18329 9720 22320
rect 10244 20618 10272 22320
rect 10244 20590 10732 20618
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 9770 19816 9826 19825
rect 9770 19751 9772 19760
rect 9824 19751 9826 19760
rect 9772 19722 9824 19728
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9678 18320 9734 18329
rect 9220 18284 9272 18290
rect 9678 18255 9734 18264
rect 9220 18226 9272 18232
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9692 17882 9720 18090
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9128 17808 9180 17814
rect 9128 17750 9180 17756
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8772 16590 8800 17138
rect 9140 16998 9168 17750
rect 9508 17202 9536 17818
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9048 16794 9076 16934
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8864 15094 8892 15914
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 9048 14414 9076 15030
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8956 12986 8984 13806
rect 9140 13682 9168 16934
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9048 13654 9168 13682
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8864 8498 8892 9454
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8404 6254 8432 7278
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8404 5778 8432 6190
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 8404 4078 8432 5714
rect 8956 4146 8984 12922
rect 9048 10266 9076 13654
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11286 9168 12038
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9140 10674 9168 11222
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9232 10470 9260 16594
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16114 9444 16458
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14618 9352 14758
rect 9508 14618 9536 16594
rect 9692 16250 9720 16934
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9784 15570 9812 18838
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 16998 9904 18022
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9508 13394 9536 14554
rect 9692 14550 9720 15506
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9876 15162 9904 15438
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9784 14482 9812 14826
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 13530 9720 14350
rect 9876 14278 9904 14962
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 13938 9904 14214
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9692 13394 9720 13466
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 12782 9720 13330
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9600 12374 9628 12582
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9692 12306 9720 12718
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 12102 9720 12242
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11354 9444 11630
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7484 3126 7512 3946
rect 7576 3670 7604 4014
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7484 480 7512 2926
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 762 8248 3946
rect 8404 3534 8432 4014
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 9048 3194 9076 10202
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8036 734 8248 762
rect 8036 480 8064 734
rect 8588 480 8616 2858
rect 9140 480 9168 10406
rect 9324 10198 9352 11018
rect 9692 10810 9720 11086
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9518 9352 9862
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 8974 9260 9318
rect 9692 9178 9720 9998
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 9110 9812 10542
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9876 9042 9904 9386
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9232 4078 9260 8910
rect 9876 8430 9904 8978
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7002 9720 7890
rect 9784 7546 9812 8298
rect 9968 8022 9996 18770
rect 10060 18222 10088 19654
rect 10244 19514 10272 19858
rect 10508 19848 10560 19854
rect 10428 19796 10508 19802
rect 10428 19790 10560 19796
rect 10428 19774 10548 19790
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10152 18442 10180 19246
rect 10336 19009 10364 19246
rect 10428 19242 10456 19774
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 10322 19000 10378 19009
rect 10322 18935 10378 18944
rect 10322 18864 10378 18873
rect 10322 18799 10378 18808
rect 10152 18414 10272 18442
rect 10244 18358 10272 18414
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10152 17882 10180 18294
rect 10336 18170 10364 18799
rect 10244 18142 10364 18170
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10060 13977 10088 17682
rect 10244 15586 10272 18142
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 17746 10364 18022
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10428 17678 10456 19178
rect 10506 19000 10562 19009
rect 10506 18935 10562 18944
rect 10520 18766 10548 18935
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10520 17202 10548 18362
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10140 15564 10192 15570
rect 10244 15558 10364 15586
rect 10140 15506 10192 15512
rect 10046 13968 10102 13977
rect 10046 13903 10102 13912
rect 10152 13841 10180 15506
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 12850 10180 13670
rect 10244 13462 10272 14758
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10244 12442 10272 12650
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11354 10088 11494
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6934 9812 7482
rect 10152 7426 10180 8298
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7546 10272 7890
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10152 7398 10272 7426
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9692 6254 9720 6734
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9784 5914 9812 6734
rect 9876 6458 9904 7210
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9968 3466 9996 7142
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10152 5914 10180 6598
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10244 5794 10272 7398
rect 10336 6474 10364 15558
rect 10414 13968 10470 13977
rect 10414 13903 10470 13912
rect 10428 10033 10456 13903
rect 10520 11286 10548 16934
rect 10612 13716 10640 19994
rect 10704 19242 10732 20590
rect 10796 19258 10824 22320
rect 11348 20058 11376 22320
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11900 19922 11928 20266
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11900 19530 11928 19858
rect 11716 19502 11928 19530
rect 10796 19242 10916 19258
rect 10692 19236 10744 19242
rect 10796 19236 10928 19242
rect 10796 19230 10876 19236
rect 10692 19178 10744 19184
rect 10876 19178 10928 19184
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10704 18290 10732 18838
rect 10796 18290 10824 19110
rect 11624 18902 11652 19110
rect 11612 18896 11664 18902
rect 11612 18838 11664 18844
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 15026 10732 16934
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10888 16114 10916 16730
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10980 15978 11008 16730
rect 11072 15994 11100 18158
rect 11716 17542 11744 19502
rect 11992 19394 12020 22320
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 11808 19366 12020 19394
rect 11808 18970 11836 19366
rect 12084 19258 12112 19790
rect 12256 19712 12308 19718
rect 12544 19700 12572 22320
rect 13096 20058 13124 22320
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12256 19654 12308 19660
rect 12452 19672 12572 19700
rect 11992 19242 12112 19258
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 11980 19236 12112 19242
rect 12032 19230 12112 19236
rect 11980 19178 12032 19184
rect 11992 18970 12020 19178
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11164 16130 11192 17478
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11164 16102 11376 16130
rect 10968 15972 11020 15978
rect 11072 15966 11284 15994
rect 10968 15914 11020 15920
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15570 10824 15846
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10888 15162 10916 15438
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10980 15026 11008 15914
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10966 14920 11022 14929
rect 11072 14890 11100 15846
rect 11256 15450 11284 15966
rect 11348 15706 11376 16102
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11164 15422 11284 15450
rect 10966 14855 11022 14864
rect 11060 14884 11112 14890
rect 10980 13938 11008 14855
rect 11060 14826 11112 14832
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10692 13728 10744 13734
rect 10612 13688 10692 13716
rect 10692 13670 10744 13676
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 11762 10640 12242
rect 10704 11830 10732 13670
rect 10888 13190 10916 13874
rect 11072 13394 11100 14214
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12442 10916 13126
rect 11164 12986 11192 15422
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11520 14952 11572 14958
rect 11624 14929 11652 17070
rect 11716 16658 11744 17138
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11716 16114 11744 16594
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11900 15638 11928 16594
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 15026 11836 15506
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11520 14894 11572 14900
rect 11610 14920 11666 14929
rect 11532 14482 11560 14894
rect 11610 14855 11666 14864
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11348 13530 11376 13806
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10888 12238 10916 12378
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10980 12170 11008 12582
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10704 11370 10732 11766
rect 10612 11342 10732 11370
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10612 11132 10640 11342
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10520 11104 10640 11132
rect 10414 10024 10470 10033
rect 10414 9959 10470 9968
rect 10428 8634 10456 9959
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10336 6446 10456 6474
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10060 5766 10272 5794
rect 10060 4010 10088 5766
rect 10336 5710 10364 6258
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10244 5370 10272 5646
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10152 3602 10180 4082
rect 10428 4010 10456 6446
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3602 10364 3878
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 10232 3120 10284 3126
rect 10230 3088 10232 3097
rect 10284 3088 10286 3097
rect 10336 3058 10364 3538
rect 10230 3023 10286 3032
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10520 2836 10548 11104
rect 10704 10538 10732 11222
rect 10888 11218 10916 12038
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10612 9518 10640 9998
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10612 8634 10640 8978
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10612 7410 10640 8570
rect 10704 7426 10732 10474
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8401 10824 8774
rect 10888 8634 10916 8978
rect 10980 8906 11008 9386
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10980 8498 11008 8842
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10782 8392 10838 8401
rect 10782 8327 10838 8336
rect 10980 7954 11008 8434
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10796 7546 10824 7754
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10600 7404 10652 7410
rect 10704 7398 10824 7426
rect 10600 7346 10652 7352
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10704 6934 10732 7142
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10612 2990 10640 6190
rect 10796 5234 10824 7398
rect 10888 6730 10916 7822
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10888 5778 10916 6666
rect 10980 6322 11008 6734
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 6186 11008 6258
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10888 5370 10916 5714
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10980 5234 11008 6122
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3194 10916 3878
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10520 2808 10824 2836
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9692 480 9720 1362
rect 10232 1148 10284 1154
rect 10232 1090 10284 1096
rect 10244 480 10272 1090
rect 10796 480 10824 2808
rect 10888 1601 10916 2926
rect 10874 1592 10930 1601
rect 10874 1527 10930 1536
rect 10980 1426 11008 3130
rect 10968 1420 11020 1426
rect 10968 1362 11020 1368
rect 11072 1306 11100 12242
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10742 11192 10950
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 10810 11652 14855
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11716 14074 11744 14758
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11808 14006 11836 14758
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11900 13938 11928 14418
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9654 11192 10066
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11164 9110 11192 9590
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11440 9178 11468 9454
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11624 8838 11652 10406
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11716 9178 11744 10134
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11334 6896 11390 6905
rect 11334 6831 11336 6840
rect 11388 6831 11390 6840
rect 11336 6802 11388 6808
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11164 4146 11192 6190
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11256 3738 11284 4150
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11440 3738 11468 4082
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11624 2990 11652 8502
rect 11716 5166 11744 9114
rect 11808 8022 11836 13670
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11900 10674 11928 11154
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11900 10266 11928 10610
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11992 9586 12020 18158
rect 12084 17762 12112 19110
rect 12176 18970 12204 19246
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12084 17734 12204 17762
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12084 16794 12112 17614
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12176 16266 12204 17734
rect 12268 17202 12296 19654
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12360 19009 12388 19110
rect 12346 19000 12402 19009
rect 12346 18935 12402 18944
rect 12452 18426 12480 19672
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 19174 12572 19246
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18834 12572 19110
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12254 16552 12310 16561
rect 12254 16487 12310 16496
rect 12084 16238 12204 16266
rect 12268 16250 12296 16487
rect 12256 16244 12308 16250
rect 12084 13462 12112 16238
rect 12256 16186 12308 16192
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12176 15978 12204 16118
rect 12360 15994 12388 17478
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12452 16561 12480 16662
rect 12438 16552 12494 16561
rect 12438 16487 12494 16496
rect 12544 16046 12572 17614
rect 12636 16250 12664 17682
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12728 16182 12756 17070
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12532 16040 12584 16046
rect 12164 15972 12216 15978
rect 12360 15966 12480 15994
rect 12532 15982 12584 15988
rect 12164 15914 12216 15920
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 12084 13190 12112 13398
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11762 12112 12242
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12084 11354 12112 11698
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11900 8090 11928 8910
rect 12084 8430 12112 11154
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11992 6866 12020 7686
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11971 6860 12023 6866
rect 11971 6802 12023 6808
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11808 6186 11836 6394
rect 11900 6254 11928 6598
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4690 11744 4966
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11716 3738 11744 4626
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11716 3534 11744 3674
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11348 2514 11376 2858
rect 11992 2514 12020 2858
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11072 1278 11376 1306
rect 11348 480 11376 1278
rect 11992 480 12020 2246
rect 12084 1154 12112 7414
rect 12176 1601 12204 15914
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 14226 12296 15846
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12360 14618 12388 14962
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12268 14198 12388 14226
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12268 7449 12296 13670
rect 12360 11218 12388 14198
rect 12452 13734 12480 15966
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12622 13968 12678 13977
rect 12622 13903 12678 13912
rect 12636 13870 12664 13903
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13530 12572 13670
rect 12728 13530 12756 14894
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12728 12986 12756 13330
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12820 12782 12848 19858
rect 13648 19242 13676 22320
rect 14200 20058 14228 22320
rect 14752 20346 14780 22320
rect 14568 20318 14780 20346
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 14372 19916 14424 19922
rect 14372 19858 14424 19864
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13004 18902 13032 19110
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 13096 18426 13124 18838
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13188 18290 13216 18362
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13082 18184 13138 18193
rect 13082 18119 13138 18128
rect 13096 18086 13124 18119
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13188 17898 13216 18226
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13096 17870 13216 17898
rect 13280 17882 13308 18022
rect 13268 17876 13320 17882
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12912 17270 12940 17614
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12992 17264 13044 17270
rect 12992 17206 13044 17212
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12912 15366 12940 16594
rect 13004 15910 13032 17206
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13096 15586 13124 17870
rect 13268 17818 13320 17824
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13188 15706 13216 17750
rect 13464 17338 13492 18226
rect 13556 17678 13584 19110
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13556 17202 13584 17614
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16794 13308 16934
rect 13268 16788 13320 16794
rect 13648 16776 13676 17818
rect 13268 16730 13320 16736
rect 13556 16748 13676 16776
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13280 16114 13308 16390
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13372 16046 13400 16390
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13096 15558 13216 15586
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 14414 12940 15302
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14618 13124 14758
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13433 12940 13670
rect 12898 13424 12954 13433
rect 13096 13394 13124 14214
rect 12898 13359 12954 13368
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12452 11898 12480 12582
rect 12912 11898 12940 12582
rect 13004 12306 13032 12718
rect 13096 12442 13124 12786
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12452 10810 12480 11494
rect 12912 10810 12940 11494
rect 13004 11014 13032 11494
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12360 7478 12388 10746
rect 13188 10606 13216 15558
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13268 14544 13320 14550
rect 13266 14512 13268 14521
rect 13320 14512 13322 14521
rect 13266 14447 13322 14456
rect 13464 14074 13492 14758
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13266 11248 13322 11257
rect 13266 11183 13322 11192
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12348 7472 12400 7478
rect 12254 7440 12310 7449
rect 12348 7414 12400 7420
rect 12254 7375 12310 7384
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 6390 12296 7142
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5914 12480 6054
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12452 3482 12480 3606
rect 12360 3454 12480 3482
rect 12360 3398 12388 3454
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12544 2854 12572 10542
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12162 1592 12218 1601
rect 12162 1527 12218 1536
rect 12072 1148 12124 1154
rect 12072 1090 12124 1096
rect 12544 480 12572 2586
rect 12636 2514 12664 9862
rect 12912 8922 12940 10406
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13004 9042 13032 9454
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12912 8894 13032 8922
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12728 7750 12756 8434
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12820 7546 12848 8298
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 8090 12940 8230
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13004 7970 13032 8894
rect 13176 8016 13228 8022
rect 12912 7942 13032 7970
rect 13174 7984 13176 7993
rect 13228 7984 13230 7993
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12820 7002 12848 7210
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12728 6225 12756 6938
rect 12714 6216 12770 6225
rect 12714 6151 12770 6160
rect 12820 4010 12848 6938
rect 12912 4146 12940 7942
rect 13174 7919 13230 7928
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 7546 13032 7822
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13188 7410 13216 7686
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13280 7002 13308 11183
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 6322 13216 6598
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 5370 13032 5714
rect 13096 5642 13124 6258
rect 13188 5846 13216 6258
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13096 5234 13124 5578
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4282 13032 4966
rect 13096 4758 13124 5170
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 13188 4214 13216 5782
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13280 5098 13308 5646
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13280 4826 13308 5034
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13372 4706 13400 11086
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13464 8362 13492 10202
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13464 7478 13492 7822
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13280 4678 13400 4706
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 13280 3670 13308 4678
rect 13464 4078 13492 6802
rect 13556 6458 13584 16748
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13648 16182 13676 16594
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13634 16008 13690 16017
rect 13634 15943 13690 15952
rect 13648 15910 13676 15943
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13740 15502 13768 16050
rect 13636 15496 13688 15502
rect 13634 15464 13636 15473
rect 13728 15496 13780 15502
rect 13688 15464 13690 15473
rect 13728 15438 13780 15444
rect 13634 15399 13690 15408
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14618 13768 14826
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13832 13938 13860 19858
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13924 18222 13952 18702
rect 14200 18630 14228 19246
rect 14292 18970 14320 19246
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13924 17082 13952 18158
rect 14016 17746 14044 18294
rect 14108 18222 14136 18566
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13924 17054 14044 17082
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 15706 13952 16934
rect 14016 16114 14044 17054
rect 14200 16998 14228 18022
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14016 15026 14044 16050
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14016 14618 14044 14962
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13820 13932 13872 13938
rect 13872 13892 13952 13920
rect 13820 13874 13872 13880
rect 13924 13410 13952 13892
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 13530 14044 13670
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13924 13382 14044 13410
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11082 13676 11494
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13740 10470 13768 11834
rect 13832 11762 13860 12650
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13924 11642 13952 12582
rect 14016 11898 14044 13382
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13832 11614 13952 11642
rect 14004 11620 14056 11626
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9382 13768 9998
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9110 13768 9318
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 6610 13676 8774
rect 13832 8378 13860 11614
rect 14004 11562 14056 11568
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13924 11286 13952 11494
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 14016 11121 14044 11562
rect 14002 11112 14058 11121
rect 14002 11047 14058 11056
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13924 8673 13952 10406
rect 14016 10198 14044 10406
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9722 14044 9998
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14108 9466 14136 16730
rect 14200 9586 14228 16934
rect 14292 16250 14320 18770
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14292 14362 14320 16186
rect 14384 14550 14412 19858
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14292 14334 14412 14362
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 11354 14320 13194
rect 14384 12646 14412 14334
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14292 9518 14320 11290
rect 14384 10606 14412 12106
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 9994 14412 10542
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14016 9438 14136 9466
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 13910 8664 13966 8673
rect 13910 8599 13966 8608
rect 13832 8350 13952 8378
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13818 7984 13874 7993
rect 13818 7919 13874 7928
rect 13832 7426 13860 7919
rect 13740 7410 13860 7426
rect 13728 7404 13860 7410
rect 13780 7398 13860 7404
rect 13728 7346 13780 7352
rect 13740 6882 13768 7346
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13832 7002 13860 7278
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13924 6934 13952 8350
rect 13912 6928 13964 6934
rect 13740 6854 13860 6882
rect 13912 6870 13964 6876
rect 13648 6582 13768 6610
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13372 3194 13400 3946
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12990 3088 13046 3097
rect 13188 3074 13216 3130
rect 13464 3074 13492 3606
rect 13188 3046 13492 3074
rect 12990 3023 13046 3032
rect 13004 2990 13032 3023
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13452 2508 13504 2514
rect 13556 2496 13584 5510
rect 13648 5166 13676 5646
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13504 2468 13584 2496
rect 13452 2450 13504 2456
rect 13636 2372 13688 2378
rect 13636 2314 13688 2320
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13096 480 13124 2246
rect 13648 480 13676 2314
rect 13740 649 13768 6582
rect 13832 4842 13860 6854
rect 14016 6254 14044 9438
rect 14096 9376 14148 9382
rect 14384 9364 14412 9454
rect 14096 9318 14148 9324
rect 14292 9336 14412 9364
rect 14108 9178 14136 9318
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14108 8430 14136 9114
rect 14186 8664 14242 8673
rect 14186 8599 14242 8608
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14200 8362 14228 8599
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14096 6928 14148 6934
rect 14094 6896 14096 6905
rect 14148 6896 14150 6905
rect 14094 6831 14150 6840
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13924 5574 13952 6054
rect 14016 5846 14044 6190
rect 14200 5914 14228 6190
rect 14292 6118 14320 9336
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8498 14412 8774
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14384 7954 14412 8434
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14384 6798 14412 7890
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13832 4814 14044 4842
rect 14016 4690 14044 4814
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13832 2582 13860 4626
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 3058 13952 3538
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13726 640 13782 649
rect 13726 575 13782 584
rect 14200 480 14228 4422
rect 14476 4264 14504 19246
rect 14568 18970 14596 20318
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15304 19786 15332 22320
rect 15856 20058 15884 22320
rect 16408 20074 16436 22320
rect 16408 20058 16620 20074
rect 15844 20052 15896 20058
rect 16408 20052 16632 20058
rect 16408 20046 16580 20052
rect 15844 19994 15896 20000
rect 16580 19994 16632 20000
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15580 19310 15608 19858
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15028 16538 15056 18566
rect 15120 18290 15148 18702
rect 15396 18426 15424 18770
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15396 17785 15424 18362
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15474 17912 15530 17921
rect 15474 17847 15476 17856
rect 15528 17847 15530 17856
rect 15476 17818 15528 17824
rect 15382 17776 15438 17785
rect 15382 17711 15438 17720
rect 15672 17678 15700 18158
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15212 17134 15240 17546
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15304 16658 15332 17206
rect 15488 17134 15516 17614
rect 15672 17338 15700 17614
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15200 16584 15252 16590
rect 15028 16510 15148 16538
rect 15200 16526 15252 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 16182 15056 16390
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 15028 15978 15056 16118
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15028 15502 15056 15914
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14074 14596 14758
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12850 14688 13126
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 15120 12753 15148 16510
rect 15212 15858 15240 16526
rect 15304 16522 15332 16594
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15384 15904 15436 15910
rect 15212 15830 15332 15858
rect 15384 15846 15436 15852
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15212 14550 15240 15642
rect 15304 15026 15332 15830
rect 15396 15570 15424 15846
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15396 14958 15424 15506
rect 15488 15201 15516 16934
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 15473 15608 16594
rect 15764 16590 15792 19858
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15948 18970 15976 19450
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15856 18358 15884 18770
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 16040 16980 16068 18566
rect 16132 17882 16160 19110
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16224 17338 16252 19110
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16316 18426 16344 18634
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16302 17776 16358 17785
rect 16302 17711 16358 17720
rect 16316 17678 16344 17711
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16316 17202 16344 17614
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16304 16992 16356 16998
rect 16040 16952 16304 16980
rect 16304 16934 16356 16940
rect 16210 16824 16266 16833
rect 16210 16759 16266 16768
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15764 16114 15792 16390
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15706 15700 15846
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15856 15638 15884 16390
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15660 15496 15712 15502
rect 15566 15464 15622 15473
rect 16040 15484 16068 16594
rect 16224 16590 16252 16759
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16210 16144 16266 16153
rect 16210 16079 16266 16088
rect 15712 15456 16068 15484
rect 16120 15496 16172 15502
rect 15660 15438 15712 15444
rect 16120 15438 16172 15444
rect 15566 15399 15622 15408
rect 15474 15192 15530 15201
rect 15474 15127 15530 15136
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15212 13258 15240 14350
rect 15304 14074 15332 14758
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15304 13938 15332 14010
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15488 13546 15516 14962
rect 15396 13518 15516 13546
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15200 12912 15252 12918
rect 15198 12880 15200 12889
rect 15252 12880 15254 12889
rect 15198 12815 15254 12824
rect 15106 12744 15162 12753
rect 15106 12679 15162 12688
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14568 11558 14596 12242
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11762 14688 12038
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14568 10606 14596 11494
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15120 10826 15148 12679
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11801 15240 12038
rect 15198 11792 15254 11801
rect 15198 11727 15254 11736
rect 15396 11150 15424 13518
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15488 13297 15516 13330
rect 15474 13288 15530 13297
rect 15474 13223 15530 13232
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15028 10798 15148 10826
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15028 10266 15056 10798
rect 15304 10674 15332 10950
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15120 10266 15148 10610
rect 15488 10606 15516 12174
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 14568 6798 14596 10202
rect 14646 10160 14702 10169
rect 14646 10095 14702 10104
rect 14660 9518 14688 10095
rect 15120 10062 15148 10202
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14752 9450 14780 9998
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 15028 9738 15056 9930
rect 15028 9710 15148 9738
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 15028 9382 15056 9522
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14752 7410 14780 7890
rect 14922 7440 14978 7449
rect 14740 7404 14792 7410
rect 14922 7375 14978 7384
rect 14740 7346 14792 7352
rect 14936 7342 14964 7375
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 5914 14596 6598
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14384 4236 14504 4264
rect 14384 4146 14412 4236
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3194 14412 3878
rect 14568 3738 14596 4082
rect 15028 4078 15056 9318
rect 15120 7426 15148 9710
rect 15212 9110 15240 9998
rect 15304 9178 15332 10474
rect 15580 10418 15608 15399
rect 15658 15192 15714 15201
rect 15658 15127 15714 15136
rect 15672 14006 15700 15127
rect 16132 14618 16160 15438
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16132 14482 16160 14554
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15764 13870 15792 14350
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15672 13682 15700 13738
rect 15936 13728 15988 13734
rect 15934 13696 15936 13705
rect 15988 13696 15990 13705
rect 15672 13654 15884 13682
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 10810 15700 13330
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 11898 15792 13262
rect 15856 12646 15884 13654
rect 15934 13631 15990 13640
rect 16132 13530 16160 14010
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12986 15976 13262
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15948 12374 15976 12922
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 16040 11762 16068 12650
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15750 11520 15806 11529
rect 15750 11455 15806 11464
rect 15764 11354 15792 11455
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15580 10390 15700 10418
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15396 9722 15424 10066
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15580 9586 15608 10066
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15120 7398 15240 7426
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15120 6186 15148 7210
rect 15212 7002 15240 7398
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15396 6730 15424 8230
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15304 6118 15332 6326
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 5166 15148 5646
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 15212 4826 15240 5714
rect 15304 4865 15332 6054
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15396 5166 15424 5782
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15290 4856 15346 4865
rect 15200 4820 15252 4826
rect 15290 4791 15346 4800
rect 15200 4762 15252 4768
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14372 3052 14424 3058
rect 14476 3040 14504 3538
rect 14424 3012 14504 3040
rect 14372 2994 14424 3000
rect 14568 2922 14596 3674
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15028 1442 15056 3878
rect 14752 1414 15056 1442
rect 14752 480 14780 1414
rect 15304 480 15332 4422
rect 15488 2990 15516 8230
rect 15580 6866 15608 8298
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15580 5409 15608 6666
rect 15566 5400 15622 5409
rect 15566 5335 15622 5344
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15580 3602 15608 5170
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15580 2514 15608 3130
rect 15672 2553 15700 10390
rect 15764 7970 15792 11290
rect 15856 11150 15884 11698
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15948 9382 15976 11494
rect 16040 10674 16068 11698
rect 16132 11626 16160 13466
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16224 11286 16252 16079
rect 16316 15994 16344 16934
rect 16408 16153 16436 19858
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16684 18970 16712 19314
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16500 17202 16528 18906
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16500 16697 16528 17138
rect 16486 16688 16542 16697
rect 16486 16623 16542 16632
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16394 16144 16450 16153
rect 16394 16079 16450 16088
rect 16500 16017 16528 16458
rect 16486 16008 16542 16017
rect 16316 15966 16436 15994
rect 16408 15026 16436 15966
rect 16486 15943 16542 15952
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 14657 16344 14758
rect 16302 14648 16358 14657
rect 16302 14583 16358 14592
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16316 12782 16344 13806
rect 16408 13530 16436 14826
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16316 12102 16344 12718
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11898 16344 12038
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16132 9382 16160 11018
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15948 9081 15976 9318
rect 16224 9178 16252 9522
rect 16408 9518 16436 12310
rect 16500 11694 16528 14894
rect 16592 14074 16620 18770
rect 16684 18154 16712 18906
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16776 17542 16804 19858
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16868 18630 16896 19246
rect 16960 18970 16988 22320
rect 17512 20058 17540 22320
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16868 17746 16896 18158
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16776 16017 16804 17206
rect 16762 16008 16818 16017
rect 16762 15943 16818 15952
rect 16868 15201 16896 17478
rect 16960 17338 16988 17750
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16960 16046 16988 16730
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 17052 15201 17080 19246
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17130 18184 17186 18193
rect 17130 18119 17186 18128
rect 17144 17542 17172 18119
rect 17236 17814 17264 19178
rect 17328 18834 17356 19926
rect 18064 19700 18092 22320
rect 18510 21176 18566 21185
rect 18510 21111 18566 21120
rect 18142 20632 18198 20641
rect 18142 20567 18198 20576
rect 18156 19786 18184 20567
rect 18524 20058 18552 21111
rect 18616 20058 18644 22320
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 17972 19672 18092 19700
rect 17972 18970 18000 19672
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17144 16794 17172 17002
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17328 16674 17356 18770
rect 18432 18714 18460 19246
rect 18616 19242 18644 19858
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18788 18760 18840 18766
rect 18432 18686 18736 18714
rect 18788 18702 18840 18708
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 17682 18320 17738 18329
rect 17682 18255 17738 18264
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 17134 17448 17478
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17144 16646 17356 16674
rect 17592 16652 17644 16658
rect 17144 15314 17172 16646
rect 17592 16594 17644 16600
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17328 16114 17356 16526
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17328 15706 17356 16050
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17408 15360 17460 15366
rect 17144 15286 17356 15314
rect 17408 15302 17460 15308
rect 16854 15192 16910 15201
rect 16854 15127 16910 15136
rect 17038 15192 17094 15201
rect 17038 15127 17094 15136
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16684 13530 16712 14758
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16592 11762 16620 13126
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16776 11370 16804 14418
rect 16868 12374 16896 14962
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16684 11342 16804 11370
rect 16684 10146 16712 11342
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16776 10266 16804 11154
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16684 10118 16804 10146
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16408 9194 16436 9454
rect 16212 9172 16264 9178
rect 16408 9166 16620 9194
rect 16212 9114 16264 9120
rect 15934 9072 15990 9081
rect 15934 9007 15990 9016
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16408 8498 16436 8978
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16132 8090 16160 8230
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 15764 7942 15976 7970
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7342 15792 7822
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15948 7154 15976 7942
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16040 7342 16068 7890
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15948 7126 16160 7154
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 4078 15792 6054
rect 15856 5846 15884 6734
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15856 5370 15884 5782
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15856 5250 15884 5306
rect 15856 5222 15976 5250
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15658 2544 15714 2553
rect 15568 2508 15620 2514
rect 15658 2479 15714 2488
rect 15568 2450 15620 2456
rect 15672 2446 15700 2479
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15856 480 15884 4966
rect 15948 4622 15976 5222
rect 16040 5098 16068 6802
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16132 3738 16160 7126
rect 16224 7002 16252 8230
rect 16408 7954 16436 8230
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16500 6866 16528 8570
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16132 3126 16160 3538
rect 16224 3194 16252 6734
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16132 2446 16160 3062
rect 16316 2446 16344 5578
rect 16500 5166 16528 5850
rect 16592 5642 16620 9166
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16684 6662 16712 7482
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 5710 16712 6598
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16776 4758 16804 10118
rect 16868 9518 16896 11494
rect 17052 11354 17080 15030
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17144 12986 17172 14758
rect 17236 14550 17264 14962
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17236 14074 17264 14486
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17222 13832 17278 13841
rect 17222 13767 17278 13776
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17236 12866 17264 13767
rect 17144 12838 17264 12866
rect 17144 11642 17172 12838
rect 17222 12744 17278 12753
rect 17222 12679 17224 12688
rect 17276 12679 17278 12688
rect 17224 12650 17276 12656
rect 17328 12322 17356 15286
rect 17420 14346 17448 15302
rect 17512 14618 17540 15506
rect 17604 15366 17632 16594
rect 17696 16590 17724 18255
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17696 14958 17724 15982
rect 17788 15502 17816 18566
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18524 18222 18552 18566
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18524 17882 18552 18022
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18616 17610 18644 18226
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16810 17908 17070
rect 17960 16992 18012 16998
rect 17958 16960 17960 16969
rect 18012 16960 18014 16969
rect 17958 16895 18014 16904
rect 17880 16782 18000 16810
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17512 13326 17540 14554
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17604 13002 17632 14554
rect 17788 14482 17816 15438
rect 17880 15162 17908 16594
rect 17972 16046 18000 16782
rect 18064 16561 18092 17206
rect 18616 17134 18644 17546
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18050 16552 18106 16561
rect 18050 16487 18106 16496
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17972 15910 18000 15982
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17972 15638 18000 15846
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 18524 14618 18552 16594
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 14890 18644 16390
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17420 12974 17632 13002
rect 17420 12646 17448 12974
rect 17498 12744 17554 12753
rect 17498 12679 17554 12688
rect 17408 12640 17460 12646
rect 17406 12608 17408 12617
rect 17460 12608 17462 12617
rect 17406 12543 17462 12552
rect 17328 12294 17448 12322
rect 17420 12238 17448 12294
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11762 17356 12038
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17144 11614 17264 11642
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10606 17080 10950
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 17052 9110 17080 10542
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17052 8906 17080 9046
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 17144 8498 17172 11494
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16868 7546 16896 8434
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 17236 6866 17264 11614
rect 17328 11286 17356 11698
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17420 11098 17448 12174
rect 17512 11626 17540 12679
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17604 11354 17632 11766
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17696 11234 17724 13670
rect 17788 13530 17816 14214
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17880 13258 17908 14350
rect 17972 14074 18000 14418
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18234 13832 18290 13841
rect 18234 13767 18290 13776
rect 18248 13530 18276 13767
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18142 13424 18198 13433
rect 18524 13394 18552 14282
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18616 13802 18644 13874
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18142 13359 18144 13368
rect 18196 13359 18198 13368
rect 18512 13388 18564 13394
rect 18144 13330 18196 13336
rect 18512 13330 18564 13336
rect 18616 13326 18644 13738
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18616 12782 18644 13262
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 17866 12336 17922 12345
rect 17866 12271 17868 12280
rect 17920 12271 17922 12280
rect 17868 12242 17920 12248
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17328 11070 17448 11098
rect 17512 11206 17724 11234
rect 17328 7834 17356 11070
rect 17512 10962 17540 11206
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17420 10934 17540 10962
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17420 10198 17448 10934
rect 17604 10554 17632 10950
rect 17512 10538 17632 10554
rect 17500 10532 17632 10538
rect 17552 10526 17632 10532
rect 17500 10474 17552 10480
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9722 17448 9998
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17512 9586 17540 10474
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17604 10062 17632 10406
rect 17696 10266 17724 11018
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17604 9450 17632 9998
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17420 7954 17448 8434
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17328 7806 17448 7834
rect 17314 7712 17370 7721
rect 17314 7647 17370 7656
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 16854 6216 16910 6225
rect 16854 6151 16856 6160
rect 16908 6151 16910 6160
rect 16856 6122 16908 6128
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16946 5672 17002 5681
rect 16946 5607 17002 5616
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16408 480 16436 3878
rect 16592 2514 16620 4626
rect 16960 3194 16988 5607
rect 17052 4826 17080 6054
rect 17144 5846 17172 6258
rect 17236 5914 17264 6258
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17144 5370 17172 5782
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17236 5234 17264 5646
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17328 4146 17356 7647
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17144 3058 17172 3606
rect 17236 3602 17264 3946
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17420 3505 17448 7806
rect 17512 5817 17540 9318
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17604 8634 17632 8978
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 6798 17632 7686
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17498 5808 17554 5817
rect 17498 5743 17554 5752
rect 17696 5692 17724 10066
rect 17788 9518 17816 11494
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17880 9178 17908 10542
rect 17972 10266 18000 12718
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 12238 18644 12582
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18616 11898 18644 12174
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18050 10704 18106 10713
rect 18050 10639 18106 10648
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 9976 18092 10639
rect 18524 10198 18552 10950
rect 18616 10554 18644 11562
rect 18708 11370 18736 18686
rect 18800 18426 18828 18702
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18800 17746 18828 18362
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18800 17610 18828 17682
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 18892 16946 18920 19858
rect 18984 19242 19012 22471
rect 19154 22320 19210 22800
rect 19706 22320 19762 22800
rect 20258 22320 20314 22800
rect 20810 22320 20866 22800
rect 21362 22320 21418 22800
rect 21914 22320 21970 22800
rect 22466 22320 22522 22800
rect 19062 21584 19118 21593
rect 19062 21519 19118 21528
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 19076 19174 19104 21519
rect 19168 20618 19196 22320
rect 19168 20590 19380 20618
rect 19352 20058 19380 20590
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19248 19848 19300 19854
rect 19154 19816 19210 19825
rect 19248 19790 19300 19796
rect 19154 19751 19210 19760
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19168 18850 19196 19751
rect 19260 19689 19288 19790
rect 19246 19680 19302 19689
rect 19246 19615 19302 19624
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19076 18822 19196 18850
rect 18970 18184 19026 18193
rect 18970 18119 19026 18128
rect 18984 17882 19012 18119
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18892 16918 19012 16946
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18800 15638 18828 15846
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18800 15026 18828 15574
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18892 14958 18920 16730
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18800 13190 18828 13806
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18892 12306 18920 14758
rect 18984 12986 19012 16918
rect 19076 16130 19104 18822
rect 19154 18728 19210 18737
rect 19154 18663 19210 18672
rect 19168 18426 19196 18663
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19260 18329 19288 18566
rect 19246 18320 19302 18329
rect 19246 18255 19302 18264
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19168 16833 19196 17682
rect 19352 17338 19380 19110
rect 19444 17921 19472 19858
rect 19720 18986 19748 22320
rect 20166 20224 20222 20233
rect 20166 20159 20222 20168
rect 20180 20058 20208 20159
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19628 18958 19748 18986
rect 19628 18698 19656 18958
rect 19706 18864 19762 18873
rect 19706 18799 19708 18808
rect 19760 18799 19762 18808
rect 19708 18770 19760 18776
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 19430 17912 19486 17921
rect 19430 17847 19486 17856
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19154 16824 19210 16833
rect 19154 16759 19210 16768
rect 19352 16590 19380 16934
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19076 16102 19288 16130
rect 19062 15056 19118 15065
rect 19062 14991 19118 15000
rect 19076 13530 19104 14991
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19076 12986 19104 13262
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19168 12646 19196 14418
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 18892 11830 18920 12242
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 18708 11342 18828 11370
rect 18800 11234 18828 11342
rect 18696 11212 18748 11218
rect 18800 11206 18920 11234
rect 18696 11154 18748 11160
rect 18708 10674 18736 11154
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18616 10526 18736 10554
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18616 10266 18644 10406
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 17972 9948 18092 9976
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17866 8392 17922 8401
rect 17866 8327 17868 8336
rect 17920 8327 17922 8336
rect 17868 8298 17920 8304
rect 17512 5664 17724 5692
rect 17406 3496 17462 3505
rect 17406 3431 17462 3440
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16776 2582 16804 2790
rect 16960 2650 16988 2790
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17512 2582 17540 5664
rect 17880 5352 17908 8298
rect 17972 6186 18000 9948
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18052 9512 18104 9518
rect 18708 9489 18736 10526
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18800 10062 18828 10474
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18052 9454 18104 9460
rect 18694 9480 18750 9489
rect 18064 8906 18092 9454
rect 18694 9415 18750 9424
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18708 8242 18736 9415
rect 18708 8214 18828 8242
rect 18694 8120 18750 8129
rect 18694 8055 18750 8064
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18510 7576 18566 7585
rect 18510 7511 18566 7520
rect 18234 7304 18290 7313
rect 18234 7239 18290 7248
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 7002 18092 7142
rect 18248 7002 18276 7239
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18524 6934 18552 7511
rect 18616 7410 18644 7890
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 18616 6798 18644 7346
rect 18708 7274 18736 8055
rect 18800 7342 18828 8214
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17696 5324 17908 5352
rect 17696 4078 17724 5324
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4554 17816 4966
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17604 2990 17632 3334
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17788 2514 17816 4490
rect 17880 4078 17908 5170
rect 17972 4758 18000 5714
rect 18524 5710 18552 6190
rect 18616 5914 18644 6734
rect 18800 6225 18828 7142
rect 18786 6216 18842 6225
rect 18786 6151 18842 6160
rect 18696 6112 18748 6118
rect 18892 6066 18920 11206
rect 19076 10690 19104 11494
rect 19168 10810 19196 12242
rect 19260 12102 19288 16102
rect 19352 15978 19380 16526
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19444 15706 19472 16594
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19536 14634 19564 17002
rect 19628 14822 19656 17138
rect 19812 15994 19840 19178
rect 19996 18902 20024 19858
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19904 16794 19932 17070
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19720 15966 19840 15994
rect 19720 15094 19748 15966
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19708 15088 19760 15094
rect 19708 15030 19760 15036
rect 19812 15026 19840 15846
rect 19904 15706 19932 16050
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19904 15094 19932 15642
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19996 14906 20024 16934
rect 20088 15162 20116 18158
rect 20180 15978 20208 19858
rect 20272 18834 20300 22320
rect 20626 22128 20682 22137
rect 20626 22063 20682 22072
rect 20640 20058 20668 22063
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20626 19272 20682 19281
rect 20626 19207 20682 19216
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20442 17912 20498 17921
rect 20442 17847 20498 17856
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20260 16720 20312 16726
rect 20260 16662 20312 16668
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20180 15366 20208 15914
rect 20272 15570 20300 16662
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19904 14878 20024 14906
rect 20074 14920 20130 14929
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19536 14606 19656 14634
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19430 14104 19486 14113
rect 19430 14039 19486 14048
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19352 13462 19380 13738
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19352 11762 19380 12582
rect 19444 11898 19472 14039
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19076 10662 19196 10690
rect 19260 10674 19288 11018
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18984 9926 19012 10406
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 19076 9738 19104 10406
rect 18984 9710 19104 9738
rect 18984 6322 19012 9710
rect 19168 9602 19196 10662
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19260 10130 19288 10610
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19352 10198 19380 10542
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19076 9574 19196 9602
rect 19076 7206 19104 9574
rect 19352 9518 19380 10134
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19352 9042 19380 9454
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9110 19472 9318
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8090 19380 8978
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19246 7168 19302 7177
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 19076 6254 19104 6734
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 18696 6054 18748 6060
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18524 5234 18552 5646
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17880 3074 17908 3878
rect 17972 3194 18000 4558
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18616 4321 18644 5034
rect 18708 4758 18736 6054
rect 18800 6038 18920 6066
rect 18800 4826 18828 6038
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18602 4312 18658 4321
rect 18602 4247 18658 4256
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18616 3738 18644 3946
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17880 3046 18000 3074
rect 18616 3058 18644 3674
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 16960 480 16988 2246
rect 17512 480 17540 2246
rect 17972 1442 18000 3046
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18708 2961 18736 4014
rect 18984 3505 19012 5850
rect 19168 4826 19196 7142
rect 19246 7103 19302 7112
rect 19260 6118 19288 7103
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 4826 19288 6054
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19076 3602 19104 4422
rect 19168 3942 19196 4558
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19444 3602 19472 8502
rect 19536 5914 19564 14486
rect 19628 6458 19656 14606
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19708 13388 19760 13394
rect 19708 13330 19760 13336
rect 19720 12442 19748 13330
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19812 11286 19840 13738
rect 19904 13530 19932 14878
rect 20074 14855 20130 14864
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19996 14074 20024 14758
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 20088 13802 20116 14855
rect 20180 14550 20208 15302
rect 20364 15178 20392 16934
rect 20456 15706 20484 17847
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20272 15150 20392 15178
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20180 13870 20208 14350
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19890 12880 19946 12889
rect 19890 12815 19946 12824
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19720 8906 19748 10066
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19706 7440 19762 7449
rect 19706 7375 19762 7384
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19720 6338 19748 7375
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19628 6310 19748 6338
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19524 3528 19576 3534
rect 18970 3496 19026 3505
rect 19524 3470 19576 3476
rect 18970 3431 19026 3440
rect 18694 2952 18750 2961
rect 18694 2887 18696 2896
rect 18748 2887 18750 2896
rect 18696 2858 18748 2864
rect 18708 2827 18736 2858
rect 18418 2680 18474 2689
rect 18418 2615 18474 2624
rect 18432 2514 18460 2615
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18616 2009 18644 2518
rect 19536 2514 19564 3470
rect 19628 2990 19656 6310
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19720 4282 19748 4626
rect 19812 4622 19840 6802
rect 19904 6474 19932 12815
rect 19996 12714 20024 13262
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19996 12442 20024 12650
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19996 9178 20024 11154
rect 20088 10470 20116 11562
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20272 10418 20300 15150
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20364 14482 20392 15030
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20456 14618 20484 14962
rect 20548 14958 20576 18090
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20456 14521 20484 14554
rect 20442 14512 20498 14521
rect 20352 14476 20404 14482
rect 20442 14447 20498 14456
rect 20352 14418 20404 14424
rect 20364 13938 20392 14418
rect 20640 14074 20668 19207
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 18290 20760 18702
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20824 17490 20852 22320
rect 21376 19854 21404 22320
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21928 19174 21956 22320
rect 22480 20262 22508 22320
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20916 17882 20944 18906
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20732 17462 20852 17490
rect 20732 16454 20760 17462
rect 20810 17368 20866 17377
rect 20810 17303 20866 17312
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20456 12782 20484 13126
rect 20732 12850 20760 16186
rect 20824 15162 20852 17303
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20916 15502 20944 15914
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15609 21036 15846
rect 20994 15600 21050 15609
rect 20994 15535 21050 15544
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20824 11121 20852 13806
rect 20810 11112 20866 11121
rect 20810 11047 20866 11056
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20350 10432 20406 10441
rect 20272 10390 20350 10418
rect 20350 10367 20406 10376
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19996 8294 20024 8774
rect 20088 8430 20116 9318
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19996 6769 20024 8230
rect 20180 8090 20208 8434
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20364 7342 20392 10367
rect 20548 10266 20576 10474
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20534 10024 20590 10033
rect 20534 9959 20590 9968
rect 20548 9518 20576 9959
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 8090 20484 9318
rect 20548 9110 20576 9454
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20640 8498 20668 9522
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20640 8022 20668 8434
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19904 6446 20208 6474
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19904 5370 19932 6190
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19812 4078 19840 4422
rect 19904 4214 19932 5306
rect 19892 4208 19944 4214
rect 19892 4150 19944 4156
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19996 2990 20024 5510
rect 20180 5250 20208 6446
rect 20272 5914 20300 7142
rect 20456 6254 20484 7346
rect 20640 7002 20668 7958
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 6458 20668 6802
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20088 5222 20208 5250
rect 20088 5098 20116 5222
rect 20272 5166 20300 5510
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20260 5160 20312 5166
rect 20312 5108 20392 5114
rect 20260 5102 20392 5108
rect 20076 5092 20128 5098
rect 20272 5086 20392 5102
rect 20076 5034 20128 5040
rect 20364 4622 20392 5086
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20272 3913 20300 4558
rect 20456 4078 20484 5238
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20258 3904 20314 3913
rect 20258 3839 20314 3848
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 18602 2000 18658 2009
rect 18602 1935 18658 1944
rect 17972 1414 18092 1442
rect 18064 480 18092 1414
rect 18708 1170 18736 2314
rect 19064 2304 19116 2310
rect 19616 2304 19668 2310
rect 19116 2264 19196 2292
rect 19064 2246 19116 2252
rect 18616 1142 18736 1170
rect 18616 480 18644 1142
rect 19168 480 19196 2264
rect 19668 2264 19748 2292
rect 19616 2246 19668 2252
rect 19720 480 19748 2264
rect 20272 480 20300 3062
rect 20364 2514 20392 3470
rect 20548 2990 20576 4490
rect 20732 4078 20760 5034
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20824 480 20852 2246
rect 21376 480 21404 2858
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21928 480 21956 2790
rect 22480 480 22508 3878
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7470 0 7526 480
rect 8022 0 8078 480
rect 8574 0 8630 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10230 0 10286 480
rect 10782 0 10838 480
rect 11334 0 11390 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14186 0 14242 480
rect 14738 0 14794 480
rect 15290 0 15346 480
rect 15842 0 15898 480
rect 16394 0 16450 480
rect 16946 0 17002 480
rect 17498 0 17554 480
rect 18050 0 18106 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19706 0 19762 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
<< via2 >>
rect 18970 22480 19026 22536
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3422 17176 3478 17232
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 8482 19116 8484 19136
rect 8484 19116 8536 19136
rect 8536 19116 8538 19136
rect 8482 19080 8538 19116
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4066 5752 4122 5808
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 6366 3440 6422 3496
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 9770 19780 9826 19816
rect 9770 19760 9772 19780
rect 9772 19760 9824 19780
rect 9824 19760 9826 19780
rect 9678 18264 9734 18320
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 10322 18944 10378 19000
rect 10322 18808 10378 18864
rect 10506 18944 10562 19000
rect 10046 13912 10102 13968
rect 10138 13776 10194 13832
rect 10414 13912 10470 13968
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 10966 14864 11022 14920
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11610 14864 11666 14920
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 10414 9968 10470 10024
rect 10230 3068 10232 3088
rect 10232 3068 10284 3088
rect 10284 3068 10286 3088
rect 10230 3032 10286 3068
rect 10782 8336 10838 8392
rect 10874 1536 10930 1592
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11334 6860 11390 6896
rect 11334 6840 11336 6860
rect 11336 6840 11388 6860
rect 11388 6840 11390 6860
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 12346 18944 12402 19000
rect 12254 16496 12310 16552
rect 12438 16496 12494 16552
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12622 13912 12678 13968
rect 13082 18128 13138 18184
rect 12898 13368 12954 13424
rect 13266 14492 13268 14512
rect 13268 14492 13320 14512
rect 13320 14492 13322 14512
rect 13266 14456 13322 14492
rect 13266 11192 13322 11248
rect 12254 7384 12310 7440
rect 12162 1536 12218 1592
rect 13174 7964 13176 7984
rect 13176 7964 13228 7984
rect 13228 7964 13230 7984
rect 12714 6160 12770 6216
rect 13174 7928 13230 7964
rect 13634 15952 13690 16008
rect 13634 15444 13636 15464
rect 13636 15444 13688 15464
rect 13688 15444 13690 15464
rect 13634 15408 13690 15444
rect 14002 11056 14058 11112
rect 13910 8608 13966 8664
rect 13818 7928 13874 7984
rect 12990 3032 13046 3088
rect 14186 8608 14242 8664
rect 14094 6876 14096 6896
rect 14096 6876 14148 6896
rect 14148 6876 14150 6896
rect 14094 6840 14150 6876
rect 13726 584 13782 640
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 15474 17876 15530 17912
rect 15474 17856 15476 17876
rect 15476 17856 15528 17876
rect 15528 17856 15530 17876
rect 15382 17720 15438 17776
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 16302 17720 16358 17776
rect 16210 16768 16266 16824
rect 15566 15408 15622 15464
rect 16210 16088 16266 16144
rect 15474 15136 15530 15192
rect 15198 12860 15200 12880
rect 15200 12860 15252 12880
rect 15252 12860 15254 12880
rect 15198 12824 15254 12860
rect 15106 12688 15162 12744
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 15198 11736 15254 11792
rect 15474 13232 15530 13288
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14646 10104 14702 10160
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14922 7384 14978 7440
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 15658 15136 15714 15192
rect 15934 13676 15936 13696
rect 15936 13676 15988 13696
rect 15988 13676 15990 13696
rect 15934 13640 15990 13676
rect 15750 11464 15806 11520
rect 15290 4800 15346 4856
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15566 5344 15622 5400
rect 16486 16632 16542 16688
rect 16394 16088 16450 16144
rect 16486 15952 16542 16008
rect 16302 14592 16358 14648
rect 16762 15952 16818 16008
rect 17130 18128 17186 18184
rect 18510 21120 18566 21176
rect 18142 20576 18198 20632
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17682 18264 17738 18320
rect 16854 15136 16910 15192
rect 17038 15136 17094 15192
rect 15934 9016 15990 9072
rect 15658 2488 15714 2544
rect 17222 13776 17278 13832
rect 17222 12708 17278 12744
rect 17222 12688 17224 12708
rect 17224 12688 17276 12708
rect 17276 12688 17278 12708
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 16940 17960 16960
rect 17960 16940 18012 16960
rect 18012 16940 18014 16960
rect 17958 16904 18014 16940
rect 18050 16496 18106 16552
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 17498 12688 17554 12744
rect 17406 12588 17408 12608
rect 17408 12588 17460 12608
rect 17460 12588 17462 12608
rect 17406 12552 17462 12588
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18234 13776 18290 13832
rect 18142 13388 18198 13424
rect 18142 13368 18144 13388
rect 18144 13368 18196 13388
rect 18196 13368 18198 13388
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17866 12300 17922 12336
rect 17866 12280 17868 12300
rect 17868 12280 17920 12300
rect 17920 12280 17922 12300
rect 17314 7656 17370 7712
rect 16854 6180 16910 6216
rect 16854 6160 16856 6180
rect 16856 6160 16908 6180
rect 16908 6160 16910 6180
rect 16946 5616 17002 5672
rect 17498 5752 17554 5808
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18050 10648 18106 10704
rect 19062 21528 19118 21584
rect 19154 19760 19210 19816
rect 19246 19624 19302 19680
rect 18970 18128 19026 18184
rect 19154 18672 19210 18728
rect 19246 18264 19302 18320
rect 20166 20168 20222 20224
rect 19706 18828 19762 18864
rect 19706 18808 19708 18828
rect 19708 18808 19760 18828
rect 19760 18808 19762 18828
rect 19430 17856 19486 17912
rect 19154 16768 19210 16824
rect 19062 15000 19118 15056
rect 17866 8356 17922 8392
rect 17866 8336 17868 8356
rect 17868 8336 17920 8356
rect 17920 8336 17922 8356
rect 17406 3440 17462 3496
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18694 9424 18750 9480
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18694 8064 18750 8120
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18510 7520 18566 7576
rect 18234 7248 18290 7304
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18786 6160 18842 6216
rect 20626 22072 20682 22128
rect 20626 19216 20682 19272
rect 20442 17856 20498 17912
rect 19430 14048 19486 14104
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18602 4256 18658 4312
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 19246 7112 19302 7168
rect 20074 14864 20130 14920
rect 19890 12824 19946 12880
rect 19706 7384 19762 7440
rect 18970 3440 19026 3496
rect 18694 2916 18750 2952
rect 18694 2896 18696 2916
rect 18696 2896 18748 2916
rect 18748 2896 18750 2916
rect 18418 2624 18474 2680
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 20442 14456 20498 14512
rect 20810 17312 20866 17368
rect 20994 15544 21050 15600
rect 20810 11056 20866 11112
rect 20350 10376 20406 10432
rect 20534 9968 20590 10024
rect 19982 6704 20038 6760
rect 20258 3848 20314 3904
rect 18602 1944 18658 2000
<< metal3 >>
rect 18965 22538 19031 22541
rect 22320 22538 22800 22568
rect 18965 22536 22800 22538
rect 18965 22480 18970 22536
rect 19026 22480 22800 22536
rect 18965 22478 22800 22480
rect 18965 22475 19031 22478
rect 22320 22448 22800 22478
rect 20621 22130 20687 22133
rect 22320 22130 22800 22160
rect 20621 22128 22800 22130
rect 20621 22072 20626 22128
rect 20682 22072 22800 22128
rect 20621 22070 22800 22072
rect 20621 22067 20687 22070
rect 22320 22040 22800 22070
rect 19057 21586 19123 21589
rect 22320 21586 22800 21616
rect 19057 21584 22800 21586
rect 19057 21528 19062 21584
rect 19118 21528 22800 21584
rect 19057 21526 22800 21528
rect 19057 21523 19123 21526
rect 22320 21496 22800 21526
rect 18505 21178 18571 21181
rect 22320 21178 22800 21208
rect 18505 21176 22800 21178
rect 18505 21120 18510 21176
rect 18566 21120 22800 21176
rect 18505 21118 22800 21120
rect 18505 21115 18571 21118
rect 22320 21088 22800 21118
rect 18137 20634 18203 20637
rect 22320 20634 22800 20664
rect 18137 20632 22800 20634
rect 18137 20576 18142 20632
rect 18198 20576 22800 20632
rect 18137 20574 22800 20576
rect 18137 20571 18203 20574
rect 22320 20544 22800 20574
rect 20161 20226 20227 20229
rect 22320 20226 22800 20256
rect 20161 20224 22800 20226
rect 20161 20168 20166 20224
rect 20222 20168 22800 20224
rect 20161 20166 22800 20168
rect 20161 20163 20227 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 9765 19818 9831 19821
rect 19149 19818 19215 19821
rect 22320 19818 22800 19848
rect 9765 19816 18568 19818
rect 9765 19760 9770 19816
rect 9826 19760 18568 19816
rect 9765 19758 18568 19760
rect 9765 19755 9831 19758
rect 18508 19682 18568 19758
rect 19149 19816 22800 19818
rect 19149 19760 19154 19816
rect 19210 19760 22800 19816
rect 19149 19758 22800 19760
rect 19149 19755 19215 19758
rect 22320 19728 22800 19758
rect 19241 19682 19307 19685
rect 18508 19680 19307 19682
rect 18508 19624 19246 19680
rect 19302 19624 19307 19680
rect 18508 19622 19307 19624
rect 19241 19619 19307 19622
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 20621 19274 20687 19277
rect 22320 19274 22800 19304
rect 20621 19272 22800 19274
rect 20621 19216 20626 19272
rect 20682 19216 22800 19272
rect 20621 19214 22800 19216
rect 20621 19211 20687 19214
rect 22320 19184 22800 19214
rect 8477 19138 8543 19141
rect 10726 19138 10732 19140
rect 8477 19136 10732 19138
rect 8477 19080 8482 19136
rect 8538 19080 10732 19136
rect 8477 19078 10732 19080
rect 8477 19075 8543 19078
rect 10726 19076 10732 19078
rect 10796 19076 10802 19140
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 10317 19002 10383 19005
rect 10501 19002 10567 19005
rect 12341 19002 12407 19005
rect 10317 19000 12407 19002
rect 10317 18944 10322 19000
rect 10378 18944 10506 19000
rect 10562 18944 12346 19000
rect 12402 18944 12407 19000
rect 10317 18942 12407 18944
rect 10317 18939 10383 18942
rect 10501 18939 10567 18942
rect 12341 18939 12407 18942
rect 10317 18866 10383 18869
rect 19701 18866 19767 18869
rect 22320 18866 22800 18896
rect 10317 18864 19767 18866
rect 10317 18808 10322 18864
rect 10378 18808 19706 18864
rect 19762 18808 19767 18864
rect 10317 18806 19767 18808
rect 10317 18803 10383 18806
rect 19701 18803 19767 18806
rect 19934 18806 22800 18866
rect 19149 18730 19215 18733
rect 19934 18730 19994 18806
rect 22320 18776 22800 18806
rect 19149 18728 19994 18730
rect 19149 18672 19154 18728
rect 19210 18672 19994 18728
rect 19149 18670 19994 18672
rect 19149 18667 19215 18670
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 9673 18322 9739 18325
rect 14406 18322 14412 18324
rect 9673 18320 14412 18322
rect 9673 18264 9678 18320
rect 9734 18264 14412 18320
rect 9673 18262 14412 18264
rect 9673 18259 9739 18262
rect 14406 18260 14412 18262
rect 14476 18322 14482 18324
rect 17677 18322 17743 18325
rect 14476 18320 17743 18322
rect 14476 18264 17682 18320
rect 17738 18264 17743 18320
rect 14476 18262 17743 18264
rect 14476 18260 14482 18262
rect 17677 18259 17743 18262
rect 19241 18322 19307 18325
rect 22320 18322 22800 18352
rect 19241 18320 22800 18322
rect 19241 18264 19246 18320
rect 19302 18264 22800 18320
rect 19241 18262 22800 18264
rect 19241 18259 19307 18262
rect 22320 18232 22800 18262
rect 13077 18186 13143 18189
rect 17125 18186 17191 18189
rect 18965 18186 19031 18189
rect 13077 18184 19031 18186
rect 13077 18128 13082 18184
rect 13138 18128 17130 18184
rect 17186 18128 18970 18184
rect 19026 18128 19031 18184
rect 13077 18126 19031 18128
rect 13077 18123 13143 18126
rect 17125 18123 17191 18126
rect 18965 18123 19031 18126
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 15469 17914 15535 17917
rect 19425 17914 19491 17917
rect 15469 17912 19491 17914
rect 15469 17856 15474 17912
rect 15530 17856 19430 17912
rect 19486 17856 19491 17912
rect 15469 17854 19491 17856
rect 15469 17851 15535 17854
rect 19425 17851 19491 17854
rect 20437 17914 20503 17917
rect 22320 17914 22800 17944
rect 20437 17912 22800 17914
rect 20437 17856 20442 17912
rect 20498 17856 22800 17912
rect 20437 17854 22800 17856
rect 20437 17851 20503 17854
rect 22320 17824 22800 17854
rect 15377 17778 15443 17781
rect 16297 17778 16363 17781
rect 15377 17776 16363 17778
rect 15377 17720 15382 17776
rect 15438 17720 16302 17776
rect 16358 17720 16363 17776
rect 15377 17718 16363 17720
rect 15377 17715 15443 17718
rect 16297 17715 16363 17718
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 20805 17370 20871 17373
rect 22320 17370 22800 17400
rect 20805 17368 22800 17370
rect 20805 17312 20810 17368
rect 20866 17312 22800 17368
rect 20805 17310 22800 17312
rect 20805 17307 20871 17310
rect 22320 17280 22800 17310
rect 0 17234 480 17264
rect 3417 17234 3483 17237
rect 0 17232 3483 17234
rect 0 17176 3422 17232
rect 3478 17176 3483 17232
rect 0 17174 3483 17176
rect 0 17144 480 17174
rect 3417 17171 3483 17174
rect 17953 16962 18019 16965
rect 22320 16962 22800 16992
rect 17953 16960 22800 16962
rect 17953 16904 17958 16960
rect 18014 16904 22800 16960
rect 17953 16902 22800 16904
rect 17953 16899 18019 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 16205 16826 16271 16829
rect 19149 16826 19215 16829
rect 16205 16824 19215 16826
rect 16205 16768 16210 16824
rect 16266 16768 19154 16824
rect 19210 16768 19215 16824
rect 16205 16766 19215 16768
rect 16205 16763 16271 16766
rect 19149 16763 19215 16766
rect 16481 16692 16547 16693
rect 16430 16690 16436 16692
rect 16390 16630 16436 16690
rect 16500 16688 16547 16692
rect 16542 16632 16547 16688
rect 16430 16628 16436 16630
rect 16500 16628 16547 16632
rect 16481 16627 16547 16628
rect 12249 16554 12315 16557
rect 12433 16554 12499 16557
rect 12249 16552 12499 16554
rect 12249 16496 12254 16552
rect 12310 16496 12438 16552
rect 12494 16496 12499 16552
rect 12249 16494 12499 16496
rect 12249 16491 12315 16494
rect 12433 16491 12499 16494
rect 18045 16554 18111 16557
rect 22320 16554 22800 16584
rect 18045 16552 22800 16554
rect 18045 16496 18050 16552
rect 18106 16496 22800 16552
rect 18045 16494 22800 16496
rect 18045 16491 18111 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 16205 16146 16271 16149
rect 16389 16146 16455 16149
rect 16205 16144 16455 16146
rect 16205 16088 16210 16144
rect 16266 16088 16394 16144
rect 16450 16088 16455 16144
rect 16205 16086 16455 16088
rect 16205 16083 16271 16086
rect 16389 16083 16455 16086
rect 13629 16010 13695 16013
rect 16481 16010 16547 16013
rect 13629 16008 16547 16010
rect 13629 15952 13634 16008
rect 13690 15952 16486 16008
rect 16542 15952 16547 16008
rect 13629 15950 16547 15952
rect 13629 15947 13695 15950
rect 16481 15947 16547 15950
rect 16757 16010 16823 16013
rect 22320 16010 22800 16040
rect 16757 16008 22800 16010
rect 16757 15952 16762 16008
rect 16818 15952 22800 16008
rect 16757 15950 22800 15952
rect 16757 15947 16823 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 20989 15602 21055 15605
rect 22320 15602 22800 15632
rect 20989 15600 22800 15602
rect 20989 15544 20994 15600
rect 21050 15544 22800 15600
rect 20989 15542 22800 15544
rect 20989 15539 21055 15542
rect 22320 15512 22800 15542
rect 13629 15466 13695 15469
rect 15561 15466 15627 15469
rect 13629 15464 15627 15466
rect 13629 15408 13634 15464
rect 13690 15408 15566 15464
rect 15622 15408 15627 15464
rect 13629 15406 15627 15408
rect 13629 15403 13695 15406
rect 15561 15403 15627 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 15469 15194 15535 15197
rect 15653 15194 15719 15197
rect 16849 15196 16915 15197
rect 15469 15192 15719 15194
rect 15469 15136 15474 15192
rect 15530 15136 15658 15192
rect 15714 15136 15719 15192
rect 15469 15134 15719 15136
rect 15469 15131 15535 15134
rect 15653 15131 15719 15134
rect 16798 15132 16804 15196
rect 16868 15194 16915 15196
rect 17033 15194 17099 15197
rect 16868 15192 16960 15194
rect 16910 15136 16960 15192
rect 16868 15134 16960 15136
rect 17033 15192 17234 15194
rect 17033 15136 17038 15192
rect 17094 15136 17234 15192
rect 17033 15134 17234 15136
rect 16868 15132 16915 15134
rect 16849 15131 16915 15132
rect 17033 15131 17099 15134
rect 16982 14996 16988 15060
rect 17052 15058 17058 15060
rect 17174 15058 17234 15134
rect 17052 14998 17234 15058
rect 19057 15058 19123 15061
rect 22320 15058 22800 15088
rect 19057 15056 22800 15058
rect 19057 15000 19062 15056
rect 19118 15000 22800 15056
rect 19057 14998 22800 15000
rect 17052 14996 17058 14998
rect 19057 14995 19123 14998
rect 22320 14968 22800 14998
rect 10726 14860 10732 14924
rect 10796 14922 10802 14924
rect 10961 14922 11027 14925
rect 10796 14920 11027 14922
rect 10796 14864 10966 14920
rect 11022 14864 11027 14920
rect 10796 14862 11027 14864
rect 10796 14860 10802 14862
rect 10961 14859 11027 14862
rect 11605 14922 11671 14925
rect 20069 14922 20135 14925
rect 11605 14920 20135 14922
rect 11605 14864 11610 14920
rect 11666 14864 20074 14920
rect 20130 14864 20135 14920
rect 11605 14862 20135 14864
rect 11605 14859 11671 14862
rect 20069 14859 20135 14862
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 16297 14650 16363 14653
rect 22320 14650 22800 14680
rect 16297 14648 22800 14650
rect 16297 14592 16302 14648
rect 16358 14592 22800 14648
rect 16297 14590 22800 14592
rect 16297 14587 16363 14590
rect 22320 14560 22800 14590
rect 13261 14514 13327 14517
rect 20437 14514 20503 14517
rect 13261 14512 20503 14514
rect 13261 14456 13266 14512
rect 13322 14456 20442 14512
rect 20498 14456 20503 14512
rect 13261 14454 20503 14456
rect 13261 14451 13327 14454
rect 20437 14451 20503 14454
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 19425 14106 19491 14109
rect 22320 14106 22800 14136
rect 19425 14104 22800 14106
rect 19425 14048 19430 14104
rect 19486 14048 22800 14104
rect 19425 14046 22800 14048
rect 19425 14043 19491 14046
rect 22320 14016 22800 14046
rect 10041 13970 10107 13973
rect 10409 13970 10475 13973
rect 12617 13970 12683 13973
rect 10041 13968 12683 13970
rect 10041 13912 10046 13968
rect 10102 13912 10414 13968
rect 10470 13912 12622 13968
rect 12678 13912 12683 13968
rect 10041 13910 12683 13912
rect 10041 13907 10107 13910
rect 10409 13907 10475 13910
rect 12617 13907 12683 13910
rect 10133 13834 10199 13837
rect 17217 13834 17283 13837
rect 18229 13834 18295 13837
rect 10133 13832 18295 13834
rect 10133 13776 10138 13832
rect 10194 13776 17222 13832
rect 17278 13776 18234 13832
rect 18290 13776 18295 13832
rect 10133 13774 18295 13776
rect 10133 13771 10199 13774
rect 17217 13771 17283 13774
rect 18229 13771 18295 13774
rect 15929 13698 15995 13701
rect 22320 13698 22800 13728
rect 15929 13696 22800 13698
rect 15929 13640 15934 13696
rect 15990 13640 22800 13696
rect 15929 13638 22800 13640
rect 15929 13635 15995 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 12893 13426 12959 13429
rect 18137 13426 18203 13429
rect 18822 13426 18828 13428
rect 12893 13424 18828 13426
rect 12893 13368 12898 13424
rect 12954 13368 18142 13424
rect 18198 13368 18828 13424
rect 12893 13366 18828 13368
rect 12893 13363 12959 13366
rect 18137 13363 18203 13366
rect 18822 13364 18828 13366
rect 18892 13364 18898 13428
rect 15469 13290 15535 13293
rect 22320 13290 22800 13320
rect 15469 13288 22800 13290
rect 15469 13232 15474 13288
rect 15530 13232 22800 13288
rect 15469 13230 22800 13232
rect 15469 13227 15535 13230
rect 22320 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 15193 12882 15259 12885
rect 19885 12882 19951 12885
rect 15193 12880 19951 12882
rect 15193 12824 15198 12880
rect 15254 12824 19890 12880
rect 19946 12824 19951 12880
rect 15193 12822 19951 12824
rect 15193 12819 15259 12822
rect 19885 12819 19951 12822
rect 15101 12746 15167 12749
rect 17217 12746 17283 12749
rect 15101 12744 17283 12746
rect 15101 12688 15106 12744
rect 15162 12688 17222 12744
rect 17278 12688 17283 12744
rect 15101 12686 17283 12688
rect 15101 12683 15167 12686
rect 17217 12683 17283 12686
rect 17493 12746 17559 12749
rect 22320 12746 22800 12776
rect 17493 12744 22800 12746
rect 17493 12688 17498 12744
rect 17554 12688 22800 12744
rect 17493 12686 22800 12688
rect 17493 12683 17559 12686
rect 22320 12656 22800 12686
rect 17401 12612 17467 12613
rect 17350 12548 17356 12612
rect 17420 12610 17467 12612
rect 17420 12608 17512 12610
rect 17462 12552 17512 12608
rect 17420 12550 17512 12552
rect 17420 12548 17467 12550
rect 17401 12547 17467 12548
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 17861 12338 17927 12341
rect 22320 12338 22800 12368
rect 17861 12336 22800 12338
rect 17861 12280 17866 12336
rect 17922 12280 22800 12336
rect 17861 12278 22800 12280
rect 17861 12275 17927 12278
rect 22320 12248 22800 12278
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 15193 11794 15259 11797
rect 22320 11794 22800 11824
rect 15193 11792 22800 11794
rect 15193 11736 15198 11792
rect 15254 11736 22800 11792
rect 15193 11734 22800 11736
rect 15193 11731 15259 11734
rect 22320 11704 22800 11734
rect 15745 11522 15811 11525
rect 16430 11522 16436 11524
rect 15745 11520 16436 11522
rect 15745 11464 15750 11520
rect 15806 11464 16436 11520
rect 15745 11462 16436 11464
rect 15745 11459 15811 11462
rect 16430 11460 16436 11462
rect 16500 11460 16506 11524
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 22320 11386 22800 11416
rect 15702 11326 22800 11386
rect 13261 11250 13327 11253
rect 15702 11250 15762 11326
rect 22320 11296 22800 11326
rect 13261 11248 15762 11250
rect 13261 11192 13266 11248
rect 13322 11192 15762 11248
rect 13261 11190 15762 11192
rect 13261 11187 13327 11190
rect 13997 11114 14063 11117
rect 20805 11114 20871 11117
rect 13997 11112 20871 11114
rect 13997 11056 14002 11112
rect 14058 11056 20810 11112
rect 20866 11056 20871 11112
rect 13997 11054 20871 11056
rect 13997 11051 14063 11054
rect 20805 11051 20871 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 22320 10842 22800 10872
rect 18646 10782 22800 10842
rect 18045 10706 18111 10709
rect 18646 10706 18706 10782
rect 22320 10752 22800 10782
rect 18045 10704 18706 10706
rect 18045 10648 18050 10704
rect 18106 10648 18706 10704
rect 18045 10646 18706 10648
rect 18045 10643 18111 10646
rect 20345 10434 20411 10437
rect 22320 10434 22800 10464
rect 20345 10432 22800 10434
rect 20345 10376 20350 10432
rect 20406 10376 22800 10432
rect 20345 10374 22800 10376
rect 20345 10371 20411 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 14406 10100 14412 10164
rect 14476 10162 14482 10164
rect 14641 10162 14707 10165
rect 14476 10160 14707 10162
rect 14476 10104 14646 10160
rect 14702 10104 14707 10160
rect 14476 10102 14707 10104
rect 14476 10100 14482 10102
rect 14641 10099 14707 10102
rect 10409 10026 10475 10029
rect 16430 10026 16436 10028
rect 10409 10024 16436 10026
rect 10409 9968 10414 10024
rect 10470 9968 16436 10024
rect 10409 9966 16436 9968
rect 10409 9963 10475 9966
rect 16430 9964 16436 9966
rect 16500 9964 16506 10028
rect 20529 10026 20595 10029
rect 22320 10026 22800 10056
rect 20529 10024 22800 10026
rect 20529 9968 20534 10024
rect 20590 9968 22800 10024
rect 20529 9966 22800 9968
rect 20529 9963 20595 9966
rect 22320 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 18689 9482 18755 9485
rect 22320 9482 22800 9512
rect 18689 9480 22800 9482
rect 18689 9424 18694 9480
rect 18750 9424 22800 9480
rect 18689 9422 22800 9424
rect 18689 9419 18755 9422
rect 22320 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 15929 9074 15995 9077
rect 22320 9074 22800 9104
rect 15929 9072 22800 9074
rect 15929 9016 15934 9072
rect 15990 9016 22800 9072
rect 15929 9014 22800 9016
rect 15929 9011 15995 9014
rect 22320 8984 22800 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 13905 8666 13971 8669
rect 14181 8666 14247 8669
rect 13905 8664 17970 8666
rect 13905 8608 13910 8664
rect 13966 8608 14186 8664
rect 14242 8608 17970 8664
rect 13905 8606 17970 8608
rect 13905 8603 13971 8606
rect 14181 8603 14247 8606
rect 17910 8530 17970 8606
rect 22320 8530 22800 8560
rect 17910 8470 22800 8530
rect 22320 8440 22800 8470
rect 10777 8394 10843 8397
rect 17861 8394 17927 8397
rect 10777 8392 17927 8394
rect 10777 8336 10782 8392
rect 10838 8336 17866 8392
rect 17922 8336 17927 8392
rect 10777 8334 17927 8336
rect 10777 8331 10843 8334
rect 17861 8331 17927 8334
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 18689 8122 18755 8125
rect 22320 8122 22800 8152
rect 18689 8120 22800 8122
rect 18689 8064 18694 8120
rect 18750 8064 22800 8120
rect 18689 8062 22800 8064
rect 18689 8059 18755 8062
rect 22320 8032 22800 8062
rect 13169 7986 13235 7989
rect 13813 7986 13879 7989
rect 13169 7984 13879 7986
rect 13169 7928 13174 7984
rect 13230 7928 13818 7984
rect 13874 7928 13879 7984
rect 13169 7926 13879 7928
rect 13169 7923 13235 7926
rect 13813 7923 13879 7926
rect 17309 7716 17375 7717
rect 17309 7712 17356 7716
rect 17420 7714 17426 7716
rect 17309 7656 17314 7712
rect 17309 7652 17356 7656
rect 17420 7654 17466 7714
rect 17420 7652 17426 7654
rect 17309 7651 17375 7652
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 18505 7578 18571 7581
rect 22320 7578 22800 7608
rect 18505 7576 22800 7578
rect 18505 7520 18510 7576
rect 18566 7520 22800 7576
rect 18505 7518 22800 7520
rect 18505 7515 18571 7518
rect 22320 7488 22800 7518
rect 12249 7440 12315 7445
rect 12249 7384 12254 7440
rect 12310 7384 12315 7440
rect 12249 7379 12315 7384
rect 14917 7442 14983 7445
rect 16798 7442 16804 7444
rect 14917 7440 16804 7442
rect 14917 7384 14922 7440
rect 14978 7384 16804 7440
rect 14917 7382 16804 7384
rect 14917 7379 14983 7382
rect 16798 7380 16804 7382
rect 16868 7442 16874 7444
rect 19701 7442 19767 7445
rect 16868 7440 19767 7442
rect 16868 7384 19706 7440
rect 19762 7384 19767 7440
rect 16868 7382 19767 7384
rect 16868 7380 16874 7382
rect 19701 7379 19767 7382
rect 12252 7306 12312 7379
rect 17902 7306 17908 7308
rect 12252 7246 17908 7306
rect 17902 7244 17908 7246
rect 17972 7306 17978 7308
rect 18229 7306 18295 7309
rect 17972 7304 18295 7306
rect 17972 7248 18234 7304
rect 18290 7248 18295 7304
rect 17972 7246 18295 7248
rect 17972 7244 17978 7246
rect 18229 7243 18295 7246
rect 19241 7170 19307 7173
rect 22320 7170 22800 7200
rect 19241 7168 22800 7170
rect 19241 7112 19246 7168
rect 19302 7112 22800 7168
rect 19241 7110 22800 7112
rect 19241 7107 19307 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 11329 6898 11395 6901
rect 14089 6898 14155 6901
rect 11329 6896 14155 6898
rect 11329 6840 11334 6896
rect 11390 6840 14094 6896
rect 14150 6840 14155 6896
rect 11329 6838 14155 6840
rect 11329 6835 11395 6838
rect 14089 6835 14155 6838
rect 19977 6762 20043 6765
rect 22320 6762 22800 6792
rect 19977 6760 22800 6762
rect 19977 6704 19982 6760
rect 20038 6704 22800 6760
rect 19977 6702 22800 6704
rect 19977 6699 20043 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 12709 6218 12775 6221
rect 16849 6218 16915 6221
rect 12709 6216 16915 6218
rect 12709 6160 12714 6216
rect 12770 6160 16854 6216
rect 16910 6160 16915 6216
rect 12709 6158 16915 6160
rect 12709 6155 12775 6158
rect 16849 6155 16915 6158
rect 18781 6218 18847 6221
rect 22320 6218 22800 6248
rect 18781 6216 22800 6218
rect 18781 6160 18786 6216
rect 18842 6160 22800 6216
rect 18781 6158 22800 6160
rect 18781 6155 18847 6158
rect 22320 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 17493 5810 17559 5813
rect 22320 5810 22800 5840
rect 17493 5808 22800 5810
rect 17493 5752 17498 5808
rect 17554 5752 22800 5808
rect 17493 5750 22800 5752
rect 17493 5747 17559 5750
rect 22320 5720 22800 5750
rect 16941 5676 17007 5677
rect 16941 5674 16988 5676
rect 16896 5672 16988 5674
rect 16896 5616 16946 5672
rect 16896 5614 16988 5616
rect 16941 5612 16988 5614
rect 17052 5612 17058 5676
rect 16941 5611 17007 5612
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 15561 5402 15627 5405
rect 15561 5400 17970 5402
rect 15561 5344 15566 5400
rect 15622 5344 17970 5400
rect 15561 5342 17970 5344
rect 15561 5339 15627 5342
rect 17910 5266 17970 5342
rect 22320 5266 22800 5296
rect 17910 5206 22800 5266
rect 22320 5176 22800 5206
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 15285 4858 15351 4861
rect 22320 4858 22800 4888
rect 15285 4856 22800 4858
rect 15285 4800 15290 4856
rect 15346 4800 22800 4856
rect 15285 4798 22800 4800
rect 15285 4795 15351 4798
rect 22320 4768 22800 4798
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 18597 4314 18663 4317
rect 22320 4314 22800 4344
rect 18597 4312 22800 4314
rect 18597 4256 18602 4312
rect 18658 4256 22800 4312
rect 18597 4254 22800 4256
rect 18597 4251 18663 4254
rect 22320 4224 22800 4254
rect 20253 3906 20319 3909
rect 22320 3906 22800 3936
rect 20253 3904 22800 3906
rect 20253 3848 20258 3904
rect 20314 3848 22800 3904
rect 20253 3846 22800 3848
rect 20253 3843 20319 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 6361 3498 6427 3501
rect 17401 3498 17467 3501
rect 6361 3496 17467 3498
rect 6361 3440 6366 3496
rect 6422 3440 17406 3496
rect 17462 3440 17467 3496
rect 6361 3438 17467 3440
rect 6361 3435 6427 3438
rect 17401 3435 17467 3438
rect 18965 3498 19031 3501
rect 22320 3498 22800 3528
rect 18965 3496 22800 3498
rect 18965 3440 18970 3496
rect 19026 3440 22800 3496
rect 18965 3438 22800 3440
rect 18965 3435 19031 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 10225 3090 10291 3093
rect 12985 3090 13051 3093
rect 10225 3088 13051 3090
rect 10225 3032 10230 3088
rect 10286 3032 12990 3088
rect 13046 3032 13051 3088
rect 10225 3030 13051 3032
rect 10225 3027 10291 3030
rect 12985 3027 13051 3030
rect 18689 2954 18755 2957
rect 22320 2954 22800 2984
rect 18689 2952 22800 2954
rect 18689 2896 18694 2952
rect 18750 2896 22800 2952
rect 18689 2894 22800 2896
rect 18689 2891 18755 2894
rect 22320 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 17902 2620 17908 2684
rect 17972 2682 17978 2684
rect 18413 2682 18479 2685
rect 17972 2680 18479 2682
rect 17972 2624 18418 2680
rect 18474 2624 18479 2680
rect 17972 2622 18479 2624
rect 17972 2620 17978 2622
rect 18413 2619 18479 2622
rect 15653 2546 15719 2549
rect 22320 2546 22800 2576
rect 15653 2544 22800 2546
rect 15653 2488 15658 2544
rect 15714 2488 22800 2544
rect 15653 2486 22800 2488
rect 15653 2483 15719 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 18597 2002 18663 2005
rect 22320 2002 22800 2032
rect 18597 2000 22800 2002
rect 18597 1944 18602 2000
rect 18658 1944 22800 2000
rect 18597 1942 22800 1944
rect 18597 1939 18663 1942
rect 22320 1912 22800 1942
rect 10869 1594 10935 1597
rect 12157 1594 12223 1597
rect 22320 1594 22800 1624
rect 10869 1592 22800 1594
rect 10869 1536 10874 1592
rect 10930 1536 12162 1592
rect 12218 1536 22800 1592
rect 10869 1534 22800 1536
rect 10869 1531 10935 1534
rect 12157 1531 12223 1534
rect 22320 1504 22800 1534
rect 16430 988 16436 1052
rect 16500 1050 16506 1052
rect 22320 1050 22800 1080
rect 16500 990 22800 1050
rect 16500 988 16506 990
rect 22320 960 22800 990
rect 13721 642 13787 645
rect 22320 642 22800 672
rect 13721 640 22800 642
rect 13721 584 13726 640
rect 13782 584 22800 640
rect 13721 582 22800 584
rect 13721 579 13787 582
rect 22320 552 22800 582
rect 18822 172 18828 236
rect 18892 234 18898 236
rect 22320 234 22800 264
rect 18892 174 22800 234
rect 18892 172 18898 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 10732 19076 10796 19140
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 14412 18260 14476 18324
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 16436 16688 16500 16692
rect 16436 16632 16486 16688
rect 16486 16632 16500 16688
rect 16436 16628 16500 16632
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 16804 15192 16868 15196
rect 16804 15136 16854 15192
rect 16854 15136 16868 15192
rect 16804 15132 16868 15136
rect 16988 14996 17052 15060
rect 10732 14860 10796 14924
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 18828 13364 18892 13428
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 17356 12608 17420 12612
rect 17356 12552 17406 12608
rect 17406 12552 17420 12608
rect 17356 12548 17420 12552
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 16436 11460 16500 11524
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 14412 10100 14476 10164
rect 16436 9964 16500 10028
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 17356 7712 17420 7716
rect 17356 7656 17370 7712
rect 17370 7656 17420 7712
rect 17356 7652 17420 7656
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 16804 7380 16868 7444
rect 17908 7244 17972 7308
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 16988 5672 17052 5676
rect 16988 5616 17002 5672
rect 17002 5616 17052 5672
rect 16988 5612 17052 5616
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 17908 2620 17972 2684
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 16436 988 16500 1052
rect 18828 172 18892 236
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 10731 19140 10797 19141
rect 10731 19076 10732 19140
rect 10796 19076 10797 19140
rect 10731 19075 10797 19076
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 10734 14925 10794 19075
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14411 18324 14477 18325
rect 14411 18260 14412 18324
rect 14476 18260 14477 18324
rect 14411 18259 14477 18260
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 10731 14924 10797 14925
rect 10731 14860 10732 14924
rect 10796 14860 10797 14924
rect 10731 14859 10797 14860
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 14414 10165 14474 18259
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 16435 16692 16501 16693
rect 16435 16628 16436 16692
rect 16500 16628 16501 16692
rect 16435 16627 16501 16628
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 16438 11525 16498 16627
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 16803 15196 16869 15197
rect 16803 15132 16804 15196
rect 16868 15132 16869 15196
rect 16803 15131 16869 15132
rect 16435 11524 16501 11525
rect 16435 11460 16436 11524
rect 16500 11460 16501 11524
rect 16435 11459 16501 11460
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14411 10164 14477 10165
rect 14411 10100 14412 10164
rect 14476 10100 14477 10164
rect 14411 10099 14477 10100
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 9280 14992 10304
rect 16435 10028 16501 10029
rect 16435 9964 16436 10028
rect 16500 9964 16501 10028
rect 16435 9963 16501 9964
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 16438 1053 16498 9963
rect 16806 7445 16866 15131
rect 16987 15060 17053 15061
rect 16987 14996 16988 15060
rect 17052 14996 17053 15060
rect 16987 14995 17053 14996
rect 16803 7444 16869 7445
rect 16803 7380 16804 7444
rect 16868 7380 16869 7444
rect 16803 7379 16869 7380
rect 16990 5677 17050 14995
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18827 13428 18893 13429
rect 18827 13364 18828 13428
rect 18892 13364 18893 13428
rect 18827 13363 18893 13364
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 17355 12612 17421 12613
rect 17355 12548 17356 12612
rect 17420 12548 17421 12612
rect 17355 12547 17421 12548
rect 17358 7717 17418 12547
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 17355 7716 17421 7717
rect 17355 7652 17356 7716
rect 17420 7652 17421 7716
rect 17355 7651 17421 7652
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 17907 7308 17973 7309
rect 17907 7244 17908 7308
rect 17972 7244 17973 7308
rect 17907 7243 17973 7244
rect 16987 5676 17053 5677
rect 16987 5612 16988 5676
rect 17052 5612 17053 5676
rect 16987 5611 17053 5612
rect 17910 2685 17970 7243
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 17907 2684 17973 2685
rect 17907 2620 17908 2684
rect 17972 2620 17973 2684
rect 17907 2619 17973 2620
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 16435 1052 16501 1053
rect 16435 988 16436 1052
rect 16500 988 16501 1052
rect 16435 987 16501 988
rect 18830 237 18890 13363
rect 18827 236 18893 237
rect 18827 172 18828 236
rect 18892 172 18893 236
rect 18827 171 18893 172
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606256979
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606256979
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606256979
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606256979
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_98
timestamp 1606256979
transform 1 0 10120 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1606256979
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11224 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106
timestamp 1606256979
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115
timestamp 1606256979
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11592 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606256979
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606256979
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1606256979
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606256979
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14352 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12788 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13524 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13340 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp 1606256979
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1606256979
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1606256979
transform 1 0 12972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1606256979
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606256979
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1606256979
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606256979
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1606256979
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_160
timestamp 1606256979
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15548 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1606256979
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_176
timestamp 1606256979
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1606256979
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16468 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606256979
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606256979
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606256979
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606256979
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606256979
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_192
timestamp 1606256979
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606256979
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1606256979
transform 1 0 19044 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606256979
transform 1 0 18952 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_198
timestamp 1606256979
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606256979
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606256979
transform 1 0 19412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1606256979
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1606256979
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606256979
transform 1 0 19964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_208
timestamp 1606256979
transform 1 0 20240 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1606256979
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1606256979
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606256979
transform 1 0 20332 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606256979
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606256979
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1606256979
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606256979
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606256979
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10028 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11684 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1606256979
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13340 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_131
timestamp 1606256979
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15548 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606256979
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17204 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1606256979
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19044 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19780 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1606256979
transform 1 0 18676 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1606256979
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1606256979
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1606256979
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606256979
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606256979
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606256979
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606256979
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9108 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_86
timestamp 1606256979
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_103
timestamp 1606256979
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606256979
transform 1 0 11776 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1606256979
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606256979
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12788 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1606256979
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606256979
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15732 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1606256979
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1606256979
transform 1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1606256979
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606256979
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606256979
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_171
timestamp 1606256979
transform 1 0 16836 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606256979
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1606256979
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606256979
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1606256979
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1606256979
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606256979
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606256979
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606256979
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606256979
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12236 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606256979
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1606256979
transform 1 0 11868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606256979
transform 1 0 13892 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1606256979
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_143
timestamp 1606256979
transform 1 0 14260 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606256979
transform 1 0 16284 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606256979
transform 1 0 14536 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1606256979
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1606256979
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606256979
transform 1 0 17296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1606256979
transform 1 0 17756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_168
timestamp 1606256979
transform 1 0 16560 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_179
timestamp 1606256979
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 19780 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18768 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1606256979
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1606256979
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606256979
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606256979
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606256979
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606256979
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606256979
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606256979
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_98
timestamp 1606256979
transform 1 0 10120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11408 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1606256979
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1606256979
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1606256979
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13708 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_133
timestamp 1606256979
transform 1 0 13340 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606256979
transform 1 0 15364 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15916 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_153
timestamp 1606256979
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_159
timestamp 1606256979
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_177
timestamp 1606256979
transform 1 0 17388 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18492 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 20148 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_188
timestamp 1606256979
transform 1 0 18400 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_205
timestamp 1606256979
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1606256979
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606256979
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606256979
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606256979
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606256979
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606256979
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606256979
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606256979
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8464 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606256979
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606256979
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1606256979
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1606256979
transform 1 0 10580 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1606256979
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10948 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12604 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_123
timestamp 1606256979
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1606256979
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606256979
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606256979
transform 1 0 13616 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13432 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1606256979
transform 1 0 14444 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_134
timestamp 1606256979
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_139
timestamp 1606256979
transform 1 0 13892 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1606256979
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_143
timestamp 1606256979
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15640 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606256979
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1606256979
transform 1 0 15272 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_167
timestamp 1606256979
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_174
timestamp 1606256979
transform 1 0 17112 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1606256979
transform 1 0 16744 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16652 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1606256979
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1606256979
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18216 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17204 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18860 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 19228 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1606256979
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1606256979
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1606256979
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1606256979
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_218
timestamp 1606256979
transform 1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_213
timestamp 1606256979
transform 1 0 20700 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1606256979
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606256979
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606256979
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606256979
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606256979
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_80
timestamp 1606256979
transform 1 0 8464 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606256979
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 10672 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_86
timestamp 1606256979
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606256979
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1606256979
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11684 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_113
timestamp 1606256979
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13800 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_131
timestamp 1606256979
transform 1 0 13156 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_137
timestamp 1606256979
transform 1 0 13708 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 16284 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_147
timestamp 1606256979
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606256979
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17848 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp 1606256979
transform 1 0 16560 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1606256979
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1606256979
transform 1 0 18676 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1606256979
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1606256979
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606256979
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606256979
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1606256979
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1606256979
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1606256979
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606256979
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1606256979
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_78
timestamp 1606256979
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1606256979
transform 1 0 9844 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1606256979
transform 1 0 10212 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1606256979
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606256979
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13800 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12788 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1606256979
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1606256979
transform 1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15456 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_147
timestamp 1606256979
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1606256979
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606256979
transform 1 0 17112 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1606256979
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1606256979
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_193
timestamp 1606256979
transform 1 0 18860 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_201
timestamp 1606256979
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_213
timestamp 1606256979
transform 1 0 20700 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606256979
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606256979
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606256979
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606256979
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1606256979
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1606256979
transform 1 0 8464 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9844 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606256979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1606256979
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10856 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12512 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1606256979
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1606256979
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15640 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606256979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16652 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_167
timestamp 1606256979
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1606256979
transform 1 0 18124 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18860 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1606256979
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1606256979
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1606256979
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606256979
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606256979
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606256979
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1606256979
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8188 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_74
timestamp 1606256979
transform 1 0 7912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9200 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1606256979
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_104
timestamp 1606256979
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606256979
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10856 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1606256979
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606256979
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13800 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_147
timestamp 1606256979
transform 1 0 14628 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp 1606256979
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 16744 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1606256979
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1606256979
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18584 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_199
timestamp 1606256979
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_210
timestamp 1606256979
transform 1 0 20424 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_218
timestamp 1606256979
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606256979
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606256979
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606256979
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606256979
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606256979
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1606256979
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9752 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606256979
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11408 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 12420 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1606256979
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1606256979
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12972 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_126
timestamp 1606256979
transform 1 0 12696 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1606256979
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15732 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1606256979
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17664 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 17388 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1606256979
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18676 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1606256979
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1606256979
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606256979
transform 1 0 20332 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1606256979
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606256979
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606256979
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1606256979
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1606256979
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606256979
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1606256979
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1606256979
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8188 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_13_74
timestamp 1606256979
transform 1 0 7912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_68
timestamp 1606256979
transform 1 0 7360 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9936 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_93
timestamp 1606256979
transform 1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_96
timestamp 1606256979
transform 1 0 9936 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11592 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1606256979
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606256979
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_119
timestamp 1606256979
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13156 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1606256979
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1606256979
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1606256979
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14536 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15548 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1606256979
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_166
timestamp 1606256979
transform 1 0 16376 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606256979
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16928 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18124 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606256979
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1606256979
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1606256979
transform 1 0 17756 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 19136 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1606256979
transform 1 0 20056 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_200
timestamp 1606256979
transform 1 0 19504 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1606256979
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606256979
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606256979
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1606256979
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606256979
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1606256979
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1606256979
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1606256979
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8740 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_74
timestamp 1606256979
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_82
timestamp 1606256979
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9752 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1606256979
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_100
timestamp 1606256979
transform 1 0 10304 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_108
timestamp 1606256979
transform 1 0 11040 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_143
timestamp 1606256979
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14536 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_164
timestamp 1606256979
transform 1 0 16192 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606256979
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp 1606256979
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19596 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1606256979
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_217
timestamp 1606256979
transform 1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606256979
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606256979
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1606256979
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1606256979
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_16_68
timestamp 1606256979
transform 1 0 7360 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606256979
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1606256979
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10856 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_16_122
timestamp 1606256979
transform 1 0 12328 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12972 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_16_128
timestamp 1606256979
transform 1 0 12880 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16100 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606256979
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16652 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18308 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1606256979
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19596 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_196
timestamp 1606256979
transform 1 0 19136 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_200
timestamp 1606256979
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1606256979
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606256979
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606256979
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606256979
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606256979
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606256979
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1606256979
transform 1 0 7912 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_82
timestamp 1606256979
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606256979
transform 1 0 10580 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606256979
transform 1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9384 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1606256979
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_96
timestamp 1606256979
transform 1 0 9936 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_102
timestamp 1606256979
transform 1 0 10488 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606256979
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_106
timestamp 1606256979
transform 1 0 10856 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13432 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 14260 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_133
timestamp 1606256979
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15456 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1606256979
transform 1 0 15088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_165
timestamp 1606256979
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16836 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 16468 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_170
timestamp 1606256979
transform 1 0 16744 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1606256979
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606256979
transform 1 0 19136 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 19688 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_193
timestamp 1606256979
transform 1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1606256979
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1606256979
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606256979
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606256979
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1606256979
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1606256979
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7728 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1606256979
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10304 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1606256979
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1606256979
transform 1 0 10212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 11408 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_109
timestamp 1606256979
transform 1 0 11132 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13064 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1606256979
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15916 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_146
timestamp 1606256979
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1606256979
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1606256979
transform 1 0 15548 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1606256979
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1606256979
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606256979
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18584 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1606256979
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1606256979
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606256979
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606256979
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606256979
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606256979
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606256979
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606256979
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606256979
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606256979
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606256979
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1606256979
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1606256979
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_74
timestamp 1606256979
transform 1 0 7912 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_82
timestamp 1606256979
transform 1 0 8648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1606256979
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_80
timestamp 1606256979
transform 1 0 8464 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8924 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1606256979
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_88
timestamp 1606256979
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11316 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11592 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1606256979
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606256979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1606256979
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_120
timestamp 1606256979
transform 1 0 12144 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606256979
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13064 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 12696 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_132
timestamp 1606256979
transform 1 0 13248 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_129
timestamp 1606256979
transform 1 0 12972 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1606256979
transform 1 0 13616 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_143
timestamp 1606256979
transform 1 0 14260 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606256979
transform 1 0 16284 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606256979
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15180 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1606256979
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606256979
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606256979
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17756 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 16836 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16744 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1606256979
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1606256979
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1606256979
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1606256979
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606256979
transform 1 0 18768 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18768 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1606256979
transform 1 0 19320 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1606256979
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1606256979
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1606256979
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_196
timestamp 1606256979
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1606256979
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 20424 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_216
timestamp 1606256979
transform 1 0 20976 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1606256979
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1606256979
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1606256979
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606256979
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606256979
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8464 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_74
timestamp 1606256979
transform 1 0 7912 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606256979
transform 1 0 9476 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1606256979
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_94
timestamp 1606256979
transform 1 0 9752 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1606256979
transform 1 0 10948 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1606256979
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1606256979
transform 1 0 13616 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1606256979
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1606256979
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606256979
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16284 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 14628 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_156
timestamp 1606256979
transform 1 0 15456 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1606256979
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606256979
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19044 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1606256979
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1606256979
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_201
timestamp 1606256979
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606256979
transform 1 0 20792 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1606256979
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1606256979
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606256979
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606256979
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1606256979
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8464 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1606256979
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1606256979
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11592 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 11316 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1606256979
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13248 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14260 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1606256979
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1606256979
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16100 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1606256979
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_160
timestamp 1606256979
transform 1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 17756 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_179
timestamp 1606256979
transform 1 0 17572 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 19044 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_190
timestamp 1606256979
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_194
timestamp 1606256979
transform 1 0 18952 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1606256979
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1606256979
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606256979
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1606256979
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_39
timestamp 1606256979
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1606256979
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606256979
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7636 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_70
timestamp 1606256979
transform 1 0 7544 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10304 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9292 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_87
timestamp 1606256979
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1606256979
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1606256979
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606256979
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14260 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13064 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1606256979
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606256979
transform 1 0 16100 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1606256979
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16652 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_167
timestamp 1606256979
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1606256979
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1606256979
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18492 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19596 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_188
timestamp 1606256979
transform 1 0 18400 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_198
timestamp 1606256979
transform 1 0 19320 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606256979
transform 1 0 20608 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1606256979
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_216
timestamp 1606256979
transform 1 0 20976 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1606256979
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606256979
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6164 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_44
timestamp 1606256979
transform 1 0 5152 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_52
timestamp 1606256979
transform 1 0 5888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_71
timestamp 1606256979
transform 1 0 7636 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1606256979
transform 1 0 8740 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10396 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8832 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606256979
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_99
timestamp 1606256979
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 11500 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_110
timestamp 1606256979
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13156 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1606256979
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_140
timestamp 1606256979
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16376 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1606256979
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_163
timestamp 1606256979
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606256979
transform 1 0 18032 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1606256979
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_187
timestamp 1606256979
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606256979
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18492 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_205
timestamp 1606256979
transform 1 0 19964 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606256979
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1606256979
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1606256979
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1606256979
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1606256979
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606256979
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8648 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1606256979
transform 1 0 8280 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9384 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_88
timestamp 1606256979
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1606256979
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1606256979
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606256979
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606256979
transform 1 0 13432 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 13984 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1606256979
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1606256979
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15640 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1606256979
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1606256979
transform 1 0 16652 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_167
timestamp 1606256979
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_178
timestamp 1606256979
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19780 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_200
timestamp 1606256979
transform 1 0 19504 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606256979
transform 1 0 20792 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1606256979
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_218
timestamp 1606256979
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606256979
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1606256979
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1606256979
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1606256979
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1606256979
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606256979
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_56
timestamp 1606256979
transform 1 0 6256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1606256979
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606256979
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6992 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6992 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8188 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8648 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_73
timestamp 1606256979
transform 1 0 7820 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1606256979
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1606256979
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_86
timestamp 1606256979
transform 1 0 9016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1606256979
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_96
timestamp 1606256979
transform 1 0 9936 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10212 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606256979
transform 1 0 11776 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11868 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12604 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1606256979
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_113
timestamp 1606256979
transform 1 0 11500 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1606256979
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13892 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1606256979
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_134
timestamp 1606256979
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_138
timestamp 1606256979
transform 1 0 13800 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_152
timestamp 1606256979
transform 1 0 15088 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1606256979
transform 1 0 14720 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606256979
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606256979
transform 1 0 15180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1606256979
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1606256979
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1606256979
transform 1 0 15732 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15732 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1606256979
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_168
timestamp 1606256979
transform 1 0 16560 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1606256979
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16744 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606256979
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606256979
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1606256979
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_179
timestamp 1606256979
transform 1 0 17572 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17848 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18584 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1606256979
transform 1 0 19596 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19964 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1606256979
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1606256979
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1606256979
transform 1 0 19504 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1606256979
transform 1 0 19872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1606256979
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606256979
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_214
timestamp 1606256979
transform 1 0 20792 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1606256979
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1606256979
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606256979
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606256979
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7452 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_68
timestamp 1606256979
transform 1 0 7360 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1606256979
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1606256979
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_102
timestamp 1606256979
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606256979
transform 1 0 12512 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10764 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11500 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1606256979
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1606256979
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12972 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13984 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1606256979
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1606256979
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606256979
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15732 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1606256979
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606256979
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_157
timestamp 1606256979
transform 1 0 15548 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17112 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_28_168
timestamp 1606256979
transform 1 0 16560 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19780 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18768 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1606256979
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1606256979
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1606256979
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1606256979
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_218
timestamp 1606256979
transform 1 0 21160 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1606256979
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1606256979
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1606256979
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1606256979
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_74
timestamp 1606256979
transform 1 0 7912 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_82
timestamp 1606256979
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10028 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_93
timestamp 1606256979
transform 1 0 9660 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1606256979
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11040 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1606256979
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1606256979
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606256979
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13984 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12972 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_127
timestamp 1606256979
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_138
timestamp 1606256979
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606256979
transform 1 0 15732 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16284 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_156
timestamp 1606256979
transform 1 0 15456 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_163
timestamp 1606256979
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606256979
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606256979
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19688 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_193
timestamp 1606256979
transform 1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1606256979
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_208
timestamp 1606256979
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 20424 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_216
timestamp 1606256979
transform 1 0 20976 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1606256979
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1606256979
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606256979
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1606256979
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7820 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1606256979
transform 1 0 7360 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_72
timestamp 1606256979
transform 1 0 7728 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1606256979
transform 1 0 10028 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10580 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_89
timestamp 1606256979
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_101
timestamp 1606256979
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_119
timestamp 1606256979
transform 1 0 12052 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1606256979
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12696 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_142
timestamp 1606256979
transform 1 0 14168 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1606256979
transform 1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1606256979
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606256979
transform 1 0 17572 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606256979
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18124 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1606256979
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_176
timestamp 1606256979
transform 1 0 17296 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1606256979
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606256979
transform 1 0 19136 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19688 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1606256979
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_200
timestamp 1606256979
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1606256979
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606256979
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1606256979
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1606256979
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1606256979
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606256979
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8556 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_74
timestamp 1606256979
transform 1 0 7912 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1606256979
transform 1 0 8464 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10212 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1606256979
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_115
timestamp 1606256979
transform 1 0 11684 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1606256979
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1606256979
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606256979
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_145
timestamp 1606256979
transform 1 0 14444 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15732 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14720 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1606256979
transform 1 0 15272 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_158
timestamp 1606256979
transform 1 0 15640 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17020 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18216 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_168
timestamp 1606256979
transform 1 0 16560 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_172
timestamp 1606256979
transform 1 0 16928 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1606256979
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606256979
transform 1 0 19044 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 19596 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_192
timestamp 1606256979
transform 1 0 18768 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_199
timestamp 1606256979
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_213
timestamp 1606256979
transform 1 0 20700 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606256979
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606256979
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606256979
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606256979
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606256979
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606256979
transform 1 0 8556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_75
timestamp 1606256979
transform 1 0 8004 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606256979
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10028 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1606256979
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1606256979
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_94
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606256979
transform 1 0 11040 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_106
timestamp 1606256979
transform 1 0 10856 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_111
timestamp 1606256979
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606256979
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1606256979
transform 1 0 13800 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1606256979
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1606256979
transform 1 0 12788 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_131
timestamp 1606256979
transform 1 0 13156 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_137
timestamp 1606256979
transform 1 0 13708 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_142
timestamp 1606256979
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606256979
transform 1 0 15548 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1606256979
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_148
timestamp 1606256979
transform 1 0 14720 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1606256979
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_156
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1606256979
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606256979
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1606256979
transform 1 0 16652 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1606256979
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1606256979
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_179
timestamp 1606256979
transform 1 0 17572 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1606256979
transform 1 0 18124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606256979
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606256979
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1606256979
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1606256979
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1606256979
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606256979
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1606256979
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606256979
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 5720 480 5840 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 17144 480 17264 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 22320 3816 22800 3936 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 846 0 902 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 1950 0 2006 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2502 0 2558 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 846 22320 902 22800 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 6366 22320 6422 22800 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 6918 22320 6974 22800 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 7470 22320 7526 22800 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 8022 22320 8078 22800 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 8574 22320 8630 22800 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 9126 22320 9182 22800 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 9678 22320 9734 22800 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 10230 22320 10286 22800 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 10782 22320 10838 22800 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 11334 22320 11390 22800 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1398 22320 1454 22800 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 1950 22320 2006 22800 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2502 22320 2558 22800 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3054 22320 3110 22800 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 3606 22320 3662 22800 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4158 22320 4214 22800 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 5262 22320 5318 22800 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 5814 22320 5870 22800 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 18050 22320 18106 22800 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 18602 22320 18658 22800 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 19706 22320 19762 22800 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 20258 22320 20314 22800 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 20810 22320 20866 22800 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 21362 22320 21418 22800 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 21914 22320 21970 22800 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 22466 22320 22522 22800 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 12530 22320 12586 22800 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 13082 22320 13138 22800 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 13634 22320 13690 22800 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 14186 22320 14242 22800 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 14738 22320 14794 22800 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 15290 22320 15346 22800 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 15842 22320 15898 22800 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 16394 22320 16450 22800 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 16946 22320 17002 22800 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 22320 22448 22800 22568 6 prog_clk_0_E_in
port 123 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 124 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 125 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 126 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 127 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 128 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 129 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 130 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 131 nsew default input
rlabel metal2 s 294 22320 350 22800 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 133 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
