* NGSPICE file created from cby_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

.subckt cby_0__1_ ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] left_grid_pin_0_ prog_clk right_grid_pin_52_
+ vpwr vgnd
XFILLER_22_133 vgnd vpwr scs8hd_decap_12
XFILLER_3_78 vgnd vpwr scs8hd_decap_12
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_1__A1 mux_left_ipin_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_0__S mux_left_ipin_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_23_86 vgnd vpwr scs8hd_decap_12
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l3_in_0__A1 mux_left_ipin_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_56_117 vgnd vpwr scs8hd_decap_12
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XFILLER_34_85 vgnd vpwr scs8hd_decap_6
XFILLER_18_86 vgnd vpwr scs8hd_decap_3
XFILLER_55_29 vgnd vpwr scs8hd_decap_4
XFILLER_29_41 vgnd vpwr scs8hd_decap_8
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_40_145 vgnd vpwr scs8hd_fill_1
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XFILLER_31_112 vgnd vpwr scs8hd_decap_8
XFILLER_31_75 vgnd vpwr scs8hd_decap_12
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l2_in_3__S mux_left_ipin_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_22_145 vgnd vpwr scs8hd_fill_1
XFILLER_42_30 vgnd vpwr scs8hd_fill_1
XFILLER_13_101 vgnd vpwr scs8hd_decap_12
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_53_95 vpwr vgnd scs8hd_fill_2
XFILLER_45_6 vpwr vgnd scs8hd_fill_2
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_23_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_36 vpwr vgnd scs8hd_fill_2
XFILLER_56_129 vgnd vpwr scs8hd_decap_12
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_61_143 vgnd vpwr scs8hd_decap_3
XFILLER_61_110 vgnd vpwr scs8hd_decap_12
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_52_143 vgnd vpwr scs8hd_decap_3
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
XFILLER_43_143 vgnd vpwr scs8hd_decap_3
XFILLER_43_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_25_143 vgnd vpwr scs8hd_decap_3
XFILLER_25_110 vgnd vpwr scs8hd_decap_12
XFILLER_31_135 vgnd vpwr scs8hd_decap_8
XFILLER_31_87 vgnd vpwr scs8hd_decap_6
XFILLER_31_54 vgnd vpwr scs8hd_fill_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0__S mux_right_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_113 vgnd vpwr scs8hd_decap_8
XFILLER_13_135 vgnd vpwr scs8hd_decap_8
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_4_90 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vgnd vpwr scs8hd_fill_1
XFILLER_0_48 vpwr vgnd scs8hd_fill_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_47_108 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_4
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_59_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_46_141 vgnd vpwr scs8hd_decap_4
XFILLER_52_111 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A0 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_61_74 vgnd vpwr scs8hd_decap_12
XFILLER_45_75 vgnd vpwr scs8hd_decap_12
XFILLER_45_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_54 vpwr vgnd scs8hd_fill_2
XFILLER_28_141 vgnd vpwr scs8hd_decap_4
XANTENNA__04__A chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A0 mux_right_ipin_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_42_21 vgnd vpwr scs8hd_fill_1
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_53_75 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.mux_l3_in_1__S mux_left_ipin_0.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA__12__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_131 vgnd vpwr scs8hd_decap_12
XANTENNA__07__A chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XFILLER_59_74 vgnd vpwr scs8hd_decap_12
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
XFILLER_52_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A1 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
X_29_ chany_top_in[11] chany_bottom_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_61_86 vgnd vpwr scs8hd_decap_12
XFILLER_45_87 vgnd vpwr scs8hd_decap_12
XFILLER_45_10 vgnd vpwr scs8hd_decap_12
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_66 vgnd vpwr scs8hd_decap_12
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_145 vgnd vpwr scs8hd_fill_1
XANTENNA__20__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_31_23 vpwr vgnd scs8hd_fill_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_79 vgnd vpwr scs8hd_decap_12
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A1 mux_right_ipin_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_145 vgnd vpwr scs8hd_fill_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XANTENNA__15__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_53_87 vgnd vpwr scs8hd_decap_4
XFILLER_53_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_111 vgnd vpwr scs8hd_decap_8
XFILLER_48_32 vgnd vpwr scs8hd_decap_12
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_55_143 vgnd vpwr scs8hd_decap_3
XFILLER_55_121 vgnd vpwr scs8hd_fill_1
XFILLER_18_68 vgnd vpwr scs8hd_decap_4
XFILLER_61_135 vgnd vpwr scs8hd_decap_8
XFILLER_59_86 vgnd vpwr scs8hd_decap_12
XFILLER_50_44 vgnd vpwr scs8hd_decap_12
XANTENNA__23__A chany_top_in[17] vgnd vpwr scs8hd_diode_2
X_28_ chany_top_in[12] chany_bottom_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_52_135 vgnd vpwr scs8hd_decap_8
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_143 vgnd vpwr scs8hd_decap_3
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XFILLER_61_98 vgnd vpwr scs8hd_decap_12
XANTENNA__18__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_45_99 vgnd vpwr scs8hd_decap_12
XFILLER_45_22 vgnd vpwr scs8hd_decap_12
XFILLER_43_135 vgnd vpwr scs8hd_decap_8
XFILLER_29_78 vgnd vpwr scs8hd_decap_12
XFILLER_19_143 vgnd vpwr scs8hd_decap_3
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_8
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__31__A chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_1__S mux_right_ipin_0.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_53_99 vpwr vgnd scs8hd_fill_2
XFILLER_53_66 vpwr vgnd scs8hd_fill_2
XFILLER_53_33 vpwr vgnd scs8hd_fill_2
XANTENNA__26__A chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_58_141 vgnd vpwr scs8hd_decap_4
XFILLER_48_99 vgnd vpwr scs8hd_fill_1
XFILLER_48_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_59_98 vgnd vpwr scs8hd_decap_12
XFILLER_50_56 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_27_ chany_top_in[13] chany_bottom_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_45_34 vgnd vpwr scs8hd_decap_12
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__D mux_left_ipin_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A0 _03_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__34__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_decap_3
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__29__A chany_top_in[11] vgnd vpwr scs8hd_diode_2
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_42_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_24 vgnd vpwr scs8hd_decap_6
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_121 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XANTENNA__42__A chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_53_45 vpwr vgnd scs8hd_fill_2
XFILLER_5_135 vgnd vpwr scs8hd_decap_8
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_48_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA__37__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_64_145 vgnd vpwr scs8hd_fill_1
X_43_ chany_bottom_in[17] chany_top_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_55_101 vpwr vgnd scs8hd_fill_2
XFILLER_50_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_46_145 vgnd vpwr scs8hd_fill_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
X_26_ chany_top_in[14] chany_bottom_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_0.scs8hd_buf_4_0__A mux_left_ipin_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_58 vgnd vpwr scs8hd_decap_3
XFILLER_28_145 vgnd vpwr scs8hd_fill_1
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_62 vgnd vpwr scs8hd_decap_4
XFILLER_1_51 vgnd vpwr scs8hd_decap_4
XFILLER_45_57 vpwr vgnd scs8hd_fill_2
XFILLER_45_46 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
X_09_ chany_bottom_in[11] chany_top_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XPHY_121 vgnd vpwr scs8hd_decap_3
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_15 vgnd vpwr scs8hd_decap_8
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_92 vgnd vpwr scs8hd_fill_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_50 vgnd vpwr scs8hd_decap_8
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_133 vgnd vpwr scs8hd_decap_12
XFILLER_53_57 vgnd vpwr scs8hd_fill_1
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
XFILLER_48_68 vgnd vpwr scs8hd_decap_12
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
X_42_ chany_bottom_in[18] chany_top_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_49_143 vgnd vpwr scs8hd_decap_3
XFILLER_13_60 vgnd vpwr scs8hd_fill_1
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_25_ chany_top_in[15] chany_bottom_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_8
XFILLER_29_15 vgnd vpwr scs8hd_decap_4
XFILLER_19_102 vpwr vgnd scs8hd_fill_2
X_08_ chany_bottom_in[12] chany_top_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_135 vgnd vpwr scs8hd_decap_8
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_decap_3
XFILLER_31_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_15 vgnd vpwr scs8hd_decap_6
XFILLER_30_141 vgnd vpwr scs8hd_decap_4
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_145 vgnd vpwr scs8hd_fill_1
XFILLER_12_141 vgnd vpwr scs8hd_decap_4
XFILLER_53_25 vpwr vgnd scs8hd_fill_2
XFILLER_53_14 vgnd vpwr scs8hd_fill_1
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
X_41_ chany_bottom_in[19] chany_top_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_49_111 vgnd vpwr scs8hd_decap_8
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XFILLER_34_38 vgnd vpwr scs8hd_decap_12
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_75 vgnd vpwr scs8hd_decap_12
X_24_ chany_top_in[16] chany_bottom_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_29_49 vgnd vpwr scs8hd_decap_3
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
X_07_ chany_bottom_in[13] chany_top_out[13] vgnd vpwr scs8hd_buf_2
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_46_80 vgnd vpwr scs8hd_decap_12
XFILLER_22_109 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_32_93 vgnd vpwr scs8hd_fill_1
XFILLER_53_37 vpwr vgnd scs8hd_fill_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_97 vgnd vpwr scs8hd_fill_1
XFILLER_58_145 vgnd vpwr scs8hd_fill_1
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
X_40_ chany_top_in[0] chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_13_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_0__S mux_left_ipin_0.mux_l1_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_13_73 vpwr vgnd scs8hd_fill_2
XFILLER_64_137 vgnd vpwr scs8hd_decap_8
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_23_ chany_top_in[17] chany_bottom_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_1_87 vgnd vpwr scs8hd_decap_12
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_51_92 vgnd vpwr scs8hd_fill_1
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XFILLER_19_94 vpwr vgnd scs8hd_fill_2
X_06_ chany_bottom_in[14] chany_top_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_31 vgnd vpwr scs8hd_fill_1
XFILLER_7_86 vgnd vpwr scs8hd_decap_3
XFILLER_21_143 vgnd vpwr scs8hd_decap_3
XFILLER_53_49 vgnd vpwr scs8hd_decap_8
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_0__A0 mux_left_ipin_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_76 vgnd vpwr scs8hd_decap_12
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l4_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_13_52 vpwr vgnd scs8hd_fill_2
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XFILLER_54_70 vgnd vpwr scs8hd_decap_3
XFILLER_49_135 vgnd vpwr scs8hd_decap_8
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__D mux_right_ipin_0.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_59_59 vpwr vgnd scs8hd_fill_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_127 vpwr vgnd scs8hd_fill_2
XFILLER_55_105 vgnd vpwr scs8hd_decap_12
XFILLER_46_105 vgnd vpwr scs8hd_decap_12
X_22_ chany_top_in[18] chany_bottom_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_1_99 vgnd vpwr scs8hd_decap_12
XFILLER_1_66 vgnd vpwr scs8hd_fill_1
XFILLER_1_55 vgnd vpwr scs8hd_fill_1
XFILLER_60_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.scs8hd_buf_4_0__A mux_right_ipin_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
X_05_ chany_bottom_in[15] chany_top_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XPHY_103 vgnd vpwr scs8hd_decap_3
XFILLER_24_141 vgnd vpwr scs8hd_decap_4
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_46_93 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_16_74 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.scs8hd_buf_4_0_ mux_left_ipin_0.mux_l4_in_0_/X right_grid_pin_52_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_ipin_0.mux_l2_in_0__A1 mux_left_ipin_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_107 vpwr vgnd scs8hd_fill_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_1_143 vgnd vpwr scs8hd_decap_3
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XFILLER_55_117 vgnd vpwr scs8hd_decap_4
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_21_ chany_top_in[19] chany_bottom_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_46_117 vgnd vpwr scs8hd_decap_12
XFILLER_1_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_19 vgnd vpwr scs8hd_fill_1
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_19_106 vgnd vpwr scs8hd_decap_12
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
X_04_ chany_bottom_in[16] chany_top_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_145 vgnd vpwr scs8hd_fill_1
XFILLER_21_86 vgnd vpwr scs8hd_decap_6
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
XFILLER_16_86 vgnd vpwr scs8hd_decap_3
XFILLER_12_145 vgnd vpwr scs8hd_fill_1
XFILLER_5_119 vgnd vpwr scs8hd_decap_3
XFILLER_43_62 vgnd vpwr scs8hd_decap_12
XFILLER_43_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_fill_1
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XFILLER_54_50 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.mux_l2_in_1__S mux_left_ipin_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_1_111 vgnd vpwr scs8hd_decap_8
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_59_39 vgnd vpwr scs8hd_decap_12
XFILLER_46_129 vgnd vpwr scs8hd_decap_12
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
X_20_ chany_bottom_in[0] chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_1_35 vpwr vgnd scs8hd_fill_2
XFILLER_51_143 vgnd vpwr scs8hd_decap_3
XFILLER_51_121 vgnd vpwr scs8hd_fill_1
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XFILLER_19_118 vgnd vpwr scs8hd_decap_4
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_51_62 vgnd vpwr scs8hd_decap_12
X_03_ _03_/HI _03_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_19_86 vgnd vpwr scs8hd_decap_8
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XFILLER_33_143 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_121 vgnd vpwr scs8hd_fill_1
XFILLER_15_143 vgnd vpwr scs8hd_decap_3
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.mux_l2_in_3__A0 _02_/HI vgnd vpwr scs8hd_diode_2
XFILLER_7_34 vpwr vgnd scs8hd_fill_2
XFILLER_32_75 vpwr vgnd scs8hd_fill_2
XFILLER_32_64 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_43_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
XFILLER_4_131 vgnd vpwr scs8hd_decap_12
XFILLER_58_105 vgnd vpwr scs8hd_decap_12
XFILLER_54_62 vgnd vpwr scs8hd_decap_8
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XFILLER_13_66 vgnd vpwr scs8hd_fill_1
XFILLER_13_77 vgnd vpwr scs8hd_decap_12
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_53_3 vgnd vpwr scs8hd_decap_3
XFILLER_49_62 vgnd vpwr scs8hd_decap_12
XFILLER_49_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_58 vgnd vpwr scs8hd_decap_3
XFILLER_1_47 vpwr vgnd scs8hd_fill_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_51_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_122 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_19_98 vpwr vgnd scs8hd_fill_2
XFILLER_18_141 vgnd vpwr scs8hd_decap_4
X_02_ _02_/HI _02_/LO vgnd vpwr scs8hd_conb_1
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_114 vgnd vpwr scs8hd_decap_8
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_3__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_43_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1__S mux_right_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_143 vgnd vpwr scs8hd_decap_3
XFILLER_58_117 vgnd vpwr scs8hd_decap_12
XFILLER_49_106 vgnd vpwr scs8hd_decap_3
XFILLER_1_135 vgnd vpwr scs8hd_decap_8
XFILLER_13_56 vpwr vgnd scs8hd_fill_2
XFILLER_13_89 vgnd vpwr scs8hd_decap_12
XFILLER_54_30 vgnd vpwr scs8hd_fill_1
XFILLER_60_145 vgnd vpwr scs8hd_fill_1
XFILLER_49_74 vgnd vpwr scs8hd_decap_12
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_40_21 vgnd vpwr scs8hd_fill_1
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_15 vgnd vpwr scs8hd_decap_4
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_51_86 vgnd vpwr scs8hd_decap_6
XFILLER_51_31 vgnd vpwr scs8hd_fill_1
XFILLER_42_134 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XANTENNA__10__A chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vgnd vpwr scs8hd_fill_1
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_7_58 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XFILLER_57_74 vgnd vpwr scs8hd_decap_12
XANTENNA__05__A chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_3
XFILLER_16_56 vgnd vpwr scs8hd_decap_3
XFILLER_43_98 vgnd vpwr scs8hd_decap_12
XFILLER_43_43 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_0.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_0.mux_l3_in_1_/S ccff_tail
+ mem_right_ipin_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_58_129 vgnd vpwr scs8hd_decap_12
XFILLER_54_97 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_63_143 vgnd vpwr scs8hd_decap_3
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XFILLER_54_121 vgnd vpwr scs8hd_fill_1
XFILLER_48_140 vgnd vpwr scs8hd_decap_6
XANTENNA__13__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_49_86 vgnd vpwr scs8hd_decap_12
XFILLER_45_143 vgnd vpwr scs8hd_decap_3
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_135 vgnd vpwr scs8hd_decap_8
XFILLER_51_113 vpwr vgnd scs8hd_fill_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XANTENNA__08__A chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_35_33 vgnd vpwr scs8hd_fill_1
XFILLER_27_143 vgnd vpwr scs8hd_decap_3
XFILLER_27_110 vgnd vpwr scs8hd_decap_12
XFILLER_33_135 vgnd vpwr scs8hd_decap_8
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_46_32 vgnd vpwr scs8hd_decap_12
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_135 vgnd vpwr scs8hd_decap_8
XFILLER_57_86 vgnd vpwr scs8hd_decap_12
XANTENNA__21__A chany_top_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_4
XFILLER_8_109 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA__16__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_0.mux_l2_in_3_/S mux_right_ipin_0.mux_l3_in_1_/S
+ mem_right_ipin_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_0.mux_l2_in_3_ _03_/HI chany_top_in[17] mux_right_ipin_0.mux_l2_in_3_/S
+ mux_right_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_47 vgnd vpwr scs8hd_decap_3
XFILLER_13_69 vpwr vgnd scs8hd_fill_2
XFILLER_54_10 vgnd vpwr scs8hd_decap_8
XFILLER_49_119 vgnd vpwr scs8hd_decap_3
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_49_98 vgnd vpwr scs8hd_decap_8
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XFILLER_45_111 vgnd vpwr scs8hd_decap_8
XFILLER_1_39 vpwr vgnd scs8hd_fill_2
XFILLER_51_103 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ ccff_tail mux_right_ipin_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_45 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_51_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A0 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA__24__A chany_top_in[16] vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XFILLER_2_60 vgnd vpwr scs8hd_decap_12
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XANTENNA__19__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_46_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_7_27 vgnd vpwr scs8hd_decap_4
XFILLER_7_38 vgnd vpwr scs8hd_decap_12
XFILLER_15_103 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A0 mux_right_ipin_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_79 vgnd vpwr scs8hd_decap_12
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_57_98 vgnd vpwr scs8hd_decap_12
XFILLER_7_143 vgnd vpwr scs8hd_decap_3
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_0.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_0.mux_l1_in_2_/S mux_right_ipin_0.mux_l2_in_3_/S
+ mem_right_ipin_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XANTENNA__32__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_2__S mux_right_ipin_0.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[11] mux_right_ipin_0.mux_l2_in_3_/S
+ mux_right_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A0 mux_right_ipin_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_77 vgnd vpwr scs8hd_decap_12
XFILLER_54_44 vpwr vgnd scs8hd_fill_2
XFILLER_54_22 vgnd vpwr scs8hd_decap_8
XANTENNA__27__A chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_40_24 vgnd vpwr scs8hd_decap_6
XFILLER_45_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_145 vgnd vpwr scs8hd_fill_1
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_51_34 vgnd vpwr scs8hd_decap_12
XFILLER_35_57 vgnd vpwr scs8hd_decap_4
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l4_in_0__S mux_left_ipin_0.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_18_145 vgnd vpwr scs8hd_fill_1
XANTENNA__40__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A1 chany_top_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_72 vgnd vpwr scs8hd_decap_12
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XFILLER_46_56 vgnd vpwr scs8hd_decap_3
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__D mux_left_ipin_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XANTENNA__35__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_15_115 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A1 mux_right_ipin_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_58 vgnd vpwr scs8hd_decap_4
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_80 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_0.scs8hd_dfxbp_1_0_ prog_clk mux_left_ipin_0.mux_l4_in_0_/S mux_right_ipin_0.mux_l1_in_2_/S
+ mem_right_ipin_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_93 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l2_in_1_ chany_bottom_in[11] mux_right_ipin_0.mux_l1_in_2_/X
+ mux_right_ipin_0.mux_l2_in_3_/S mux_right_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A1 mux_right_ipin_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_143 vgnd vpwr scs8hd_decap_3
XFILLER_57_110 vgnd vpwr scs8hd_decap_12
XFILLER_54_89 vgnd vpwr scs8hd_decap_3
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_63_135 vgnd vpwr scs8hd_decap_8
XANTENNA__43__A chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_39_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_60_105 vgnd vpwr scs8hd_decap_12
XFILLER_53_8 vgnd vpwr scs8hd_decap_6
XFILLER_45_135 vgnd vpwr scs8hd_decap_8
XANTENNA__38__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_51_46 vgnd vpwr scs8hd_decap_12
XFILLER_42_105 vgnd vpwr scs8hd_decap_12
XFILLER_27_135 vgnd vpwr scs8hd_decap_8
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_84 vgnd vpwr scs8hd_decap_8
XFILLER_46_68 vgnd vpwr scs8hd_decap_12
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_141 vgnd vpwr scs8hd_decap_4
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_43_47 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_3_/S mux_right_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_81 vgnd vpwr scs8hd_decap_6
XFILLER_13_39 vgnd vpwr scs8hd_decap_8
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_60_117 vgnd vpwr scs8hd_decap_12
XFILLER_40_15 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_0.mux_l3_in_0__S mux_right_ipin_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_51_117 vgnd vpwr scs8hd_decap_4
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_51_58 vgnd vpwr scs8hd_decap_3
XFILLER_42_117 vpwr vgnd scs8hd_fill_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_0.scs8hd_buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X left_grid_pin_0_
+ vgnd vpwr scs8hd_buf_1
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
X_39_ chany_top_in[1] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_135 vgnd vpwr scs8hd_decap_8
XFILLER_8_51 vgnd vpwr scs8hd_decap_12
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_119 vgnd vpwr scs8hd_decap_3
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_123 vgnd vpwr scs8hd_decap_12
XFILLER_54_36 vgnd vpwr scs8hd_decap_8
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_126 vgnd vpwr scs8hd_decap_8
XFILLER_44_80 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_60_129 vgnd vpwr scs8hd_decap_12
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_27 vgnd vpwr scs8hd_decap_6
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
X_38_ chany_top_in[2] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XFILLER_11_143 vgnd vpwr scs8hd_decap_3
XFILLER_43_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_8_63 vgnd vpwr scs8hd_decap_12
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_57_135 vgnd vpwr scs8hd_decap_8
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_60_80 vgnd vpwr scs8hd_decap_12
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_54_138 vgnd vpwr scs8hd_decap_8
XFILLER_49_59 vpwr vgnd scs8hd_fill_2
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_8
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_1__S mux_left_ipin_0.mux_l1_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_51_27 vgnd vpwr scs8hd_decap_4
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_33_108 vgnd vpwr scs8hd_decap_12
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__D mux_left_ipin_0.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vgnd vpwr scs8hd_decap_4
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
X_37_ chany_top_in[3] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_104 vgnd vpwr scs8hd_decap_12
XFILLER_8_75 vgnd vpwr scs8hd_decap_12
XFILLER_8_97 vgnd vpwr scs8hd_decap_12
XFILLER_43_39 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vgnd vpwr scs8hd_decap_8
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_4_107 vgnd vpwr scs8hd_decap_12
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_80 vgnd vpwr scs8hd_decap_12
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_50 vpwr vgnd scs8hd_fill_2
XFILLER_44_93 vgnd vpwr scs8hd_decap_12
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_73 vgnd vpwr scs8hd_decap_12
XFILLER_30_51 vpwr vgnd scs8hd_fill_2
XFILLER_55_70 vgnd vpwr scs8hd_decap_12
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__D mux_right_ipin_0.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_117 vgnd vpwr scs8hd_decap_12
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XFILLER_52_93 vpwr vgnd scs8hd_fill_2
XFILLER_52_60 vgnd vpwr scs8hd_decap_12
XFILLER_36_50 vgnd vpwr scs8hd_decap_12
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_145 vgnd vpwr scs8hd_fill_1
X_36_ chany_top_in[4] chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XFILLER_7_116 vgnd vpwr scs8hd_decap_6
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_8_87 vgnd vpwr scs8hd_decap_4
X_19_ chany_bottom_in[1] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_4_119 vgnd vpwr scs8hd_decap_12
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_48_104 vgnd vpwr scs8hd_decap_12
XFILLER_44_50 vgnd vpwr scs8hd_decap_12
XFILLER_60_93 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_49_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_64 vgnd vpwr scs8hd_decap_3
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_93 vgnd vpwr scs8hd_decap_4
XFILLER_55_82 vgnd vpwr scs8hd_decap_3
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_30_85 vgnd vpwr scs8hd_decap_6
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vgnd vpwr scs8hd_decap_3
XFILLER_41_121 vgnd vpwr scs8hd_fill_1
XFILLER_41_110 vgnd vpwr scs8hd_decap_8
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_36_62 vgnd vpwr scs8hd_decap_12
XFILLER_23_143 vgnd vpwr scs8hd_decap_3
XFILLER_23_110 vgnd vpwr scs8hd_decap_12
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_52_72 vgnd vpwr scs8hd_decap_12
X_35_ chany_top_in[5] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_11_135 vgnd vpwr scs8hd_decap_8
XFILLER_22_97 vgnd vpwr scs8hd_decap_12
X_18_ chany_bottom_in[2] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_96 vgnd vpwr scs8hd_decap_12
XFILLER_33_74 vgnd vpwr scs8hd_fill_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l3_in_1__A0 mux_left_ipin_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_58_93 vgnd vpwr scs8hd_decap_12
XFILLER_48_116 vgnd vpwr scs8hd_decap_12
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XFILLER_0_145 vgnd vpwr scs8hd_fill_1
XFILLER_62_141 vgnd vpwr scs8hd_decap_4
XFILLER_44_40 vgnd vpwr scs8hd_fill_1
XFILLER_45_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.mux_l4_in_0__A0 mux_left_ipin_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_76 vgnd vpwr scs8hd_decap_12
XFILLER_44_141 vgnd vpwr scs8hd_decap_4
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.mux_l2_in_2__S mux_left_ipin_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_4
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_86 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_0.scs8hd_dfxbp_1_3_ prog_clk mux_left_ipin_0.mux_l3_in_0_/S mux_left_ipin_0.mux_l4_in_0_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_52_84 vgnd vpwr scs8hd_decap_8
XFILLER_36_74 vgnd vpwr scs8hd_decap_12
X_34_ chany_top_in[6] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_47_51 vgnd vpwr scs8hd_decap_8
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
X_17_ chany_bottom_in[3] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_140 vgnd vpwr scs8hd_decap_6
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.mux_l3_in_1__A1 mux_left_ipin_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_48_128 vgnd vpwr scs8hd_decap_12
XFILLER_54_109 vgnd vpwr scs8hd_decap_12
XFILLER_53_131 vgnd vpwr scs8hd_decap_3
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_30_65 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l4_in_0__A1 mux_left_ipin_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_6
XFILLER_14_88 vgnd vpwr scs8hd_decap_4
XFILLER_50_145 vgnd vpwr scs8hd_fill_1
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XFILLER_41_31 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_98 vgnd vpwr scs8hd_decap_12
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_0.scs8hd_dfxbp_1_2_ prog_clk mux_left_ipin_0.mux_l2_in_1_/S mux_left_ipin_0.mux_l3_in_0_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_145 vgnd vpwr scs8hd_fill_1
XFILLER_2_36 vgnd vpwr scs8hd_decap_8
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
X_33_ chany_top_in[7] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_36_86 vgnd vpwr scs8hd_decap_6
XFILLER_14_145 vgnd vpwr scs8hd_fill_1
XFILLER_3_90 vgnd vpwr scs8hd_decap_4
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
X_16_ chany_bottom_in[4] chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_54 vpwr vgnd scs8hd_fill_2
XFILLER_44_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_2__S mux_right_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_28_21 vgnd vpwr scs8hd_fill_1
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_55_41 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_30_55 vgnd vpwr scs8hd_fill_1
XFILLER_30_44 vgnd vpwr scs8hd_decap_4
XFILLER_50_113 vgnd vpwr scs8hd_decap_12
XFILLER_35_143 vgnd vpwr scs8hd_decap_3
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XPHY_99 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_8
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_0.scs8hd_dfxbp_1_1_ prog_clk mux_left_ipin_0.mux_l1_in_2_/S mux_left_ipin_0.mux_l2_in_1_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XFILLER_6_90 vpwr vgnd scs8hd_fill_2
XPHY_22 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_41_43 vgnd vpwr scs8hd_decap_12
XFILLER_32_113 vgnd vpwr scs8hd_decap_12
XFILLER_17_143 vgnd vpwr scs8hd_decap_3
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
XFILLER_2_48 vgnd vpwr scs8hd_decap_8
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_135 vgnd vpwr scs8hd_decap_8
XFILLER_36_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l3_in_0__S mux_left_ipin_0.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
X_32_ chany_top_in[8] chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
XANTENNA__11__A chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
X_15_ chany_bottom_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_47_97 vgnd vpwr scs8hd_fill_1
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__06__A chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_56_141 vgnd vpwr scs8hd_decap_4
XFILLER_44_32 vgnd vpwr scs8hd_decap_8
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_137 vgnd vpwr scs8hd_decap_8
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_53_144 vpwr vgnd scs8hd_fill_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A0 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_55_53 vgnd vpwr scs8hd_decap_8
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_50_125 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_6_80 vgnd vpwr scs8hd_decap_8
Xmem_left_ipin_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_left_ipin_0.mux_l1_in_2_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_55 vgnd vpwr scs8hd_decap_6
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_32_125 vgnd vpwr scs8hd_decap_12
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XANTENNA__14__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
X_31_ chany_top_in[9] chany_bottom_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A0 mux_right_ipin_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_47_65 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_14_ chany_bottom_in[6] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__22__A chany_top_in[18] vgnd vpwr scs8hd_diode_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_135 vgnd vpwr scs8hd_decap_8
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_71 vpwr vgnd scs8hd_fill_2
XFILLER_0_60 vpwr vgnd scs8hd_fill_2
XANTENNA__17__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_62_145 vgnd vpwr scs8hd_fill_1
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XFILLER_47_120 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l2_in_3_ _02_/HI chany_top_in[16] mux_left_ipin_0.mux_l2_in_1_/S
+ mux_left_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_44_145 vgnd vpwr scs8hd_fill_1
XFILLER_50_137 vgnd vpwr scs8hd_decap_8
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_0__S mux_right_ipin_0.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_26_145 vgnd vpwr scs8hd_fill_1
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__30__A chany_top_in[10] vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A1 mux_right_ipin_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_137 vgnd vpwr scs8hd_decap_8
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XANTENNA__25__A chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_52_99 vgnd vpwr scs8hd_decap_12
XFILLER_20_129 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.mux_l4_in_0_ mux_left_ipin_0.mux_l3_in_1_/X mux_left_ipin_0.mux_l3_in_0_/X
+ mux_left_ipin_0.mux_l4_in_0_/S mux_left_ipin_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
X_30_ chany_top_in[10] chany_bottom_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XFILLER_47_77 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A1 mux_right_ipin_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_7 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
X_13_ chany_bottom_in[7] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_103 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l3_in_1_ mux_left_ipin_0.mux_l2_in_3_/X mux_left_ipin_0.mux_l2_in_2_/X
+ mux_left_ipin_0.mux_l3_in_0_/S mux_left_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XFILLER_28_24 vgnd vpwr scs8hd_decap_6
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__D mux_left_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XANTENNA__33__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_47_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_3__S mux_right_ipin_0.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_left_ipin_0.mux_l2_in_1_/S
+ mux_left_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_59 vgnd vpwr scs8hd_decap_3
XANTENNA__28__A chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_55_66 vpwr vgnd scs8hd_fill_2
XFILLER_30_69 vpwr vgnd scs8hd_fill_2
XFILLER_29_143 vgnd vpwr scs8hd_decap_3
XFILLER_50_105 vgnd vpwr scs8hd_decap_4
XFILLER_35_135 vgnd vpwr scs8hd_decap_8
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XFILLER_17_135 vgnd vpwr scs8hd_decap_8
XFILLER_15_91 vgnd vpwr scs8hd_decap_12
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XANTENNA__41__A chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XFILLER_54_3 vgnd vpwr scs8hd_decap_3
XFILLER_47_89 vgnd vpwr scs8hd_decap_8
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA__36__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_141 vgnd vpwr scs8hd_decap_4
X_12_ chany_bottom_in[8] chany_top_out[8] vgnd vpwr scs8hd_buf_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_decap_3
XFILLER_33_47 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_0.mux_l3_in_0_ mux_left_ipin_0.mux_l2_in_1_/X mux_left_ipin_0.mux_l2_in_0_/X
+ mux_left_ipin_0.mux_l3_in_0_/S mux_left_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_0_40 vgnd vpwr scs8hd_decap_4
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XFILLER_44_68 vgnd vpwr scs8hd_decap_12
XFILLER_53_136 vgnd vpwr scs8hd_decap_8
XFILLER_53_103 vgnd vpwr scs8hd_decap_12
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_0.mux_l2_in_1_ chany_bottom_in[10] mux_left_ipin_0.mux_l1_in_2_/X mux_left_ipin_0.mux_l2_in_1_/S
+ mux_left_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_55_89 vpwr vgnd scs8hd_fill_2
XFILLER_30_48 vgnd vpwr scs8hd_fill_1
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_90 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA__39__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_left_ipin_0.mux_l1_in_2_/S
+ mux_left_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_6
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
X_11_ chany_bottom_in[9] chany_top_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
XFILLER_0_63 vgnd vpwr scs8hd_decap_4
XFILLER_0_52 vgnd vpwr scs8hd_decap_8
XFILLER_60_68 vgnd vpwr scs8hd_decap_12
XFILLER_56_145 vgnd vpwr scs8hd_fill_1
XFILLER_28_15 vgnd vpwr scs8hd_decap_6
XFILLER_47_123 vgnd vpwr scs8hd_decap_12
XFILLER_38_145 vgnd vpwr scs8hd_fill_1
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_0.mux_l2_in_0_ mux_left_ipin_0.mux_l1_in_1_/X mux_left_ipin_0.mux_l1_in_0_/X
+ mux_left_ipin_0.mux_l2_in_1_/S mux_left_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_53_115 vgnd vpwr scs8hd_decap_4
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XFILLER_41_118 vgnd vpwr scs8hd_fill_1
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l3_in_1__S mux_right_ipin_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_0.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_left_ipin_0.mux_l1_in_2_/S
+ mux_left_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_52_36 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_42_80 vgnd vpwr scs8hd_decap_12
XFILLER_3_96 vpwr vgnd scs8hd_fill_2
X_10_ chany_bottom_in[10] chany_top_out[10] vgnd vpwr scs8hd_buf_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_59_143 vgnd vpwr scs8hd_decap_3
XFILLER_59_110 vgnd vpwr scs8hd_decap_12
XFILLER_58_68 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XFILLER_50_80 vgnd vpwr scs8hd_decap_12
XFILLER_47_135 vgnd vpwr scs8hd_decap_8
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_53_127 vpwr vgnd scs8hd_fill_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_102 vgnd vpwr scs8hd_decap_12
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_25 vpwr vgnd scs8hd_fill_2
XFILLER_44_105 vgnd vpwr scs8hd_decap_12
XFILLER_29_135 vgnd vpwr scs8hd_decap_8
XFILLER_26_105 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_left_ipin_0.mux_l1_in_2_/S
+ mux_left_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_141 vgnd vpwr scs8hd_decap_4
XFILLER_31_93 vgnd vpwr scs8hd_fill_1
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XFILLER_52_48 vgnd vpwr scs8hd_decap_12
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_38 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_104 vgnd vpwr scs8hd_decap_12
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_39 vgnd vpwr scs8hd_decap_8
XFILLER_3_107 vgnd vpwr scs8hd_decap_12
XFILLER_48_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_62_117 vgnd vpwr scs8hd_decap_12
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_37 vpwr vgnd scs8hd_fill_2
XFILLER_55_15 vgnd vpwr scs8hd_decap_6
XFILLER_44_117 vgnd vpwr scs8hd_decap_12
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vgnd vpwr scs8hd_decap_8
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
XFILLER_31_50 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_2__S mux_left_ipin_0.mux_l1_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_31_120 vpwr vgnd scs8hd_fill_2
XFILLER_9_135 vgnd vpwr scs8hd_decap_8
XFILLER_42_93 vgnd vpwr scs8hd_decap_12
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_27 vgnd vpwr scs8hd_decap_12
XFILLER_6_116 vgnd vpwr scs8hd_decap_12
XFILLER_10_145 vgnd vpwr scs8hd_fill_1
XFILLER_53_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__D mux_right_ipin_0.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_59_123 vgnd vpwr scs8hd_decap_12
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_119 vgnd vpwr scs8hd_decap_3
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_2_141 vgnd vpwr scs8hd_decap_4
XFILLER_0_11 vgnd vpwr scs8hd_decap_8
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_62_129 vgnd vpwr scs8hd_decap_12
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XFILLER_47_104 vpwr vgnd scs8hd_fill_2
XFILLER_34_61 vgnd vpwr scs8hd_decap_12
XFILLER_34_50 vpwr vgnd scs8hd_fill_2
XFILLER_50_93 vgnd vpwr scs8hd_decap_12
XFILLER_44_129 vgnd vpwr scs8hd_decap_12
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_45_71 vpwr vgnd scs8hd_fill_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_129 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A0 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_31_143 vgnd vpwr scs8hd_decap_3
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_121 vgnd vpwr scs8hd_decap_12
XFILLER_3_66 vgnd vpwr scs8hd_decap_12
XFILLER_13_121 vgnd vpwr scs8hd_fill_1
XFILLER_13_143 vgnd vpwr scs8hd_decap_3
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_47_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_1__A0 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_53_60 vgnd vpwr scs8hd_fill_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_128 vgnd vpwr scs8hd_decap_12
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_59_135 vgnd vpwr scs8hd_decap_8
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
XFILLER_56_105 vgnd vpwr scs8hd_decap_12
XFILLER_48_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_0.mux_l3_in_0__A0 mux_left_ipin_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_74 vgnd vpwr scs8hd_decap_12
XFILLER_53_119 vgnd vpwr scs8hd_fill_1
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_34_73 vgnd vpwr scs8hd_decap_12
XFILLER_45_50 vgnd vpwr scs8hd_fill_1
XFILLER_29_62 vpwr vgnd scs8hd_fill_2
XFILLER_41_19 vgnd vpwr scs8hd_fill_1
XFILLER_34_141 vgnd vpwr scs8hd_decap_4
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_31_96 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XFILLER_56_93 vgnd vpwr scs8hd_decap_12
XFILLER_31_100 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_141 vgnd vpwr scs8hd_decap_4
.ends

