VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__2_
  CLASS BLOCK ;
  FOREIGN sb_2__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 138.000 ;
  PIN bottom_left_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END bottom_left_grid_pin_34_
  PIN bottom_left_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 2.400 ;
    END
  END bottom_left_grid_pin_35_
  PIN bottom_left_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END bottom_left_grid_pin_36_
  PIN bottom_left_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.400 ;
    END
  END bottom_left_grid_pin_37_
  PIN bottom_left_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.400 ;
    END
  END bottom_left_grid_pin_38_
  PIN bottom_left_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 2.400 ;
    END
  END bottom_left_grid_pin_39_
  PIN bottom_left_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END bottom_left_grid_pin_40_
  PIN bottom_left_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END bottom_left_grid_pin_41_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.400 ;
    END
  END bottom_right_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 116.320 140.000 116.920 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 2.400 12.200 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.400 29.200 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 2.400 32.600 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 2.400 104.000 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 2.400 107.400 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 2.400 114.200 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 2.400 117.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 2.400 121.000 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 2.400 124.400 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 2.400 127.800 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 2.400 134.600 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 2.400 76.800 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.400 93.800 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 2.400 97.200 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chany_bottom_out[9]
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 2.400 138.000 ;
    END
  END left_top_grid_pin_1_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.160 140.000 23.760 ;
    END
  END prog_clk
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 1.450 2.760 134.320 128.080 ;
      LAYER met2 ;
        RECT 1.480 2.680 138.370 137.885 ;
        RECT 2.030 1.515 3.950 2.680 ;
        RECT 4.790 1.515 6.710 2.680 ;
        RECT 7.550 1.515 9.470 2.680 ;
        RECT 10.310 1.515 12.230 2.680 ;
        RECT 13.070 1.515 15.450 2.680 ;
        RECT 16.290 1.515 18.210 2.680 ;
        RECT 19.050 1.515 20.970 2.680 ;
        RECT 21.810 1.515 23.730 2.680 ;
        RECT 24.570 1.515 26.490 2.680 ;
        RECT 27.330 1.515 29.710 2.680 ;
        RECT 30.550 1.515 32.470 2.680 ;
        RECT 33.310 1.515 35.230 2.680 ;
        RECT 36.070 1.515 37.990 2.680 ;
        RECT 38.830 1.515 40.750 2.680 ;
        RECT 41.590 1.515 43.970 2.680 ;
        RECT 44.810 1.515 46.730 2.680 ;
        RECT 47.570 1.515 49.490 2.680 ;
        RECT 50.330 1.515 52.250 2.680 ;
        RECT 53.090 1.515 55.010 2.680 ;
        RECT 55.850 1.515 58.230 2.680 ;
        RECT 59.070 1.515 60.990 2.680 ;
        RECT 61.830 1.515 63.750 2.680 ;
        RECT 64.590 1.515 66.510 2.680 ;
        RECT 67.350 1.515 69.270 2.680 ;
        RECT 70.110 1.515 72.490 2.680 ;
        RECT 73.330 1.515 75.250 2.680 ;
        RECT 76.090 1.515 78.010 2.680 ;
        RECT 78.850 1.515 80.770 2.680 ;
        RECT 81.610 1.515 83.530 2.680 ;
        RECT 84.370 1.515 86.750 2.680 ;
        RECT 87.590 1.515 89.510 2.680 ;
        RECT 90.350 1.515 92.270 2.680 ;
        RECT 93.110 1.515 95.030 2.680 ;
        RECT 95.870 1.515 97.790 2.680 ;
        RECT 98.630 1.515 101.010 2.680 ;
        RECT 101.850 1.515 103.770 2.680 ;
        RECT 104.610 1.515 106.530 2.680 ;
        RECT 107.370 1.515 109.290 2.680 ;
        RECT 110.130 1.515 112.050 2.680 ;
        RECT 112.890 1.515 115.270 2.680 ;
        RECT 116.110 1.515 118.030 2.680 ;
        RECT 118.870 1.515 120.790 2.680 ;
        RECT 121.630 1.515 123.550 2.680 ;
        RECT 124.390 1.515 126.310 2.680 ;
        RECT 127.150 1.515 129.530 2.680 ;
        RECT 130.370 1.515 132.290 2.680 ;
        RECT 133.130 1.515 135.050 2.680 ;
        RECT 135.890 1.515 137.810 2.680 ;
      LAYER met3 ;
        RECT 2.800 137.000 138.395 137.865 ;
        RECT 2.400 135.000 138.395 137.000 ;
        RECT 2.800 133.600 138.395 135.000 ;
        RECT 2.400 131.600 138.395 133.600 ;
        RECT 2.800 130.200 138.395 131.600 ;
        RECT 2.400 128.200 138.395 130.200 ;
        RECT 2.800 126.800 138.395 128.200 ;
        RECT 2.400 124.800 138.395 126.800 ;
        RECT 2.800 123.400 138.395 124.800 ;
        RECT 2.400 121.400 138.395 123.400 ;
        RECT 2.800 120.000 138.395 121.400 ;
        RECT 2.400 118.000 138.395 120.000 ;
        RECT 2.800 117.320 138.395 118.000 ;
        RECT 2.800 116.600 137.200 117.320 ;
        RECT 2.400 115.920 137.200 116.600 ;
        RECT 2.400 114.600 138.395 115.920 ;
        RECT 2.800 113.200 138.395 114.600 ;
        RECT 2.400 111.200 138.395 113.200 ;
        RECT 2.800 109.800 138.395 111.200 ;
        RECT 2.400 107.800 138.395 109.800 ;
        RECT 2.800 106.400 138.395 107.800 ;
        RECT 2.400 104.400 138.395 106.400 ;
        RECT 2.800 103.000 138.395 104.400 ;
        RECT 2.400 101.000 138.395 103.000 ;
        RECT 2.800 99.600 138.395 101.000 ;
        RECT 2.400 97.600 138.395 99.600 ;
        RECT 2.800 96.200 138.395 97.600 ;
        RECT 2.400 94.200 138.395 96.200 ;
        RECT 2.800 92.800 138.395 94.200 ;
        RECT 2.400 90.800 138.395 92.800 ;
        RECT 2.800 89.400 138.395 90.800 ;
        RECT 2.400 87.400 138.395 89.400 ;
        RECT 2.800 86.000 138.395 87.400 ;
        RECT 2.400 84.000 138.395 86.000 ;
        RECT 2.800 82.600 138.395 84.000 ;
        RECT 2.400 80.600 138.395 82.600 ;
        RECT 2.800 79.200 138.395 80.600 ;
        RECT 2.400 77.200 138.395 79.200 ;
        RECT 2.800 75.800 138.395 77.200 ;
        RECT 2.400 73.800 138.395 75.800 ;
        RECT 2.800 72.400 138.395 73.800 ;
        RECT 2.400 70.400 138.395 72.400 ;
        RECT 2.800 69.000 137.200 70.400 ;
        RECT 2.400 67.000 138.395 69.000 ;
        RECT 2.800 65.600 138.395 67.000 ;
        RECT 2.400 63.600 138.395 65.600 ;
        RECT 2.800 62.200 138.395 63.600 ;
        RECT 2.400 60.200 138.395 62.200 ;
        RECT 2.800 58.800 138.395 60.200 ;
        RECT 2.400 56.800 138.395 58.800 ;
        RECT 2.800 55.400 138.395 56.800 ;
        RECT 2.400 53.400 138.395 55.400 ;
        RECT 2.800 52.000 138.395 53.400 ;
        RECT 2.400 50.000 138.395 52.000 ;
        RECT 2.800 48.600 138.395 50.000 ;
        RECT 2.400 46.600 138.395 48.600 ;
        RECT 2.800 45.200 138.395 46.600 ;
        RECT 2.400 43.200 138.395 45.200 ;
        RECT 2.800 41.800 138.395 43.200 ;
        RECT 2.400 39.800 138.395 41.800 ;
        RECT 2.800 38.400 138.395 39.800 ;
        RECT 2.400 36.400 138.395 38.400 ;
        RECT 2.800 35.000 138.395 36.400 ;
        RECT 2.400 33.000 138.395 35.000 ;
        RECT 2.800 31.600 138.395 33.000 ;
        RECT 2.400 29.600 138.395 31.600 ;
        RECT 2.800 28.200 138.395 29.600 ;
        RECT 2.400 26.200 138.395 28.200 ;
        RECT 2.800 24.800 138.395 26.200 ;
        RECT 2.400 24.160 138.395 24.800 ;
        RECT 2.400 22.800 137.200 24.160 ;
        RECT 2.800 22.760 137.200 22.800 ;
        RECT 2.800 21.400 138.395 22.760 ;
        RECT 2.400 19.400 138.395 21.400 ;
        RECT 2.800 18.000 138.395 19.400 ;
        RECT 2.400 16.000 138.395 18.000 ;
        RECT 2.800 14.600 138.395 16.000 ;
        RECT 2.400 12.600 138.395 14.600 ;
        RECT 2.800 11.200 138.395 12.600 ;
        RECT 2.400 9.200 138.395 11.200 ;
        RECT 2.800 7.800 138.395 9.200 ;
        RECT 2.400 5.800 138.395 7.800 ;
        RECT 2.800 4.400 138.395 5.800 ;
        RECT 2.400 2.400 138.395 4.400 ;
        RECT 2.800 1.535 138.395 2.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_2__2_
END LIBRARY

