VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__1_
  CLASS BLOCK ;
  FOREIGN cbx_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 80.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 2.400 ;
    END
  END address[5]
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 2.400 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 2.400 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 2.400 ;
    END
  END bottom_grid_pin_8_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 2.400 6.760 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.400 11.520 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.400 29.200 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 2.400 51.640 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 2.400 78.160 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 2.080 200.000 2.680 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 6.160 200.000 6.760 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 10.920 200.000 11.520 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 15.000 200.000 15.600 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 19.760 200.000 20.360 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 23.840 200.000 24.440 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 28.600 200.000 29.200 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 32.680 200.000 33.280 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 37.440 200.000 38.040 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 42.200 200.000 42.800 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 46.280 200.000 46.880 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 51.040 200.000 51.640 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 55.120 200.000 55.720 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 59.880 200.000 60.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 63.960 200.000 64.560 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 68.720 200.000 69.320 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 72.800 200.000 73.400 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 77.560 200.000 78.160 ;
    END
  END chanx_right_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END enable
  PIN top_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.610 77.600 166.890 80.000 ;
    END
  END top_grid_pin_14_
  PIN top_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.210 77.600 33.490 80.000 ;
    END
  END top_grid_pin_2_
  PIN top_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.910 77.600 100.190 80.000 ;
    END
  END top_grid_pin_6_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 38.055 10.640 39.655 68.240 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 71.385 10.640 72.985 68.240 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 68.085 ;
      LAYER met1 ;
        RECT 5.520 0.040 194.120 68.240 ;
      LAYER met2 ;
        RECT 7.000 77.320 32.930 78.045 ;
        RECT 33.770 77.320 99.630 78.045 ;
        RECT 100.470 77.320 166.330 78.045 ;
        RECT 167.170 77.320 190.810 78.045 ;
        RECT 7.000 2.680 190.810 77.320 ;
        RECT 7.000 0.010 8.550 2.680 ;
        RECT 9.390 0.010 26.490 2.680 ;
        RECT 27.330 0.010 44.890 2.680 ;
        RECT 45.730 0.010 62.830 2.680 ;
        RECT 63.670 0.010 81.230 2.680 ;
        RECT 82.070 0.010 99.170 2.680 ;
        RECT 100.010 0.010 117.570 2.680 ;
        RECT 118.410 0.010 135.510 2.680 ;
        RECT 136.350 0.010 153.910 2.680 ;
        RECT 154.750 0.010 171.850 2.680 ;
        RECT 172.690 0.010 190.250 2.680 ;
      LAYER met3 ;
        RECT 2.800 77.160 197.200 78.025 ;
        RECT 2.400 73.800 197.600 77.160 ;
        RECT 2.800 72.400 197.200 73.800 ;
        RECT 2.400 69.720 197.600 72.400 ;
        RECT 2.800 68.320 197.200 69.720 ;
        RECT 2.400 64.960 197.600 68.320 ;
        RECT 2.800 63.560 197.200 64.960 ;
        RECT 2.400 60.880 197.600 63.560 ;
        RECT 2.800 59.480 197.200 60.880 ;
        RECT 2.400 56.120 197.600 59.480 ;
        RECT 2.800 54.720 197.200 56.120 ;
        RECT 2.400 52.040 197.600 54.720 ;
        RECT 2.800 50.640 197.200 52.040 ;
        RECT 2.400 47.280 197.600 50.640 ;
        RECT 2.800 45.880 197.200 47.280 ;
        RECT 2.400 43.200 197.600 45.880 ;
        RECT 2.800 41.800 197.200 43.200 ;
        RECT 2.400 38.440 197.600 41.800 ;
        RECT 2.800 37.040 197.200 38.440 ;
        RECT 2.400 33.680 197.600 37.040 ;
        RECT 2.800 32.280 197.200 33.680 ;
        RECT 2.400 29.600 197.600 32.280 ;
        RECT 2.800 28.200 197.200 29.600 ;
        RECT 2.400 24.840 197.600 28.200 ;
        RECT 2.800 23.440 197.200 24.840 ;
        RECT 2.400 20.760 197.600 23.440 ;
        RECT 2.800 19.360 197.200 20.760 ;
        RECT 2.400 16.000 197.600 19.360 ;
        RECT 2.800 14.600 197.200 16.000 ;
        RECT 2.400 11.920 197.600 14.600 ;
        RECT 2.800 10.520 197.200 11.920 ;
        RECT 2.400 7.160 197.600 10.520 ;
        RECT 2.800 5.760 197.200 7.160 ;
        RECT 2.400 3.080 197.600 5.760 ;
        RECT 2.800 1.680 197.200 3.080 ;
        RECT 2.400 0.175 197.600 1.680 ;
      LAYER met4 ;
        RECT 13.670 10.240 37.655 68.240 ;
        RECT 40.055 10.240 70.985 68.240 ;
        RECT 73.385 10.240 172.985 68.240 ;
        RECT 13.670 0.175 172.985 10.240 ;
      LAYER met5 ;
        RECT 13.460 17.900 145.700 19.500 ;
  END
END cbx_1__1_
END LIBRARY

