magic
tech EFS8A
magscale 1 2
timestamp 1602874355
<< locali >>
rect 9873 18071 9907 18241
rect 10695 11305 10701 11339
rect 10695 11237 10729 11305
rect 10511 3689 10517 3723
rect 10511 3621 10545 3689
<< viali >>
rect 11437 97801 11471 97835
rect 11253 97597 11287 97631
rect 11805 97597 11839 97631
rect 11345 94945 11379 94979
rect 11161 94877 11195 94911
rect 11529 94809 11563 94843
rect 11161 94537 11195 94571
rect 11529 94265 11563 94299
rect 11713 85289 11747 85323
rect 11529 85153 11563 85187
rect 11529 84745 11563 84779
rect 11805 80937 11839 80971
rect 11161 80801 11195 80835
rect 11345 80733 11379 80767
rect 11161 80393 11195 80427
rect 11529 80053 11563 80087
rect 11437 71689 11471 71723
rect 11253 71485 11287 71519
rect 11805 71485 11839 71519
rect 11805 66793 11839 66827
rect 11161 66657 11195 66691
rect 11345 66589 11379 66623
rect 11253 66249 11287 66283
rect 11529 65977 11563 66011
rect 11437 58633 11471 58667
rect 11253 58429 11287 58463
rect 11805 58429 11839 58463
rect 11805 53737 11839 53771
rect 11161 53601 11195 53635
rect 11345 53533 11379 53567
rect 11253 53193 11287 53227
rect 11621 52853 11655 52887
rect 11713 45033 11747 45067
rect 11529 44897 11563 44931
rect 11529 44489 11563 44523
rect 10793 40137 10827 40171
rect 11529 40137 11563 40171
rect 10885 40001 10919 40035
rect 11069 39933 11103 39967
rect 10977 39253 11011 39287
rect 11437 31433 11471 31467
rect 11253 31229 11287 31263
rect 11805 31229 11839 31263
rect 10793 27081 10827 27115
rect 11253 27081 11287 27115
rect 10885 26945 10919 26979
rect 11069 26877 11103 26911
rect 10885 26197 10919 26231
rect 11253 19465 11287 19499
rect 10333 19261 10367 19295
rect 10695 19193 10729 19227
rect 10241 19125 10275 19159
rect 11621 18921 11655 18955
rect 11022 18853 11056 18887
rect 10701 18717 10735 18751
rect 8585 18581 8619 18615
rect 10333 18581 10367 18615
rect 9413 18377 9447 18411
rect 11161 18377 11195 18411
rect 11805 18377 11839 18411
rect 9873 18241 9907 18275
rect 8493 18173 8527 18207
rect 8401 18105 8435 18139
rect 8855 18105 8889 18139
rect 10241 18173 10275 18207
rect 10562 18105 10596 18139
rect 9689 18037 9723 18071
rect 9873 18037 9907 18071
rect 10149 18037 10183 18071
rect 11437 18037 11471 18071
rect 11069 17833 11103 17867
rect 10511 17765 10545 17799
rect 10149 17629 10183 17663
rect 8677 17493 8711 17527
rect 10793 17289 10827 17323
rect 11437 17221 11471 17255
rect 8677 17085 8711 17119
rect 9137 17085 9171 17119
rect 9689 17085 9723 17119
rect 9873 17085 9907 17119
rect 11253 17085 11287 17119
rect 11805 17085 11839 17119
rect 8217 16949 8251 16983
rect 8493 16949 8527 16983
rect 8769 16949 8803 16983
rect 10517 16949 10551 16983
rect 11621 16745 11655 16779
rect 11022 16677 11056 16711
rect 10701 16541 10735 16575
rect 9045 16473 9079 16507
rect 8769 16405 8803 16439
rect 11069 16201 11103 16235
rect 10241 16133 10275 16167
rect 8033 16065 8067 16099
rect 8861 15997 8895 16031
rect 9321 15997 9355 16031
rect 9781 15997 9815 16031
rect 10057 15997 10091 16031
rect 8309 15929 8343 15963
rect 8769 15861 8803 15895
rect 10701 15861 10735 15895
rect 8217 15657 8251 15691
rect 9965 15657 9999 15691
rect 8401 15589 8435 15623
rect 8769 15589 8803 15623
rect 9505 15589 9539 15623
rect 9873 15589 9907 15623
rect 10057 15589 10091 15623
rect 10425 15589 10459 15623
rect 8309 15521 8343 15555
rect 8033 15453 8067 15487
rect 9689 15453 9723 15487
rect 9045 15317 9079 15351
rect 10701 15317 10735 15351
rect 7389 15113 7423 15147
rect 8125 15113 8159 15147
rect 9965 15113 9999 15147
rect 10333 15113 10367 15147
rect 8493 14977 8527 15011
rect 9689 14977 9723 15011
rect 10517 14977 10551 15011
rect 11253 14977 11287 15011
rect 8861 14909 8895 14943
rect 9137 14909 9171 14943
rect 10701 14909 10735 14943
rect 7757 14841 7791 14875
rect 8953 14841 8987 14875
rect 9321 14841 9355 14875
rect 10885 14841 10919 14875
rect 11529 14841 11563 14875
rect 9229 14773 9263 14807
rect 10793 14773 10827 14807
rect 9137 14569 9171 14603
rect 10701 14501 10735 14535
rect 8125 14433 8159 14467
rect 9505 14433 9539 14467
rect 9781 14433 9815 14467
rect 8769 14365 8803 14399
rect 9689 14365 9723 14399
rect 8033 13685 8067 13719
rect 8953 13685 8987 13719
rect 9781 13685 9815 13719
rect 10057 13685 10091 13719
rect 11805 13481 11839 13515
rect 11161 13345 11195 13379
rect 11345 13277 11379 13311
rect 11161 12937 11195 12971
rect 8217 12733 8251 12767
rect 8861 12665 8895 12699
rect 7941 12597 7975 12631
rect 11529 12597 11563 12631
rect 8769 12053 8803 12087
rect 8677 11713 8711 11747
rect 8769 11645 8803 11679
rect 9229 11645 9263 11679
rect 9597 11645 9631 11679
rect 9965 11645 9999 11679
rect 8309 11577 8343 11611
rect 10149 11509 10183 11543
rect 10701 11305 10735 11339
rect 11253 11305 11287 11339
rect 10333 11169 10367 11203
rect 8861 10965 8895 10999
rect 10701 10761 10735 10795
rect 10333 10421 10367 10455
rect 11437 4233 11471 4267
rect 9413 4165 9447 4199
rect 9229 4029 9263 4063
rect 11253 4029 11287 4063
rect 9781 3893 9815 3927
rect 11805 3893 11839 3927
rect 8677 3689 8711 3723
rect 10517 3689 10551 3723
rect 10149 3485 10183 3519
rect 11069 3349 11103 3383
rect 8125 3009 8159 3043
rect 10057 3009 10091 3043
rect 10701 3009 10735 3043
rect 8585 2941 8619 2975
rect 9045 2941 9079 2975
rect 9413 2941 9447 2975
rect 9781 2941 9815 2975
rect 8401 2805 8435 2839
rect 10425 2805 10459 2839
rect 10977 2601 11011 2635
rect 11713 2601 11747 2635
rect 10609 2465 10643 2499
rect 11253 2465 11287 2499
rect 11069 2397 11103 2431
rect 8585 2261 8619 2295
<< metal1 >>
rect 1104 106650 12880 106672
rect 1104 106598 3315 106650
rect 3367 106598 3379 106650
rect 3431 106598 3443 106650
rect 3495 106598 3507 106650
rect 3559 106598 7982 106650
rect 8034 106598 8046 106650
rect 8098 106598 8110 106650
rect 8162 106598 8174 106650
rect 8226 106598 12880 106650
rect 1104 106576 12880 106598
rect 1104 106106 12880 106128
rect 1104 106054 5648 106106
rect 5700 106054 5712 106106
rect 5764 106054 5776 106106
rect 5828 106054 5840 106106
rect 5892 106054 10315 106106
rect 10367 106054 10379 106106
rect 10431 106054 10443 106106
rect 10495 106054 10507 106106
rect 10559 106054 12880 106106
rect 1104 106032 12880 106054
rect 1104 105562 12880 105584
rect 1104 105510 3315 105562
rect 3367 105510 3379 105562
rect 3431 105510 3443 105562
rect 3495 105510 3507 105562
rect 3559 105510 7982 105562
rect 8034 105510 8046 105562
rect 8098 105510 8110 105562
rect 8162 105510 8174 105562
rect 8226 105510 12880 105562
rect 1104 105488 12880 105510
rect 1104 105018 12880 105040
rect 1104 104966 5648 105018
rect 5700 104966 5712 105018
rect 5764 104966 5776 105018
rect 5828 104966 5840 105018
rect 5892 104966 10315 105018
rect 10367 104966 10379 105018
rect 10431 104966 10443 105018
rect 10495 104966 10507 105018
rect 10559 104966 12880 105018
rect 1104 104944 12880 104966
rect 1104 104474 12880 104496
rect 1104 104422 3315 104474
rect 3367 104422 3379 104474
rect 3431 104422 3443 104474
rect 3495 104422 3507 104474
rect 3559 104422 7982 104474
rect 8034 104422 8046 104474
rect 8098 104422 8110 104474
rect 8162 104422 8174 104474
rect 8226 104422 12880 104474
rect 1104 104400 12880 104422
rect 1104 103930 12880 103952
rect 1104 103878 5648 103930
rect 5700 103878 5712 103930
rect 5764 103878 5776 103930
rect 5828 103878 5840 103930
rect 5892 103878 10315 103930
rect 10367 103878 10379 103930
rect 10431 103878 10443 103930
rect 10495 103878 10507 103930
rect 10559 103878 12880 103930
rect 1104 103856 12880 103878
rect 1104 103386 12880 103408
rect 1104 103334 3315 103386
rect 3367 103334 3379 103386
rect 3431 103334 3443 103386
rect 3495 103334 3507 103386
rect 3559 103334 7982 103386
rect 8034 103334 8046 103386
rect 8098 103334 8110 103386
rect 8162 103334 8174 103386
rect 8226 103334 12880 103386
rect 1104 103312 12880 103334
rect 1104 102842 12880 102864
rect 1104 102790 5648 102842
rect 5700 102790 5712 102842
rect 5764 102790 5776 102842
rect 5828 102790 5840 102842
rect 5892 102790 10315 102842
rect 10367 102790 10379 102842
rect 10431 102790 10443 102842
rect 10495 102790 10507 102842
rect 10559 102790 12880 102842
rect 1104 102768 12880 102790
rect 1104 102298 12880 102320
rect 1104 102246 3315 102298
rect 3367 102246 3379 102298
rect 3431 102246 3443 102298
rect 3495 102246 3507 102298
rect 3559 102246 7982 102298
rect 8034 102246 8046 102298
rect 8098 102246 8110 102298
rect 8162 102246 8174 102298
rect 8226 102246 12880 102298
rect 1104 102224 12880 102246
rect 1104 101754 12880 101776
rect 1104 101702 5648 101754
rect 5700 101702 5712 101754
rect 5764 101702 5776 101754
rect 5828 101702 5840 101754
rect 5892 101702 10315 101754
rect 10367 101702 10379 101754
rect 10431 101702 10443 101754
rect 10495 101702 10507 101754
rect 10559 101702 12880 101754
rect 1104 101680 12880 101702
rect 1104 101210 12880 101232
rect 1104 101158 3315 101210
rect 3367 101158 3379 101210
rect 3431 101158 3443 101210
rect 3495 101158 3507 101210
rect 3559 101158 7982 101210
rect 8034 101158 8046 101210
rect 8098 101158 8110 101210
rect 8162 101158 8174 101210
rect 8226 101158 12880 101210
rect 1104 101136 12880 101158
rect 1104 100666 12880 100688
rect 1104 100614 5648 100666
rect 5700 100614 5712 100666
rect 5764 100614 5776 100666
rect 5828 100614 5840 100666
rect 5892 100614 10315 100666
rect 10367 100614 10379 100666
rect 10431 100614 10443 100666
rect 10495 100614 10507 100666
rect 10559 100614 12880 100666
rect 1104 100592 12880 100614
rect 1104 100122 12880 100144
rect 1104 100070 3315 100122
rect 3367 100070 3379 100122
rect 3431 100070 3443 100122
rect 3495 100070 3507 100122
rect 3559 100070 7982 100122
rect 8034 100070 8046 100122
rect 8098 100070 8110 100122
rect 8162 100070 8174 100122
rect 8226 100070 12880 100122
rect 1104 100048 12880 100070
rect 1104 99578 12880 99600
rect 1104 99526 5648 99578
rect 5700 99526 5712 99578
rect 5764 99526 5776 99578
rect 5828 99526 5840 99578
rect 5892 99526 10315 99578
rect 10367 99526 10379 99578
rect 10431 99526 10443 99578
rect 10495 99526 10507 99578
rect 10559 99526 12880 99578
rect 1104 99504 12880 99526
rect 1104 99034 12880 99056
rect 1104 98982 3315 99034
rect 3367 98982 3379 99034
rect 3431 98982 3443 99034
rect 3495 98982 3507 99034
rect 3559 98982 7982 99034
rect 8034 98982 8046 99034
rect 8098 98982 8110 99034
rect 8162 98982 8174 99034
rect 8226 98982 12880 99034
rect 1104 98960 12880 98982
rect 1104 98490 12880 98512
rect 1104 98438 5648 98490
rect 5700 98438 5712 98490
rect 5764 98438 5776 98490
rect 5828 98438 5840 98490
rect 5892 98438 10315 98490
rect 10367 98438 10379 98490
rect 10431 98438 10443 98490
rect 10495 98438 10507 98490
rect 10559 98438 12880 98490
rect 1104 98416 12880 98438
rect 1104 97946 12880 97968
rect 1104 97894 3315 97946
rect 3367 97894 3379 97946
rect 3431 97894 3443 97946
rect 3495 97894 3507 97946
rect 3559 97894 7982 97946
rect 8034 97894 8046 97946
rect 8098 97894 8110 97946
rect 8162 97894 8174 97946
rect 8226 97894 12880 97946
rect 1104 97872 12880 97894
rect 11422 97832 11428 97844
rect 11383 97804 11428 97832
rect 11422 97792 11428 97804
rect 11480 97792 11486 97844
rect 11238 97628 11244 97640
rect 11199 97600 11244 97628
rect 11238 97588 11244 97600
rect 11296 97628 11302 97640
rect 11793 97631 11851 97637
rect 11793 97628 11805 97631
rect 11296 97600 11805 97628
rect 11296 97588 11302 97600
rect 11793 97597 11805 97600
rect 11839 97597 11851 97631
rect 11793 97591 11851 97597
rect 1104 97402 12880 97424
rect 1104 97350 5648 97402
rect 5700 97350 5712 97402
rect 5764 97350 5776 97402
rect 5828 97350 5840 97402
rect 5892 97350 10315 97402
rect 10367 97350 10379 97402
rect 10431 97350 10443 97402
rect 10495 97350 10507 97402
rect 10559 97350 12880 97402
rect 1104 97328 12880 97350
rect 1104 96858 12880 96880
rect 1104 96806 3315 96858
rect 3367 96806 3379 96858
rect 3431 96806 3443 96858
rect 3495 96806 3507 96858
rect 3559 96806 7982 96858
rect 8034 96806 8046 96858
rect 8098 96806 8110 96858
rect 8162 96806 8174 96858
rect 8226 96806 12880 96858
rect 1104 96784 12880 96806
rect 1104 96314 12880 96336
rect 1104 96262 5648 96314
rect 5700 96262 5712 96314
rect 5764 96262 5776 96314
rect 5828 96262 5840 96314
rect 5892 96262 10315 96314
rect 10367 96262 10379 96314
rect 10431 96262 10443 96314
rect 10495 96262 10507 96314
rect 10559 96262 12880 96314
rect 1104 96240 12880 96262
rect 1104 95770 12880 95792
rect 1104 95718 3315 95770
rect 3367 95718 3379 95770
rect 3431 95718 3443 95770
rect 3495 95718 3507 95770
rect 3559 95718 7982 95770
rect 8034 95718 8046 95770
rect 8098 95718 8110 95770
rect 8162 95718 8174 95770
rect 8226 95718 12880 95770
rect 1104 95696 12880 95718
rect 1104 95226 12880 95248
rect 1104 95174 5648 95226
rect 5700 95174 5712 95226
rect 5764 95174 5776 95226
rect 5828 95174 5840 95226
rect 5892 95174 10315 95226
rect 10367 95174 10379 95226
rect 10431 95174 10443 95226
rect 10495 95174 10507 95226
rect 10559 95174 12880 95226
rect 1104 95152 12880 95174
rect 11054 94936 11060 94988
rect 11112 94976 11118 94988
rect 11333 94979 11391 94985
rect 11333 94976 11345 94979
rect 11112 94948 11345 94976
rect 11112 94936 11118 94948
rect 11333 94945 11345 94948
rect 11379 94945 11391 94979
rect 11333 94939 11391 94945
rect 11146 94908 11152 94920
rect 11107 94880 11152 94908
rect 11146 94868 11152 94880
rect 11204 94868 11210 94920
rect 11238 94800 11244 94852
rect 11296 94840 11302 94852
rect 11517 94843 11575 94849
rect 11517 94840 11529 94843
rect 11296 94812 11529 94840
rect 11296 94800 11302 94812
rect 11517 94809 11529 94812
rect 11563 94809 11575 94843
rect 11517 94803 11575 94809
rect 1104 94682 12880 94704
rect 1104 94630 3315 94682
rect 3367 94630 3379 94682
rect 3431 94630 3443 94682
rect 3495 94630 3507 94682
rect 3559 94630 7982 94682
rect 8034 94630 8046 94682
rect 8098 94630 8110 94682
rect 8162 94630 8174 94682
rect 8226 94630 12880 94682
rect 1104 94608 12880 94630
rect 11146 94568 11152 94580
rect 11107 94540 11152 94568
rect 11146 94528 11152 94540
rect 11204 94528 11210 94580
rect 11054 94256 11060 94308
rect 11112 94296 11118 94308
rect 11517 94299 11575 94305
rect 11517 94296 11529 94299
rect 11112 94268 11529 94296
rect 11112 94256 11118 94268
rect 11517 94265 11529 94268
rect 11563 94265 11575 94299
rect 11517 94259 11575 94265
rect 1104 94138 12880 94160
rect 1104 94086 5648 94138
rect 5700 94086 5712 94138
rect 5764 94086 5776 94138
rect 5828 94086 5840 94138
rect 5892 94086 10315 94138
rect 10367 94086 10379 94138
rect 10431 94086 10443 94138
rect 10495 94086 10507 94138
rect 10559 94086 12880 94138
rect 1104 94064 12880 94086
rect 1104 93594 12880 93616
rect 1104 93542 3315 93594
rect 3367 93542 3379 93594
rect 3431 93542 3443 93594
rect 3495 93542 3507 93594
rect 3559 93542 7982 93594
rect 8034 93542 8046 93594
rect 8098 93542 8110 93594
rect 8162 93542 8174 93594
rect 8226 93542 12880 93594
rect 1104 93520 12880 93542
rect 1104 93050 12880 93072
rect 1104 92998 5648 93050
rect 5700 92998 5712 93050
rect 5764 92998 5776 93050
rect 5828 92998 5840 93050
rect 5892 92998 10315 93050
rect 10367 92998 10379 93050
rect 10431 92998 10443 93050
rect 10495 92998 10507 93050
rect 10559 92998 12880 93050
rect 1104 92976 12880 92998
rect 1104 92506 12880 92528
rect 1104 92454 3315 92506
rect 3367 92454 3379 92506
rect 3431 92454 3443 92506
rect 3495 92454 3507 92506
rect 3559 92454 7982 92506
rect 8034 92454 8046 92506
rect 8098 92454 8110 92506
rect 8162 92454 8174 92506
rect 8226 92454 12880 92506
rect 1104 92432 12880 92454
rect 1104 91962 12880 91984
rect 1104 91910 5648 91962
rect 5700 91910 5712 91962
rect 5764 91910 5776 91962
rect 5828 91910 5840 91962
rect 5892 91910 10315 91962
rect 10367 91910 10379 91962
rect 10431 91910 10443 91962
rect 10495 91910 10507 91962
rect 10559 91910 12880 91962
rect 1104 91888 12880 91910
rect 1104 91418 12880 91440
rect 1104 91366 3315 91418
rect 3367 91366 3379 91418
rect 3431 91366 3443 91418
rect 3495 91366 3507 91418
rect 3559 91366 7982 91418
rect 8034 91366 8046 91418
rect 8098 91366 8110 91418
rect 8162 91366 8174 91418
rect 8226 91366 12880 91418
rect 1104 91344 12880 91366
rect 1104 90874 12880 90896
rect 1104 90822 5648 90874
rect 5700 90822 5712 90874
rect 5764 90822 5776 90874
rect 5828 90822 5840 90874
rect 5892 90822 10315 90874
rect 10367 90822 10379 90874
rect 10431 90822 10443 90874
rect 10495 90822 10507 90874
rect 10559 90822 12880 90874
rect 1104 90800 12880 90822
rect 1104 90330 12880 90352
rect 1104 90278 3315 90330
rect 3367 90278 3379 90330
rect 3431 90278 3443 90330
rect 3495 90278 3507 90330
rect 3559 90278 7982 90330
rect 8034 90278 8046 90330
rect 8098 90278 8110 90330
rect 8162 90278 8174 90330
rect 8226 90278 12880 90330
rect 1104 90256 12880 90278
rect 1104 89786 12880 89808
rect 1104 89734 5648 89786
rect 5700 89734 5712 89786
rect 5764 89734 5776 89786
rect 5828 89734 5840 89786
rect 5892 89734 10315 89786
rect 10367 89734 10379 89786
rect 10431 89734 10443 89786
rect 10495 89734 10507 89786
rect 10559 89734 12880 89786
rect 1104 89712 12880 89734
rect 1104 89242 12880 89264
rect 1104 89190 3315 89242
rect 3367 89190 3379 89242
rect 3431 89190 3443 89242
rect 3495 89190 3507 89242
rect 3559 89190 7982 89242
rect 8034 89190 8046 89242
rect 8098 89190 8110 89242
rect 8162 89190 8174 89242
rect 8226 89190 12880 89242
rect 1104 89168 12880 89190
rect 1104 88698 12880 88720
rect 1104 88646 5648 88698
rect 5700 88646 5712 88698
rect 5764 88646 5776 88698
rect 5828 88646 5840 88698
rect 5892 88646 10315 88698
rect 10367 88646 10379 88698
rect 10431 88646 10443 88698
rect 10495 88646 10507 88698
rect 10559 88646 12880 88698
rect 1104 88624 12880 88646
rect 1104 88154 12880 88176
rect 1104 88102 3315 88154
rect 3367 88102 3379 88154
rect 3431 88102 3443 88154
rect 3495 88102 3507 88154
rect 3559 88102 7982 88154
rect 8034 88102 8046 88154
rect 8098 88102 8110 88154
rect 8162 88102 8174 88154
rect 8226 88102 12880 88154
rect 1104 88080 12880 88102
rect 1104 87610 12880 87632
rect 1104 87558 5648 87610
rect 5700 87558 5712 87610
rect 5764 87558 5776 87610
rect 5828 87558 5840 87610
rect 5892 87558 10315 87610
rect 10367 87558 10379 87610
rect 10431 87558 10443 87610
rect 10495 87558 10507 87610
rect 10559 87558 12880 87610
rect 1104 87536 12880 87558
rect 1104 87066 12880 87088
rect 1104 87014 3315 87066
rect 3367 87014 3379 87066
rect 3431 87014 3443 87066
rect 3495 87014 3507 87066
rect 3559 87014 7982 87066
rect 8034 87014 8046 87066
rect 8098 87014 8110 87066
rect 8162 87014 8174 87066
rect 8226 87014 12880 87066
rect 1104 86992 12880 87014
rect 1104 86522 12880 86544
rect 1104 86470 5648 86522
rect 5700 86470 5712 86522
rect 5764 86470 5776 86522
rect 5828 86470 5840 86522
rect 5892 86470 10315 86522
rect 10367 86470 10379 86522
rect 10431 86470 10443 86522
rect 10495 86470 10507 86522
rect 10559 86470 12880 86522
rect 1104 86448 12880 86470
rect 1104 85978 12880 86000
rect 1104 85926 3315 85978
rect 3367 85926 3379 85978
rect 3431 85926 3443 85978
rect 3495 85926 3507 85978
rect 3559 85926 7982 85978
rect 8034 85926 8046 85978
rect 8098 85926 8110 85978
rect 8162 85926 8174 85978
rect 8226 85926 12880 85978
rect 1104 85904 12880 85926
rect 1104 85434 12880 85456
rect 1104 85382 5648 85434
rect 5700 85382 5712 85434
rect 5764 85382 5776 85434
rect 5828 85382 5840 85434
rect 5892 85382 10315 85434
rect 10367 85382 10379 85434
rect 10431 85382 10443 85434
rect 10495 85382 10507 85434
rect 10559 85382 12880 85434
rect 1104 85360 12880 85382
rect 10686 85280 10692 85332
rect 10744 85320 10750 85332
rect 11701 85323 11759 85329
rect 11701 85320 11713 85323
rect 10744 85292 11713 85320
rect 10744 85280 10750 85292
rect 11701 85289 11713 85292
rect 11747 85289 11759 85323
rect 11701 85283 11759 85289
rect 11514 85184 11520 85196
rect 11475 85156 11520 85184
rect 11514 85144 11520 85156
rect 11572 85144 11578 85196
rect 1104 84890 12880 84912
rect 1104 84838 3315 84890
rect 3367 84838 3379 84890
rect 3431 84838 3443 84890
rect 3495 84838 3507 84890
rect 3559 84838 7982 84890
rect 8034 84838 8046 84890
rect 8098 84838 8110 84890
rect 8162 84838 8174 84890
rect 8226 84838 12880 84890
rect 1104 84816 12880 84838
rect 11514 84776 11520 84788
rect 11475 84748 11520 84776
rect 11514 84736 11520 84748
rect 11572 84776 11578 84788
rect 11790 84776 11796 84788
rect 11572 84748 11796 84776
rect 11572 84736 11578 84748
rect 11790 84736 11796 84748
rect 11848 84736 11854 84788
rect 1104 84346 12880 84368
rect 1104 84294 5648 84346
rect 5700 84294 5712 84346
rect 5764 84294 5776 84346
rect 5828 84294 5840 84346
rect 5892 84294 10315 84346
rect 10367 84294 10379 84346
rect 10431 84294 10443 84346
rect 10495 84294 10507 84346
rect 10559 84294 12880 84346
rect 1104 84272 12880 84294
rect 1104 83802 12880 83824
rect 1104 83750 3315 83802
rect 3367 83750 3379 83802
rect 3431 83750 3443 83802
rect 3495 83750 3507 83802
rect 3559 83750 7982 83802
rect 8034 83750 8046 83802
rect 8098 83750 8110 83802
rect 8162 83750 8174 83802
rect 8226 83750 12880 83802
rect 1104 83728 12880 83750
rect 1104 83258 12880 83280
rect 1104 83206 5648 83258
rect 5700 83206 5712 83258
rect 5764 83206 5776 83258
rect 5828 83206 5840 83258
rect 5892 83206 10315 83258
rect 10367 83206 10379 83258
rect 10431 83206 10443 83258
rect 10495 83206 10507 83258
rect 10559 83206 12880 83258
rect 1104 83184 12880 83206
rect 1104 82714 12880 82736
rect 1104 82662 3315 82714
rect 3367 82662 3379 82714
rect 3431 82662 3443 82714
rect 3495 82662 3507 82714
rect 3559 82662 7982 82714
rect 8034 82662 8046 82714
rect 8098 82662 8110 82714
rect 8162 82662 8174 82714
rect 8226 82662 12880 82714
rect 1104 82640 12880 82662
rect 1104 82170 12880 82192
rect 1104 82118 5648 82170
rect 5700 82118 5712 82170
rect 5764 82118 5776 82170
rect 5828 82118 5840 82170
rect 5892 82118 10315 82170
rect 10367 82118 10379 82170
rect 10431 82118 10443 82170
rect 10495 82118 10507 82170
rect 10559 82118 12880 82170
rect 1104 82096 12880 82118
rect 1104 81626 12880 81648
rect 1104 81574 3315 81626
rect 3367 81574 3379 81626
rect 3431 81574 3443 81626
rect 3495 81574 3507 81626
rect 3559 81574 7982 81626
rect 8034 81574 8046 81626
rect 8098 81574 8110 81626
rect 8162 81574 8174 81626
rect 8226 81574 12880 81626
rect 1104 81552 12880 81574
rect 1104 81082 12880 81104
rect 1104 81030 5648 81082
rect 5700 81030 5712 81082
rect 5764 81030 5776 81082
rect 5828 81030 5840 81082
rect 5892 81030 10315 81082
rect 10367 81030 10379 81082
rect 10431 81030 10443 81082
rect 10495 81030 10507 81082
rect 10559 81030 12880 81082
rect 1104 81008 12880 81030
rect 11790 80968 11796 80980
rect 11751 80940 11796 80968
rect 11790 80928 11796 80940
rect 11848 80928 11854 80980
rect 11146 80832 11152 80844
rect 11107 80804 11152 80832
rect 11146 80792 11152 80804
rect 11204 80792 11210 80844
rect 11330 80764 11336 80776
rect 11291 80736 11336 80764
rect 11330 80724 11336 80736
rect 11388 80724 11394 80776
rect 1104 80538 12880 80560
rect 1104 80486 3315 80538
rect 3367 80486 3379 80538
rect 3431 80486 3443 80538
rect 3495 80486 3507 80538
rect 3559 80486 7982 80538
rect 8034 80486 8046 80538
rect 8098 80486 8110 80538
rect 8162 80486 8174 80538
rect 8226 80486 12880 80538
rect 1104 80464 12880 80486
rect 11146 80424 11152 80436
rect 11107 80396 11152 80424
rect 11146 80384 11152 80396
rect 11204 80384 11210 80436
rect 11146 80044 11152 80096
rect 11204 80084 11210 80096
rect 11330 80084 11336 80096
rect 11204 80056 11336 80084
rect 11204 80044 11210 80056
rect 11330 80044 11336 80056
rect 11388 80084 11394 80096
rect 11517 80087 11575 80093
rect 11517 80084 11529 80087
rect 11388 80056 11529 80084
rect 11388 80044 11394 80056
rect 11517 80053 11529 80056
rect 11563 80053 11575 80087
rect 11517 80047 11575 80053
rect 1104 79994 12880 80016
rect 1104 79942 5648 79994
rect 5700 79942 5712 79994
rect 5764 79942 5776 79994
rect 5828 79942 5840 79994
rect 5892 79942 10315 79994
rect 10367 79942 10379 79994
rect 10431 79942 10443 79994
rect 10495 79942 10507 79994
rect 10559 79942 12880 79994
rect 1104 79920 12880 79942
rect 1104 79450 12880 79472
rect 1104 79398 3315 79450
rect 3367 79398 3379 79450
rect 3431 79398 3443 79450
rect 3495 79398 3507 79450
rect 3559 79398 7982 79450
rect 8034 79398 8046 79450
rect 8098 79398 8110 79450
rect 8162 79398 8174 79450
rect 8226 79398 12880 79450
rect 1104 79376 12880 79398
rect 1104 78906 12880 78928
rect 1104 78854 5648 78906
rect 5700 78854 5712 78906
rect 5764 78854 5776 78906
rect 5828 78854 5840 78906
rect 5892 78854 10315 78906
rect 10367 78854 10379 78906
rect 10431 78854 10443 78906
rect 10495 78854 10507 78906
rect 10559 78854 12880 78906
rect 1104 78832 12880 78854
rect 1104 78362 12880 78384
rect 1104 78310 3315 78362
rect 3367 78310 3379 78362
rect 3431 78310 3443 78362
rect 3495 78310 3507 78362
rect 3559 78310 7982 78362
rect 8034 78310 8046 78362
rect 8098 78310 8110 78362
rect 8162 78310 8174 78362
rect 8226 78310 12880 78362
rect 1104 78288 12880 78310
rect 1104 77818 12880 77840
rect 1104 77766 5648 77818
rect 5700 77766 5712 77818
rect 5764 77766 5776 77818
rect 5828 77766 5840 77818
rect 5892 77766 10315 77818
rect 10367 77766 10379 77818
rect 10431 77766 10443 77818
rect 10495 77766 10507 77818
rect 10559 77766 12880 77818
rect 1104 77744 12880 77766
rect 1104 77274 12880 77296
rect 1104 77222 3315 77274
rect 3367 77222 3379 77274
rect 3431 77222 3443 77274
rect 3495 77222 3507 77274
rect 3559 77222 7982 77274
rect 8034 77222 8046 77274
rect 8098 77222 8110 77274
rect 8162 77222 8174 77274
rect 8226 77222 12880 77274
rect 1104 77200 12880 77222
rect 1104 76730 12880 76752
rect 1104 76678 5648 76730
rect 5700 76678 5712 76730
rect 5764 76678 5776 76730
rect 5828 76678 5840 76730
rect 5892 76678 10315 76730
rect 10367 76678 10379 76730
rect 10431 76678 10443 76730
rect 10495 76678 10507 76730
rect 10559 76678 12880 76730
rect 1104 76656 12880 76678
rect 1104 76186 12880 76208
rect 1104 76134 3315 76186
rect 3367 76134 3379 76186
rect 3431 76134 3443 76186
rect 3495 76134 3507 76186
rect 3559 76134 7982 76186
rect 8034 76134 8046 76186
rect 8098 76134 8110 76186
rect 8162 76134 8174 76186
rect 8226 76134 12880 76186
rect 1104 76112 12880 76134
rect 1104 75642 12880 75664
rect 1104 75590 5648 75642
rect 5700 75590 5712 75642
rect 5764 75590 5776 75642
rect 5828 75590 5840 75642
rect 5892 75590 10315 75642
rect 10367 75590 10379 75642
rect 10431 75590 10443 75642
rect 10495 75590 10507 75642
rect 10559 75590 12880 75642
rect 1104 75568 12880 75590
rect 1104 75098 12880 75120
rect 1104 75046 3315 75098
rect 3367 75046 3379 75098
rect 3431 75046 3443 75098
rect 3495 75046 3507 75098
rect 3559 75046 7982 75098
rect 8034 75046 8046 75098
rect 8098 75046 8110 75098
rect 8162 75046 8174 75098
rect 8226 75046 12880 75098
rect 1104 75024 12880 75046
rect 1104 74554 12880 74576
rect 1104 74502 5648 74554
rect 5700 74502 5712 74554
rect 5764 74502 5776 74554
rect 5828 74502 5840 74554
rect 5892 74502 10315 74554
rect 10367 74502 10379 74554
rect 10431 74502 10443 74554
rect 10495 74502 10507 74554
rect 10559 74502 12880 74554
rect 1104 74480 12880 74502
rect 1104 74010 12880 74032
rect 1104 73958 3315 74010
rect 3367 73958 3379 74010
rect 3431 73958 3443 74010
rect 3495 73958 3507 74010
rect 3559 73958 7982 74010
rect 8034 73958 8046 74010
rect 8098 73958 8110 74010
rect 8162 73958 8174 74010
rect 8226 73958 12880 74010
rect 1104 73936 12880 73958
rect 1104 73466 12880 73488
rect 1104 73414 5648 73466
rect 5700 73414 5712 73466
rect 5764 73414 5776 73466
rect 5828 73414 5840 73466
rect 5892 73414 10315 73466
rect 10367 73414 10379 73466
rect 10431 73414 10443 73466
rect 10495 73414 10507 73466
rect 10559 73414 12880 73466
rect 1104 73392 12880 73414
rect 1104 72922 12880 72944
rect 1104 72870 3315 72922
rect 3367 72870 3379 72922
rect 3431 72870 3443 72922
rect 3495 72870 3507 72922
rect 3559 72870 7982 72922
rect 8034 72870 8046 72922
rect 8098 72870 8110 72922
rect 8162 72870 8174 72922
rect 8226 72870 12880 72922
rect 1104 72848 12880 72870
rect 1104 72378 12880 72400
rect 1104 72326 5648 72378
rect 5700 72326 5712 72378
rect 5764 72326 5776 72378
rect 5828 72326 5840 72378
rect 5892 72326 10315 72378
rect 10367 72326 10379 72378
rect 10431 72326 10443 72378
rect 10495 72326 10507 72378
rect 10559 72326 12880 72378
rect 1104 72304 12880 72326
rect 1104 71834 12880 71856
rect 1104 71782 3315 71834
rect 3367 71782 3379 71834
rect 3431 71782 3443 71834
rect 3495 71782 3507 71834
rect 3559 71782 7982 71834
rect 8034 71782 8046 71834
rect 8098 71782 8110 71834
rect 8162 71782 8174 71834
rect 8226 71782 12880 71834
rect 1104 71760 12880 71782
rect 10962 71680 10968 71732
rect 11020 71720 11026 71732
rect 11425 71723 11483 71729
rect 11425 71720 11437 71723
rect 11020 71692 11437 71720
rect 11020 71680 11026 71692
rect 11425 71689 11437 71692
rect 11471 71689 11483 71723
rect 11425 71683 11483 71689
rect 11238 71516 11244 71528
rect 11199 71488 11244 71516
rect 11238 71476 11244 71488
rect 11296 71516 11302 71528
rect 11790 71516 11796 71528
rect 11296 71488 11796 71516
rect 11296 71476 11302 71488
rect 11790 71476 11796 71488
rect 11848 71476 11854 71528
rect 1104 71290 12880 71312
rect 1104 71238 5648 71290
rect 5700 71238 5712 71290
rect 5764 71238 5776 71290
rect 5828 71238 5840 71290
rect 5892 71238 10315 71290
rect 10367 71238 10379 71290
rect 10431 71238 10443 71290
rect 10495 71238 10507 71290
rect 10559 71238 12880 71290
rect 1104 71216 12880 71238
rect 1104 70746 12880 70768
rect 1104 70694 3315 70746
rect 3367 70694 3379 70746
rect 3431 70694 3443 70746
rect 3495 70694 3507 70746
rect 3559 70694 7982 70746
rect 8034 70694 8046 70746
rect 8098 70694 8110 70746
rect 8162 70694 8174 70746
rect 8226 70694 12880 70746
rect 1104 70672 12880 70694
rect 1104 70202 12880 70224
rect 1104 70150 5648 70202
rect 5700 70150 5712 70202
rect 5764 70150 5776 70202
rect 5828 70150 5840 70202
rect 5892 70150 10315 70202
rect 10367 70150 10379 70202
rect 10431 70150 10443 70202
rect 10495 70150 10507 70202
rect 10559 70150 12880 70202
rect 1104 70128 12880 70150
rect 1104 69658 12880 69680
rect 1104 69606 3315 69658
rect 3367 69606 3379 69658
rect 3431 69606 3443 69658
rect 3495 69606 3507 69658
rect 3559 69606 7982 69658
rect 8034 69606 8046 69658
rect 8098 69606 8110 69658
rect 8162 69606 8174 69658
rect 8226 69606 12880 69658
rect 1104 69584 12880 69606
rect 1104 69114 12880 69136
rect 1104 69062 5648 69114
rect 5700 69062 5712 69114
rect 5764 69062 5776 69114
rect 5828 69062 5840 69114
rect 5892 69062 10315 69114
rect 10367 69062 10379 69114
rect 10431 69062 10443 69114
rect 10495 69062 10507 69114
rect 10559 69062 12880 69114
rect 1104 69040 12880 69062
rect 1104 68570 12880 68592
rect 1104 68518 3315 68570
rect 3367 68518 3379 68570
rect 3431 68518 3443 68570
rect 3495 68518 3507 68570
rect 3559 68518 7982 68570
rect 8034 68518 8046 68570
rect 8098 68518 8110 68570
rect 8162 68518 8174 68570
rect 8226 68518 12880 68570
rect 1104 68496 12880 68518
rect 1104 68026 12880 68048
rect 1104 67974 5648 68026
rect 5700 67974 5712 68026
rect 5764 67974 5776 68026
rect 5828 67974 5840 68026
rect 5892 67974 10315 68026
rect 10367 67974 10379 68026
rect 10431 67974 10443 68026
rect 10495 67974 10507 68026
rect 10559 67974 12880 68026
rect 1104 67952 12880 67974
rect 1104 67482 12880 67504
rect 1104 67430 3315 67482
rect 3367 67430 3379 67482
rect 3431 67430 3443 67482
rect 3495 67430 3507 67482
rect 3559 67430 7982 67482
rect 8034 67430 8046 67482
rect 8098 67430 8110 67482
rect 8162 67430 8174 67482
rect 8226 67430 12880 67482
rect 1104 67408 12880 67430
rect 1104 66938 12880 66960
rect 1104 66886 5648 66938
rect 5700 66886 5712 66938
rect 5764 66886 5776 66938
rect 5828 66886 5840 66938
rect 5892 66886 10315 66938
rect 10367 66886 10379 66938
rect 10431 66886 10443 66938
rect 10495 66886 10507 66938
rect 10559 66886 12880 66938
rect 1104 66864 12880 66886
rect 11790 66824 11796 66836
rect 11751 66796 11796 66824
rect 11790 66784 11796 66796
rect 11848 66784 11854 66836
rect 11149 66691 11207 66697
rect 11149 66657 11161 66691
rect 11195 66688 11207 66691
rect 11422 66688 11428 66700
rect 11195 66660 11428 66688
rect 11195 66657 11207 66660
rect 11149 66651 11207 66657
rect 11422 66648 11428 66660
rect 11480 66648 11486 66700
rect 11330 66620 11336 66632
rect 11291 66592 11336 66620
rect 11330 66580 11336 66592
rect 11388 66580 11394 66632
rect 1104 66394 12880 66416
rect 1104 66342 3315 66394
rect 3367 66342 3379 66394
rect 3431 66342 3443 66394
rect 3495 66342 3507 66394
rect 3559 66342 7982 66394
rect 8034 66342 8046 66394
rect 8098 66342 8110 66394
rect 8162 66342 8174 66394
rect 8226 66342 12880 66394
rect 1104 66320 12880 66342
rect 11241 66283 11299 66289
rect 11241 66249 11253 66283
rect 11287 66280 11299 66283
rect 11422 66280 11428 66292
rect 11287 66252 11428 66280
rect 11287 66249 11299 66252
rect 11241 66243 11299 66249
rect 11422 66240 11428 66252
rect 11480 66240 11486 66292
rect 10134 65968 10140 66020
rect 10192 66008 10198 66020
rect 11330 66008 11336 66020
rect 10192 65980 11336 66008
rect 10192 65968 10198 65980
rect 11330 65968 11336 65980
rect 11388 66008 11394 66020
rect 11517 66011 11575 66017
rect 11517 66008 11529 66011
rect 11388 65980 11529 66008
rect 11388 65968 11394 65980
rect 11517 65977 11529 65980
rect 11563 65977 11575 66011
rect 11517 65971 11575 65977
rect 1104 65850 12880 65872
rect 1104 65798 5648 65850
rect 5700 65798 5712 65850
rect 5764 65798 5776 65850
rect 5828 65798 5840 65850
rect 5892 65798 10315 65850
rect 10367 65798 10379 65850
rect 10431 65798 10443 65850
rect 10495 65798 10507 65850
rect 10559 65798 12880 65850
rect 1104 65776 12880 65798
rect 1104 65306 12880 65328
rect 1104 65254 3315 65306
rect 3367 65254 3379 65306
rect 3431 65254 3443 65306
rect 3495 65254 3507 65306
rect 3559 65254 7982 65306
rect 8034 65254 8046 65306
rect 8098 65254 8110 65306
rect 8162 65254 8174 65306
rect 8226 65254 12880 65306
rect 1104 65232 12880 65254
rect 1104 64762 12880 64784
rect 1104 64710 5648 64762
rect 5700 64710 5712 64762
rect 5764 64710 5776 64762
rect 5828 64710 5840 64762
rect 5892 64710 10315 64762
rect 10367 64710 10379 64762
rect 10431 64710 10443 64762
rect 10495 64710 10507 64762
rect 10559 64710 12880 64762
rect 1104 64688 12880 64710
rect 1104 64218 12880 64240
rect 1104 64166 3315 64218
rect 3367 64166 3379 64218
rect 3431 64166 3443 64218
rect 3495 64166 3507 64218
rect 3559 64166 7982 64218
rect 8034 64166 8046 64218
rect 8098 64166 8110 64218
rect 8162 64166 8174 64218
rect 8226 64166 12880 64218
rect 1104 64144 12880 64166
rect 1104 63674 12880 63696
rect 1104 63622 5648 63674
rect 5700 63622 5712 63674
rect 5764 63622 5776 63674
rect 5828 63622 5840 63674
rect 5892 63622 10315 63674
rect 10367 63622 10379 63674
rect 10431 63622 10443 63674
rect 10495 63622 10507 63674
rect 10559 63622 12880 63674
rect 1104 63600 12880 63622
rect 1104 63130 12880 63152
rect 1104 63078 3315 63130
rect 3367 63078 3379 63130
rect 3431 63078 3443 63130
rect 3495 63078 3507 63130
rect 3559 63078 7982 63130
rect 8034 63078 8046 63130
rect 8098 63078 8110 63130
rect 8162 63078 8174 63130
rect 8226 63078 12880 63130
rect 1104 63056 12880 63078
rect 1104 62586 12880 62608
rect 1104 62534 5648 62586
rect 5700 62534 5712 62586
rect 5764 62534 5776 62586
rect 5828 62534 5840 62586
rect 5892 62534 10315 62586
rect 10367 62534 10379 62586
rect 10431 62534 10443 62586
rect 10495 62534 10507 62586
rect 10559 62534 12880 62586
rect 1104 62512 12880 62534
rect 1104 62042 12880 62064
rect 1104 61990 3315 62042
rect 3367 61990 3379 62042
rect 3431 61990 3443 62042
rect 3495 61990 3507 62042
rect 3559 61990 7982 62042
rect 8034 61990 8046 62042
rect 8098 61990 8110 62042
rect 8162 61990 8174 62042
rect 8226 61990 12880 62042
rect 1104 61968 12880 61990
rect 1104 61498 12880 61520
rect 1104 61446 5648 61498
rect 5700 61446 5712 61498
rect 5764 61446 5776 61498
rect 5828 61446 5840 61498
rect 5892 61446 10315 61498
rect 10367 61446 10379 61498
rect 10431 61446 10443 61498
rect 10495 61446 10507 61498
rect 10559 61446 12880 61498
rect 1104 61424 12880 61446
rect 1104 60954 12880 60976
rect 1104 60902 3315 60954
rect 3367 60902 3379 60954
rect 3431 60902 3443 60954
rect 3495 60902 3507 60954
rect 3559 60902 7982 60954
rect 8034 60902 8046 60954
rect 8098 60902 8110 60954
rect 8162 60902 8174 60954
rect 8226 60902 12880 60954
rect 1104 60880 12880 60902
rect 1104 60410 12880 60432
rect 1104 60358 5648 60410
rect 5700 60358 5712 60410
rect 5764 60358 5776 60410
rect 5828 60358 5840 60410
rect 5892 60358 10315 60410
rect 10367 60358 10379 60410
rect 10431 60358 10443 60410
rect 10495 60358 10507 60410
rect 10559 60358 12880 60410
rect 1104 60336 12880 60358
rect 1104 59866 12880 59888
rect 1104 59814 3315 59866
rect 3367 59814 3379 59866
rect 3431 59814 3443 59866
rect 3495 59814 3507 59866
rect 3559 59814 7982 59866
rect 8034 59814 8046 59866
rect 8098 59814 8110 59866
rect 8162 59814 8174 59866
rect 8226 59814 12880 59866
rect 1104 59792 12880 59814
rect 1104 59322 12880 59344
rect 1104 59270 5648 59322
rect 5700 59270 5712 59322
rect 5764 59270 5776 59322
rect 5828 59270 5840 59322
rect 5892 59270 10315 59322
rect 10367 59270 10379 59322
rect 10431 59270 10443 59322
rect 10495 59270 10507 59322
rect 10559 59270 12880 59322
rect 1104 59248 12880 59270
rect 1104 58778 12880 58800
rect 1104 58726 3315 58778
rect 3367 58726 3379 58778
rect 3431 58726 3443 58778
rect 3495 58726 3507 58778
rect 3559 58726 7982 58778
rect 8034 58726 8046 58778
rect 8098 58726 8110 58778
rect 8162 58726 8174 58778
rect 8226 58726 12880 58778
rect 1104 58704 12880 58726
rect 11422 58664 11428 58676
rect 11383 58636 11428 58664
rect 11422 58624 11428 58636
rect 11480 58624 11486 58676
rect 11238 58460 11244 58472
rect 11199 58432 11244 58460
rect 11238 58420 11244 58432
rect 11296 58460 11302 58472
rect 11790 58460 11796 58472
rect 11296 58432 11796 58460
rect 11296 58420 11302 58432
rect 11790 58420 11796 58432
rect 11848 58420 11854 58472
rect 1104 58234 12880 58256
rect 1104 58182 5648 58234
rect 5700 58182 5712 58234
rect 5764 58182 5776 58234
rect 5828 58182 5840 58234
rect 5892 58182 10315 58234
rect 10367 58182 10379 58234
rect 10431 58182 10443 58234
rect 10495 58182 10507 58234
rect 10559 58182 12880 58234
rect 1104 58160 12880 58182
rect 1104 57690 12880 57712
rect 1104 57638 3315 57690
rect 3367 57638 3379 57690
rect 3431 57638 3443 57690
rect 3495 57638 3507 57690
rect 3559 57638 7982 57690
rect 8034 57638 8046 57690
rect 8098 57638 8110 57690
rect 8162 57638 8174 57690
rect 8226 57638 12880 57690
rect 1104 57616 12880 57638
rect 1104 57146 12880 57168
rect 1104 57094 5648 57146
rect 5700 57094 5712 57146
rect 5764 57094 5776 57146
rect 5828 57094 5840 57146
rect 5892 57094 10315 57146
rect 10367 57094 10379 57146
rect 10431 57094 10443 57146
rect 10495 57094 10507 57146
rect 10559 57094 12880 57146
rect 1104 57072 12880 57094
rect 1104 56602 12880 56624
rect 1104 56550 3315 56602
rect 3367 56550 3379 56602
rect 3431 56550 3443 56602
rect 3495 56550 3507 56602
rect 3559 56550 7982 56602
rect 8034 56550 8046 56602
rect 8098 56550 8110 56602
rect 8162 56550 8174 56602
rect 8226 56550 12880 56602
rect 1104 56528 12880 56550
rect 1104 56058 12880 56080
rect 1104 56006 5648 56058
rect 5700 56006 5712 56058
rect 5764 56006 5776 56058
rect 5828 56006 5840 56058
rect 5892 56006 10315 56058
rect 10367 56006 10379 56058
rect 10431 56006 10443 56058
rect 10495 56006 10507 56058
rect 10559 56006 12880 56058
rect 1104 55984 12880 56006
rect 1104 55514 12880 55536
rect 1104 55462 3315 55514
rect 3367 55462 3379 55514
rect 3431 55462 3443 55514
rect 3495 55462 3507 55514
rect 3559 55462 7982 55514
rect 8034 55462 8046 55514
rect 8098 55462 8110 55514
rect 8162 55462 8174 55514
rect 8226 55462 12880 55514
rect 1104 55440 12880 55462
rect 1104 54970 12880 54992
rect 1104 54918 5648 54970
rect 5700 54918 5712 54970
rect 5764 54918 5776 54970
rect 5828 54918 5840 54970
rect 5892 54918 10315 54970
rect 10367 54918 10379 54970
rect 10431 54918 10443 54970
rect 10495 54918 10507 54970
rect 10559 54918 12880 54970
rect 1104 54896 12880 54918
rect 1104 54426 12880 54448
rect 1104 54374 3315 54426
rect 3367 54374 3379 54426
rect 3431 54374 3443 54426
rect 3495 54374 3507 54426
rect 3559 54374 7982 54426
rect 8034 54374 8046 54426
rect 8098 54374 8110 54426
rect 8162 54374 8174 54426
rect 8226 54374 12880 54426
rect 1104 54352 12880 54374
rect 1104 53882 12880 53904
rect 1104 53830 5648 53882
rect 5700 53830 5712 53882
rect 5764 53830 5776 53882
rect 5828 53830 5840 53882
rect 5892 53830 10315 53882
rect 10367 53830 10379 53882
rect 10431 53830 10443 53882
rect 10495 53830 10507 53882
rect 10559 53830 12880 53882
rect 1104 53808 12880 53830
rect 11790 53768 11796 53780
rect 11751 53740 11796 53768
rect 11790 53728 11796 53740
rect 11848 53728 11854 53780
rect 11149 53635 11207 53641
rect 11149 53601 11161 53635
rect 11195 53632 11207 53635
rect 11422 53632 11428 53644
rect 11195 53604 11428 53632
rect 11195 53601 11207 53604
rect 11149 53595 11207 53601
rect 11422 53592 11428 53604
rect 11480 53592 11486 53644
rect 11333 53567 11391 53573
rect 11333 53533 11345 53567
rect 11379 53564 11391 53567
rect 11606 53564 11612 53576
rect 11379 53536 11612 53564
rect 11379 53533 11391 53536
rect 11333 53527 11391 53533
rect 11606 53524 11612 53536
rect 11664 53524 11670 53576
rect 1104 53338 12880 53360
rect 1104 53286 3315 53338
rect 3367 53286 3379 53338
rect 3431 53286 3443 53338
rect 3495 53286 3507 53338
rect 3559 53286 7982 53338
rect 8034 53286 8046 53338
rect 8098 53286 8110 53338
rect 8162 53286 8174 53338
rect 8226 53286 12880 53338
rect 1104 53264 12880 53286
rect 11241 53227 11299 53233
rect 11241 53193 11253 53227
rect 11287 53224 11299 53227
rect 11422 53224 11428 53236
rect 11287 53196 11428 53224
rect 11287 53193 11299 53196
rect 11241 53187 11299 53193
rect 11422 53184 11428 53196
rect 11480 53184 11486 53236
rect 11606 52884 11612 52896
rect 11567 52856 11612 52884
rect 11606 52844 11612 52856
rect 11664 52844 11670 52896
rect 1104 52794 12880 52816
rect 1104 52742 5648 52794
rect 5700 52742 5712 52794
rect 5764 52742 5776 52794
rect 5828 52742 5840 52794
rect 5892 52742 10315 52794
rect 10367 52742 10379 52794
rect 10431 52742 10443 52794
rect 10495 52742 10507 52794
rect 10559 52742 12880 52794
rect 1104 52720 12880 52742
rect 1104 52250 12880 52272
rect 1104 52198 3315 52250
rect 3367 52198 3379 52250
rect 3431 52198 3443 52250
rect 3495 52198 3507 52250
rect 3559 52198 7982 52250
rect 8034 52198 8046 52250
rect 8098 52198 8110 52250
rect 8162 52198 8174 52250
rect 8226 52198 12880 52250
rect 1104 52176 12880 52198
rect 1104 51706 12880 51728
rect 1104 51654 5648 51706
rect 5700 51654 5712 51706
rect 5764 51654 5776 51706
rect 5828 51654 5840 51706
rect 5892 51654 10315 51706
rect 10367 51654 10379 51706
rect 10431 51654 10443 51706
rect 10495 51654 10507 51706
rect 10559 51654 12880 51706
rect 1104 51632 12880 51654
rect 1104 51162 12880 51184
rect 1104 51110 3315 51162
rect 3367 51110 3379 51162
rect 3431 51110 3443 51162
rect 3495 51110 3507 51162
rect 3559 51110 7982 51162
rect 8034 51110 8046 51162
rect 8098 51110 8110 51162
rect 8162 51110 8174 51162
rect 8226 51110 12880 51162
rect 1104 51088 12880 51110
rect 1104 50618 12880 50640
rect 1104 50566 5648 50618
rect 5700 50566 5712 50618
rect 5764 50566 5776 50618
rect 5828 50566 5840 50618
rect 5892 50566 10315 50618
rect 10367 50566 10379 50618
rect 10431 50566 10443 50618
rect 10495 50566 10507 50618
rect 10559 50566 12880 50618
rect 1104 50544 12880 50566
rect 1104 50074 12880 50096
rect 1104 50022 3315 50074
rect 3367 50022 3379 50074
rect 3431 50022 3443 50074
rect 3495 50022 3507 50074
rect 3559 50022 7982 50074
rect 8034 50022 8046 50074
rect 8098 50022 8110 50074
rect 8162 50022 8174 50074
rect 8226 50022 12880 50074
rect 1104 50000 12880 50022
rect 1104 49530 12880 49552
rect 1104 49478 5648 49530
rect 5700 49478 5712 49530
rect 5764 49478 5776 49530
rect 5828 49478 5840 49530
rect 5892 49478 10315 49530
rect 10367 49478 10379 49530
rect 10431 49478 10443 49530
rect 10495 49478 10507 49530
rect 10559 49478 12880 49530
rect 1104 49456 12880 49478
rect 1104 48986 12880 49008
rect 1104 48934 3315 48986
rect 3367 48934 3379 48986
rect 3431 48934 3443 48986
rect 3495 48934 3507 48986
rect 3559 48934 7982 48986
rect 8034 48934 8046 48986
rect 8098 48934 8110 48986
rect 8162 48934 8174 48986
rect 8226 48934 12880 48986
rect 1104 48912 12880 48934
rect 1104 48442 12880 48464
rect 1104 48390 5648 48442
rect 5700 48390 5712 48442
rect 5764 48390 5776 48442
rect 5828 48390 5840 48442
rect 5892 48390 10315 48442
rect 10367 48390 10379 48442
rect 10431 48390 10443 48442
rect 10495 48390 10507 48442
rect 10559 48390 12880 48442
rect 1104 48368 12880 48390
rect 1104 47898 12880 47920
rect 1104 47846 3315 47898
rect 3367 47846 3379 47898
rect 3431 47846 3443 47898
rect 3495 47846 3507 47898
rect 3559 47846 7982 47898
rect 8034 47846 8046 47898
rect 8098 47846 8110 47898
rect 8162 47846 8174 47898
rect 8226 47846 12880 47898
rect 1104 47824 12880 47846
rect 1104 47354 12880 47376
rect 1104 47302 5648 47354
rect 5700 47302 5712 47354
rect 5764 47302 5776 47354
rect 5828 47302 5840 47354
rect 5892 47302 10315 47354
rect 10367 47302 10379 47354
rect 10431 47302 10443 47354
rect 10495 47302 10507 47354
rect 10559 47302 12880 47354
rect 1104 47280 12880 47302
rect 1104 46810 12880 46832
rect 1104 46758 3315 46810
rect 3367 46758 3379 46810
rect 3431 46758 3443 46810
rect 3495 46758 3507 46810
rect 3559 46758 7982 46810
rect 8034 46758 8046 46810
rect 8098 46758 8110 46810
rect 8162 46758 8174 46810
rect 8226 46758 12880 46810
rect 1104 46736 12880 46758
rect 1104 46266 12880 46288
rect 1104 46214 5648 46266
rect 5700 46214 5712 46266
rect 5764 46214 5776 46266
rect 5828 46214 5840 46266
rect 5892 46214 10315 46266
rect 10367 46214 10379 46266
rect 10431 46214 10443 46266
rect 10495 46214 10507 46266
rect 10559 46214 12880 46266
rect 1104 46192 12880 46214
rect 1104 45722 12880 45744
rect 1104 45670 3315 45722
rect 3367 45670 3379 45722
rect 3431 45670 3443 45722
rect 3495 45670 3507 45722
rect 3559 45670 7982 45722
rect 8034 45670 8046 45722
rect 8098 45670 8110 45722
rect 8162 45670 8174 45722
rect 8226 45670 12880 45722
rect 1104 45648 12880 45670
rect 1104 45178 12880 45200
rect 1104 45126 5648 45178
rect 5700 45126 5712 45178
rect 5764 45126 5776 45178
rect 5828 45126 5840 45178
rect 5892 45126 10315 45178
rect 10367 45126 10379 45178
rect 10431 45126 10443 45178
rect 10495 45126 10507 45178
rect 10559 45126 12880 45178
rect 1104 45104 12880 45126
rect 11698 45064 11704 45076
rect 11659 45036 11704 45064
rect 11698 45024 11704 45036
rect 11756 45024 11762 45076
rect 11514 44928 11520 44940
rect 11475 44900 11520 44928
rect 11514 44888 11520 44900
rect 11572 44888 11578 44940
rect 1104 44634 12880 44656
rect 1104 44582 3315 44634
rect 3367 44582 3379 44634
rect 3431 44582 3443 44634
rect 3495 44582 3507 44634
rect 3559 44582 7982 44634
rect 8034 44582 8046 44634
rect 8098 44582 8110 44634
rect 8162 44582 8174 44634
rect 8226 44582 12880 44634
rect 1104 44560 12880 44582
rect 11514 44520 11520 44532
rect 11475 44492 11520 44520
rect 11514 44480 11520 44492
rect 11572 44480 11578 44532
rect 1104 44090 12880 44112
rect 1104 44038 5648 44090
rect 5700 44038 5712 44090
rect 5764 44038 5776 44090
rect 5828 44038 5840 44090
rect 5892 44038 10315 44090
rect 10367 44038 10379 44090
rect 10431 44038 10443 44090
rect 10495 44038 10507 44090
rect 10559 44038 12880 44090
rect 1104 44016 12880 44038
rect 1104 43546 12880 43568
rect 1104 43494 3315 43546
rect 3367 43494 3379 43546
rect 3431 43494 3443 43546
rect 3495 43494 3507 43546
rect 3559 43494 7982 43546
rect 8034 43494 8046 43546
rect 8098 43494 8110 43546
rect 8162 43494 8174 43546
rect 8226 43494 12880 43546
rect 1104 43472 12880 43494
rect 1104 43002 12880 43024
rect 1104 42950 5648 43002
rect 5700 42950 5712 43002
rect 5764 42950 5776 43002
rect 5828 42950 5840 43002
rect 5892 42950 10315 43002
rect 10367 42950 10379 43002
rect 10431 42950 10443 43002
rect 10495 42950 10507 43002
rect 10559 42950 12880 43002
rect 1104 42928 12880 42950
rect 1104 42458 12880 42480
rect 1104 42406 3315 42458
rect 3367 42406 3379 42458
rect 3431 42406 3443 42458
rect 3495 42406 3507 42458
rect 3559 42406 7982 42458
rect 8034 42406 8046 42458
rect 8098 42406 8110 42458
rect 8162 42406 8174 42458
rect 8226 42406 12880 42458
rect 1104 42384 12880 42406
rect 1104 41914 12880 41936
rect 1104 41862 5648 41914
rect 5700 41862 5712 41914
rect 5764 41862 5776 41914
rect 5828 41862 5840 41914
rect 5892 41862 10315 41914
rect 10367 41862 10379 41914
rect 10431 41862 10443 41914
rect 10495 41862 10507 41914
rect 10559 41862 12880 41914
rect 1104 41840 12880 41862
rect 1104 41370 12880 41392
rect 1104 41318 3315 41370
rect 3367 41318 3379 41370
rect 3431 41318 3443 41370
rect 3495 41318 3507 41370
rect 3559 41318 7982 41370
rect 8034 41318 8046 41370
rect 8098 41318 8110 41370
rect 8162 41318 8174 41370
rect 8226 41318 12880 41370
rect 1104 41296 12880 41318
rect 1104 40826 12880 40848
rect 1104 40774 5648 40826
rect 5700 40774 5712 40826
rect 5764 40774 5776 40826
rect 5828 40774 5840 40826
rect 5892 40774 10315 40826
rect 10367 40774 10379 40826
rect 10431 40774 10443 40826
rect 10495 40774 10507 40826
rect 10559 40774 12880 40826
rect 1104 40752 12880 40774
rect 1104 40282 12880 40304
rect 1104 40230 3315 40282
rect 3367 40230 3379 40282
rect 3431 40230 3443 40282
rect 3495 40230 3507 40282
rect 3559 40230 7982 40282
rect 8034 40230 8046 40282
rect 8098 40230 8110 40282
rect 8162 40230 8174 40282
rect 8226 40230 12880 40282
rect 1104 40208 12880 40230
rect 10778 40168 10784 40180
rect 10739 40140 10784 40168
rect 10778 40128 10784 40140
rect 10836 40168 10842 40180
rect 11514 40168 11520 40180
rect 10836 40140 10916 40168
rect 11475 40140 11520 40168
rect 10836 40128 10842 40140
rect 10888 40041 10916 40140
rect 11514 40128 11520 40140
rect 11572 40128 11578 40180
rect 10873 40035 10931 40041
rect 10873 40001 10885 40035
rect 10919 40001 10931 40035
rect 10873 39995 10931 40001
rect 11057 39967 11115 39973
rect 11057 39933 11069 39967
rect 11103 39964 11115 39967
rect 11238 39964 11244 39976
rect 11103 39936 11244 39964
rect 11103 39933 11115 39936
rect 11057 39927 11115 39933
rect 11238 39924 11244 39936
rect 11296 39924 11302 39976
rect 1104 39738 12880 39760
rect 1104 39686 5648 39738
rect 5700 39686 5712 39738
rect 5764 39686 5776 39738
rect 5828 39686 5840 39738
rect 5892 39686 10315 39738
rect 10367 39686 10379 39738
rect 10431 39686 10443 39738
rect 10495 39686 10507 39738
rect 10559 39686 12880 39738
rect 1104 39664 12880 39686
rect 10965 39287 11023 39293
rect 10965 39253 10977 39287
rect 11011 39284 11023 39287
rect 11238 39284 11244 39296
rect 11011 39256 11244 39284
rect 11011 39253 11023 39256
rect 10965 39247 11023 39253
rect 11238 39244 11244 39256
rect 11296 39244 11302 39296
rect 1104 39194 12880 39216
rect 1104 39142 3315 39194
rect 3367 39142 3379 39194
rect 3431 39142 3443 39194
rect 3495 39142 3507 39194
rect 3559 39142 7982 39194
rect 8034 39142 8046 39194
rect 8098 39142 8110 39194
rect 8162 39142 8174 39194
rect 8226 39142 12880 39194
rect 1104 39120 12880 39142
rect 1104 38650 12880 38672
rect 1104 38598 5648 38650
rect 5700 38598 5712 38650
rect 5764 38598 5776 38650
rect 5828 38598 5840 38650
rect 5892 38598 10315 38650
rect 10367 38598 10379 38650
rect 10431 38598 10443 38650
rect 10495 38598 10507 38650
rect 10559 38598 12880 38650
rect 1104 38576 12880 38598
rect 1104 38106 12880 38128
rect 1104 38054 3315 38106
rect 3367 38054 3379 38106
rect 3431 38054 3443 38106
rect 3495 38054 3507 38106
rect 3559 38054 7982 38106
rect 8034 38054 8046 38106
rect 8098 38054 8110 38106
rect 8162 38054 8174 38106
rect 8226 38054 12880 38106
rect 1104 38032 12880 38054
rect 1104 37562 12880 37584
rect 1104 37510 5648 37562
rect 5700 37510 5712 37562
rect 5764 37510 5776 37562
rect 5828 37510 5840 37562
rect 5892 37510 10315 37562
rect 10367 37510 10379 37562
rect 10431 37510 10443 37562
rect 10495 37510 10507 37562
rect 10559 37510 12880 37562
rect 1104 37488 12880 37510
rect 1104 37018 12880 37040
rect 1104 36966 3315 37018
rect 3367 36966 3379 37018
rect 3431 36966 3443 37018
rect 3495 36966 3507 37018
rect 3559 36966 7982 37018
rect 8034 36966 8046 37018
rect 8098 36966 8110 37018
rect 8162 36966 8174 37018
rect 8226 36966 12880 37018
rect 1104 36944 12880 36966
rect 1104 36474 12880 36496
rect 1104 36422 5648 36474
rect 5700 36422 5712 36474
rect 5764 36422 5776 36474
rect 5828 36422 5840 36474
rect 5892 36422 10315 36474
rect 10367 36422 10379 36474
rect 10431 36422 10443 36474
rect 10495 36422 10507 36474
rect 10559 36422 12880 36474
rect 1104 36400 12880 36422
rect 1104 35930 12880 35952
rect 1104 35878 3315 35930
rect 3367 35878 3379 35930
rect 3431 35878 3443 35930
rect 3495 35878 3507 35930
rect 3559 35878 7982 35930
rect 8034 35878 8046 35930
rect 8098 35878 8110 35930
rect 8162 35878 8174 35930
rect 8226 35878 12880 35930
rect 1104 35856 12880 35878
rect 1104 35386 12880 35408
rect 1104 35334 5648 35386
rect 5700 35334 5712 35386
rect 5764 35334 5776 35386
rect 5828 35334 5840 35386
rect 5892 35334 10315 35386
rect 10367 35334 10379 35386
rect 10431 35334 10443 35386
rect 10495 35334 10507 35386
rect 10559 35334 12880 35386
rect 1104 35312 12880 35334
rect 1104 34842 12880 34864
rect 1104 34790 3315 34842
rect 3367 34790 3379 34842
rect 3431 34790 3443 34842
rect 3495 34790 3507 34842
rect 3559 34790 7982 34842
rect 8034 34790 8046 34842
rect 8098 34790 8110 34842
rect 8162 34790 8174 34842
rect 8226 34790 12880 34842
rect 1104 34768 12880 34790
rect 1104 34298 12880 34320
rect 1104 34246 5648 34298
rect 5700 34246 5712 34298
rect 5764 34246 5776 34298
rect 5828 34246 5840 34298
rect 5892 34246 10315 34298
rect 10367 34246 10379 34298
rect 10431 34246 10443 34298
rect 10495 34246 10507 34298
rect 10559 34246 12880 34298
rect 1104 34224 12880 34246
rect 1104 33754 12880 33776
rect 1104 33702 3315 33754
rect 3367 33702 3379 33754
rect 3431 33702 3443 33754
rect 3495 33702 3507 33754
rect 3559 33702 7982 33754
rect 8034 33702 8046 33754
rect 8098 33702 8110 33754
rect 8162 33702 8174 33754
rect 8226 33702 12880 33754
rect 1104 33680 12880 33702
rect 1104 33210 12880 33232
rect 1104 33158 5648 33210
rect 5700 33158 5712 33210
rect 5764 33158 5776 33210
rect 5828 33158 5840 33210
rect 5892 33158 10315 33210
rect 10367 33158 10379 33210
rect 10431 33158 10443 33210
rect 10495 33158 10507 33210
rect 10559 33158 12880 33210
rect 1104 33136 12880 33158
rect 1104 32666 12880 32688
rect 1104 32614 3315 32666
rect 3367 32614 3379 32666
rect 3431 32614 3443 32666
rect 3495 32614 3507 32666
rect 3559 32614 7982 32666
rect 8034 32614 8046 32666
rect 8098 32614 8110 32666
rect 8162 32614 8174 32666
rect 8226 32614 12880 32666
rect 1104 32592 12880 32614
rect 1104 32122 12880 32144
rect 1104 32070 5648 32122
rect 5700 32070 5712 32122
rect 5764 32070 5776 32122
rect 5828 32070 5840 32122
rect 5892 32070 10315 32122
rect 10367 32070 10379 32122
rect 10431 32070 10443 32122
rect 10495 32070 10507 32122
rect 10559 32070 12880 32122
rect 1104 32048 12880 32070
rect 1104 31578 12880 31600
rect 1104 31526 3315 31578
rect 3367 31526 3379 31578
rect 3431 31526 3443 31578
rect 3495 31526 3507 31578
rect 3559 31526 7982 31578
rect 8034 31526 8046 31578
rect 8098 31526 8110 31578
rect 8162 31526 8174 31578
rect 8226 31526 12880 31578
rect 1104 31504 12880 31526
rect 11422 31464 11428 31476
rect 11383 31436 11428 31464
rect 11422 31424 11428 31436
rect 11480 31424 11486 31476
rect 10962 31288 10968 31340
rect 11020 31328 11026 31340
rect 11020 31300 11284 31328
rect 11020 31288 11026 31300
rect 11256 31269 11284 31300
rect 11241 31263 11299 31269
rect 11241 31229 11253 31263
rect 11287 31260 11299 31263
rect 11793 31263 11851 31269
rect 11793 31260 11805 31263
rect 11287 31232 11805 31260
rect 11287 31229 11299 31232
rect 11241 31223 11299 31229
rect 11793 31229 11805 31232
rect 11839 31229 11851 31263
rect 11793 31223 11851 31229
rect 1104 31034 12880 31056
rect 1104 30982 5648 31034
rect 5700 30982 5712 31034
rect 5764 30982 5776 31034
rect 5828 30982 5840 31034
rect 5892 30982 10315 31034
rect 10367 30982 10379 31034
rect 10431 30982 10443 31034
rect 10495 30982 10507 31034
rect 10559 30982 12880 31034
rect 1104 30960 12880 30982
rect 1104 30490 12880 30512
rect 1104 30438 3315 30490
rect 3367 30438 3379 30490
rect 3431 30438 3443 30490
rect 3495 30438 3507 30490
rect 3559 30438 7982 30490
rect 8034 30438 8046 30490
rect 8098 30438 8110 30490
rect 8162 30438 8174 30490
rect 8226 30438 12880 30490
rect 1104 30416 12880 30438
rect 1104 29946 12880 29968
rect 1104 29894 5648 29946
rect 5700 29894 5712 29946
rect 5764 29894 5776 29946
rect 5828 29894 5840 29946
rect 5892 29894 10315 29946
rect 10367 29894 10379 29946
rect 10431 29894 10443 29946
rect 10495 29894 10507 29946
rect 10559 29894 12880 29946
rect 1104 29872 12880 29894
rect 1104 29402 12880 29424
rect 1104 29350 3315 29402
rect 3367 29350 3379 29402
rect 3431 29350 3443 29402
rect 3495 29350 3507 29402
rect 3559 29350 7982 29402
rect 8034 29350 8046 29402
rect 8098 29350 8110 29402
rect 8162 29350 8174 29402
rect 8226 29350 12880 29402
rect 1104 29328 12880 29350
rect 1104 28858 12880 28880
rect 1104 28806 5648 28858
rect 5700 28806 5712 28858
rect 5764 28806 5776 28858
rect 5828 28806 5840 28858
rect 5892 28806 10315 28858
rect 10367 28806 10379 28858
rect 10431 28806 10443 28858
rect 10495 28806 10507 28858
rect 10559 28806 12880 28858
rect 1104 28784 12880 28806
rect 1104 28314 12880 28336
rect 1104 28262 3315 28314
rect 3367 28262 3379 28314
rect 3431 28262 3443 28314
rect 3495 28262 3507 28314
rect 3559 28262 7982 28314
rect 8034 28262 8046 28314
rect 8098 28262 8110 28314
rect 8162 28262 8174 28314
rect 8226 28262 12880 28314
rect 1104 28240 12880 28262
rect 1104 27770 12880 27792
rect 1104 27718 5648 27770
rect 5700 27718 5712 27770
rect 5764 27718 5776 27770
rect 5828 27718 5840 27770
rect 5892 27718 10315 27770
rect 10367 27718 10379 27770
rect 10431 27718 10443 27770
rect 10495 27718 10507 27770
rect 10559 27718 12880 27770
rect 1104 27696 12880 27718
rect 1104 27226 12880 27248
rect 1104 27174 3315 27226
rect 3367 27174 3379 27226
rect 3431 27174 3443 27226
rect 3495 27174 3507 27226
rect 3559 27174 7982 27226
rect 8034 27174 8046 27226
rect 8098 27174 8110 27226
rect 8162 27174 8174 27226
rect 8226 27174 12880 27226
rect 1104 27152 12880 27174
rect 10778 27112 10784 27124
rect 10739 27084 10784 27112
rect 10778 27072 10784 27084
rect 10836 27112 10842 27124
rect 10836 27084 10916 27112
rect 10836 27072 10842 27084
rect 10888 26985 10916 27084
rect 10962 27072 10968 27124
rect 11020 27112 11026 27124
rect 11241 27115 11299 27121
rect 11241 27112 11253 27115
rect 11020 27084 11253 27112
rect 11020 27072 11026 27084
rect 11241 27081 11253 27084
rect 11287 27081 11299 27115
rect 11241 27075 11299 27081
rect 10873 26979 10931 26985
rect 10873 26945 10885 26979
rect 10919 26945 10931 26979
rect 10873 26939 10931 26945
rect 10962 26868 10968 26920
rect 11020 26908 11026 26920
rect 11057 26911 11115 26917
rect 11057 26908 11069 26911
rect 11020 26880 11069 26908
rect 11020 26868 11026 26880
rect 11057 26877 11069 26880
rect 11103 26877 11115 26911
rect 11057 26871 11115 26877
rect 1104 26682 12880 26704
rect 1104 26630 5648 26682
rect 5700 26630 5712 26682
rect 5764 26630 5776 26682
rect 5828 26630 5840 26682
rect 5892 26630 10315 26682
rect 10367 26630 10379 26682
rect 10431 26630 10443 26682
rect 10495 26630 10507 26682
rect 10559 26630 12880 26682
rect 1104 26608 12880 26630
rect 9398 26188 9404 26240
rect 9456 26228 9462 26240
rect 10873 26231 10931 26237
rect 10873 26228 10885 26231
rect 9456 26200 10885 26228
rect 9456 26188 9462 26200
rect 10873 26197 10885 26200
rect 10919 26228 10931 26231
rect 10962 26228 10968 26240
rect 10919 26200 10968 26228
rect 10919 26197 10931 26200
rect 10873 26191 10931 26197
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 1104 26138 12880 26160
rect 1104 26086 3315 26138
rect 3367 26086 3379 26138
rect 3431 26086 3443 26138
rect 3495 26086 3507 26138
rect 3559 26086 7982 26138
rect 8034 26086 8046 26138
rect 8098 26086 8110 26138
rect 8162 26086 8174 26138
rect 8226 26086 12880 26138
rect 1104 26064 12880 26086
rect 1104 25594 12880 25616
rect 1104 25542 5648 25594
rect 5700 25542 5712 25594
rect 5764 25542 5776 25594
rect 5828 25542 5840 25594
rect 5892 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 12880 25594
rect 1104 25520 12880 25542
rect 1104 25050 12880 25072
rect 1104 24998 3315 25050
rect 3367 24998 3379 25050
rect 3431 24998 3443 25050
rect 3495 24998 3507 25050
rect 3559 24998 7982 25050
rect 8034 24998 8046 25050
rect 8098 24998 8110 25050
rect 8162 24998 8174 25050
rect 8226 24998 12880 25050
rect 1104 24976 12880 24998
rect 1104 24506 12880 24528
rect 1104 24454 5648 24506
rect 5700 24454 5712 24506
rect 5764 24454 5776 24506
rect 5828 24454 5840 24506
rect 5892 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 12880 24506
rect 1104 24432 12880 24454
rect 1104 23962 12880 23984
rect 1104 23910 3315 23962
rect 3367 23910 3379 23962
rect 3431 23910 3443 23962
rect 3495 23910 3507 23962
rect 3559 23910 7982 23962
rect 8034 23910 8046 23962
rect 8098 23910 8110 23962
rect 8162 23910 8174 23962
rect 8226 23910 12880 23962
rect 1104 23888 12880 23910
rect 1104 23418 12880 23440
rect 1104 23366 5648 23418
rect 5700 23366 5712 23418
rect 5764 23366 5776 23418
rect 5828 23366 5840 23418
rect 5892 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 12880 23418
rect 1104 23344 12880 23366
rect 1104 22874 12880 22896
rect 1104 22822 3315 22874
rect 3367 22822 3379 22874
rect 3431 22822 3443 22874
rect 3495 22822 3507 22874
rect 3559 22822 7982 22874
rect 8034 22822 8046 22874
rect 8098 22822 8110 22874
rect 8162 22822 8174 22874
rect 8226 22822 12880 22874
rect 1104 22800 12880 22822
rect 1104 22330 12880 22352
rect 1104 22278 5648 22330
rect 5700 22278 5712 22330
rect 5764 22278 5776 22330
rect 5828 22278 5840 22330
rect 5892 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 12880 22330
rect 1104 22256 12880 22278
rect 1104 21786 12880 21808
rect 1104 21734 3315 21786
rect 3367 21734 3379 21786
rect 3431 21734 3443 21786
rect 3495 21734 3507 21786
rect 3559 21734 7982 21786
rect 8034 21734 8046 21786
rect 8098 21734 8110 21786
rect 8162 21734 8174 21786
rect 8226 21734 12880 21786
rect 1104 21712 12880 21734
rect 1104 21242 12880 21264
rect 1104 21190 5648 21242
rect 5700 21190 5712 21242
rect 5764 21190 5776 21242
rect 5828 21190 5840 21242
rect 5892 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 12880 21242
rect 1104 21168 12880 21190
rect 1104 20698 12880 20720
rect 1104 20646 3315 20698
rect 3367 20646 3379 20698
rect 3431 20646 3443 20698
rect 3495 20646 3507 20698
rect 3559 20646 7982 20698
rect 8034 20646 8046 20698
rect 8098 20646 8110 20698
rect 8162 20646 8174 20698
rect 8226 20646 12880 20698
rect 1104 20624 12880 20646
rect 1104 20154 12880 20176
rect 1104 20102 5648 20154
rect 5700 20102 5712 20154
rect 5764 20102 5776 20154
rect 5828 20102 5840 20154
rect 5892 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 12880 20154
rect 1104 20080 12880 20102
rect 1104 19610 12880 19632
rect 1104 19558 3315 19610
rect 3367 19558 3379 19610
rect 3431 19558 3443 19610
rect 3495 19558 3507 19610
rect 3559 19558 7982 19610
rect 8034 19558 8046 19610
rect 8098 19558 8110 19610
rect 8162 19558 8174 19610
rect 8226 19558 12880 19610
rect 1104 19536 12880 19558
rect 11238 19496 11244 19508
rect 11199 19468 11244 19496
rect 11238 19456 11244 19468
rect 11296 19456 11302 19508
rect 10042 19252 10048 19304
rect 10100 19292 10106 19304
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 10100 19264 10333 19292
rect 10100 19252 10106 19264
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10321 19255 10379 19261
rect 10683 19227 10741 19233
rect 10683 19193 10695 19227
rect 10729 19193 10741 19227
rect 10683 19187 10741 19193
rect 10229 19159 10287 19165
rect 10229 19125 10241 19159
rect 10275 19156 10287 19159
rect 10698 19156 10726 19187
rect 10778 19156 10784 19168
rect 10275 19128 10784 19156
rect 10275 19125 10287 19128
rect 10229 19119 10287 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 1104 19066 12880 19088
rect 1104 19014 5648 19066
rect 5700 19014 5712 19066
rect 5764 19014 5776 19066
rect 5828 19014 5840 19066
rect 5892 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 12880 19066
rect 1104 18992 12880 19014
rect 11606 18952 11612 18964
rect 11567 18924 11612 18952
rect 11606 18912 11612 18924
rect 11664 18912 11670 18964
rect 10778 18844 10784 18896
rect 10836 18884 10842 18896
rect 11010 18887 11068 18893
rect 11010 18884 11022 18887
rect 10836 18856 11022 18884
rect 10836 18844 10842 18856
rect 11010 18853 11022 18856
rect 11056 18853 11068 18887
rect 11010 18847 11068 18853
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 10689 18751 10747 18757
rect 10689 18748 10701 18751
rect 8812 18720 10701 18748
rect 8812 18708 8818 18720
rect 10689 18717 10701 18720
rect 10735 18748 10747 18751
rect 11790 18748 11796 18760
rect 10735 18720 11796 18748
rect 10735 18717 10747 18720
rect 10689 18711 10747 18717
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 8570 18612 8576 18624
rect 8531 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 10042 18572 10048 18624
rect 10100 18612 10106 18624
rect 10321 18615 10379 18621
rect 10321 18612 10333 18615
rect 10100 18584 10333 18612
rect 10100 18572 10106 18584
rect 10321 18581 10333 18584
rect 10367 18581 10379 18615
rect 10321 18575 10379 18581
rect 1104 18522 12880 18544
rect 1104 18470 3315 18522
rect 3367 18470 3379 18522
rect 3431 18470 3443 18522
rect 3495 18470 3507 18522
rect 3559 18470 7982 18522
rect 8034 18470 8046 18522
rect 8098 18470 8110 18522
rect 8162 18470 8174 18522
rect 8226 18470 12880 18522
rect 1104 18448 12880 18470
rect 9398 18408 9404 18420
rect 9359 18380 9404 18408
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 11146 18408 11152 18420
rect 11107 18380 11152 18408
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 11790 18408 11796 18420
rect 11751 18380 11796 18408
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 8858 18244 9873 18272
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18204 8539 18207
rect 8570 18204 8576 18216
rect 8527 18176 8576 18204
rect 8527 18173 8539 18176
rect 8481 18167 8539 18173
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 8858 18145 8886 18244
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 9692 18176 10241 18204
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18136 8447 18139
rect 8843 18139 8901 18145
rect 8843 18136 8855 18139
rect 8435 18108 8855 18136
rect 8435 18105 8447 18108
rect 8389 18099 8447 18105
rect 8843 18105 8855 18108
rect 8889 18105 8901 18139
rect 8843 18099 8901 18105
rect 9692 18080 9720 18176
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 10550 18139 10608 18145
rect 10550 18105 10562 18139
rect 10596 18105 10608 18139
rect 10550 18099 10608 18105
rect 9674 18068 9680 18080
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18068 9919 18071
rect 10137 18071 10195 18077
rect 10137 18068 10149 18071
rect 9907 18040 10149 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 10137 18037 10149 18040
rect 10183 18068 10195 18071
rect 10565 18068 10593 18099
rect 10778 18068 10784 18080
rect 10183 18040 10784 18068
rect 10183 18037 10195 18040
rect 10137 18031 10195 18037
rect 10778 18028 10784 18040
rect 10836 18068 10842 18080
rect 11425 18071 11483 18077
rect 11425 18068 11437 18071
rect 10836 18040 11437 18068
rect 10836 18028 10842 18040
rect 11425 18037 11437 18040
rect 11471 18037 11483 18071
rect 11425 18031 11483 18037
rect 1104 17978 12880 18000
rect 1104 17926 5648 17978
rect 5700 17926 5712 17978
rect 5764 17926 5776 17978
rect 5828 17926 5840 17978
rect 5892 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 12880 17978
rect 1104 17904 12880 17926
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 10499 17799 10557 17805
rect 10499 17765 10511 17799
rect 10545 17796 10557 17799
rect 10778 17796 10784 17808
rect 10545 17768 10784 17796
rect 10545 17765 10557 17768
rect 10499 17759 10557 17765
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 8662 17524 8668 17536
rect 8623 17496 8668 17524
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 1104 17434 12880 17456
rect 1104 17382 3315 17434
rect 3367 17382 3379 17434
rect 3431 17382 3443 17434
rect 3495 17382 3507 17434
rect 3559 17382 7982 17434
rect 8034 17382 8046 17434
rect 8098 17382 8110 17434
rect 8162 17382 8174 17434
rect 8226 17382 12880 17434
rect 1104 17360 12880 17382
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 10781 17323 10839 17329
rect 10781 17320 10793 17323
rect 10192 17292 10793 17320
rect 10192 17280 10198 17292
rect 10781 17289 10793 17292
rect 10827 17289 10839 17323
rect 10781 17283 10839 17289
rect 10686 17212 10692 17264
rect 10744 17252 10750 17264
rect 11425 17255 11483 17261
rect 11425 17252 11437 17255
rect 10744 17224 11437 17252
rect 10744 17212 10750 17224
rect 11425 17221 11437 17224
rect 11471 17221 11483 17255
rect 11425 17215 11483 17221
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 8665 17119 8723 17125
rect 8665 17116 8677 17119
rect 8536 17088 8677 17116
rect 8536 17076 8542 17088
rect 8665 17085 8677 17088
rect 8711 17085 8723 17119
rect 8665 17079 8723 17085
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17085 9183 17119
rect 9125 17079 9183 17085
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 9766 17116 9772 17128
rect 9723 17088 9772 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9140 17048 9168 17079
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 11238 17116 11244 17128
rect 9916 17088 9961 17116
rect 11199 17088 11244 17116
rect 9916 17076 9922 17088
rect 11238 17076 11244 17088
rect 11296 17116 11302 17128
rect 11790 17116 11796 17128
rect 11296 17088 11796 17116
rect 11296 17076 11302 17088
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 8312 17020 9168 17048
rect 8312 16992 8340 17020
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 8294 16980 8300 16992
rect 8251 16952 8300 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 8478 16980 8484 16992
rect 8439 16952 8484 16980
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 8570 16940 8576 16992
rect 8628 16980 8634 16992
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8628 16952 8769 16980
rect 8628 16940 8634 16952
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 8757 16943 8815 16949
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 10778 16980 10784 16992
rect 10551 16952 10784 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 1104 16890 12880 16912
rect 1104 16838 5648 16890
rect 5700 16838 5712 16890
rect 5764 16838 5776 16890
rect 5828 16838 5840 16890
rect 5892 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 12880 16890
rect 1104 16816 12880 16838
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 11609 16779 11667 16785
rect 11609 16776 11621 16779
rect 10008 16748 11621 16776
rect 10008 16736 10014 16748
rect 11609 16745 11621 16748
rect 11655 16745 11667 16779
rect 11609 16739 11667 16745
rect 10778 16668 10784 16720
rect 10836 16708 10842 16720
rect 11010 16711 11068 16717
rect 11010 16708 11022 16711
rect 10836 16680 11022 16708
rect 10836 16668 10842 16680
rect 11010 16677 11022 16680
rect 11056 16677 11068 16711
rect 11010 16671 11068 16677
rect 10686 16572 10692 16584
rect 10647 16544 10692 16572
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 8570 16464 8576 16516
rect 8628 16504 8634 16516
rect 9033 16507 9091 16513
rect 9033 16504 9045 16507
rect 8628 16476 9045 16504
rect 8628 16464 8634 16476
rect 9033 16473 9045 16476
rect 9079 16504 9091 16507
rect 9950 16504 9956 16516
rect 9079 16476 9956 16504
rect 9079 16473 9091 16476
rect 9033 16467 9091 16473
rect 9950 16464 9956 16476
rect 10008 16464 10014 16516
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16436 8815 16439
rect 8938 16436 8944 16448
rect 8803 16408 8944 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 8938 16396 8944 16408
rect 8996 16396 9002 16448
rect 1104 16346 12880 16368
rect 1104 16294 3315 16346
rect 3367 16294 3379 16346
rect 3431 16294 3443 16346
rect 3495 16294 3507 16346
rect 3559 16294 7982 16346
rect 8034 16294 8046 16346
rect 8098 16294 8110 16346
rect 8162 16294 8174 16346
rect 8226 16294 12880 16346
rect 1104 16272 12880 16294
rect 10686 16192 10692 16244
rect 10744 16232 10750 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10744 16204 11069 16232
rect 10744 16192 10750 16204
rect 11057 16201 11069 16204
rect 11103 16232 11115 16235
rect 11238 16232 11244 16244
rect 11103 16204 11244 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 10042 16124 10048 16176
rect 10100 16164 10106 16176
rect 10229 16167 10287 16173
rect 10229 16164 10241 16167
rect 10100 16136 10241 16164
rect 10100 16124 10106 16136
rect 10229 16133 10241 16136
rect 10275 16133 10287 16167
rect 10229 16127 10287 16133
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16096 8079 16099
rect 8294 16096 8300 16108
rect 8067 16068 8300 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 8294 16056 8300 16068
rect 8352 16096 8358 16108
rect 8352 16068 9076 16096
rect 8352 16056 8358 16068
rect 9048 16040 9076 16068
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 15997 8907 16031
rect 8849 15991 8907 15997
rect 7834 15920 7840 15972
rect 7892 15960 7898 15972
rect 8297 15963 8355 15969
rect 8297 15960 8309 15963
rect 7892 15932 8309 15960
rect 7892 15920 7898 15932
rect 8297 15929 8309 15932
rect 8343 15960 8355 15963
rect 8864 15960 8892 15991
rect 9030 15988 9036 16040
rect 9088 16028 9094 16040
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 9088 16000 9321 16028
rect 9088 15988 9094 16000
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9766 16028 9772 16040
rect 9727 16000 9772 16028
rect 9309 15991 9367 15997
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 9950 15988 9956 16040
rect 10008 16028 10014 16040
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 10008 16000 10057 16028
rect 10008 15988 10014 16000
rect 10045 15997 10057 16000
rect 10091 15997 10103 16031
rect 10045 15991 10103 15997
rect 8343 15932 8892 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 8757 15895 8815 15901
rect 8757 15861 8769 15895
rect 8803 15892 8815 15895
rect 8938 15892 8944 15904
rect 8803 15864 8944 15892
rect 8803 15861 8815 15864
rect 8757 15855 8815 15861
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 10686 15892 10692 15904
rect 10647 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 1104 15802 12880 15824
rect 1104 15750 5648 15802
rect 5700 15750 5712 15802
rect 5764 15750 5776 15802
rect 5828 15750 5840 15802
rect 5892 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 12880 15802
rect 1104 15728 12880 15750
rect 8205 15691 8263 15697
rect 8205 15657 8217 15691
rect 8251 15688 8263 15691
rect 9950 15688 9956 15700
rect 8251 15660 9536 15688
rect 9911 15660 9956 15688
rect 8251 15657 8263 15660
rect 8205 15651 8263 15657
rect 7374 15580 7380 15632
rect 7432 15620 7438 15632
rect 8389 15623 8447 15629
rect 8389 15620 8401 15623
rect 7432 15592 8401 15620
rect 7432 15580 7438 15592
rect 8389 15589 8401 15592
rect 8435 15620 8447 15623
rect 8570 15620 8576 15632
rect 8435 15592 8576 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 8754 15620 8760 15632
rect 8715 15592 8760 15620
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9508 15629 9536 15660
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 9493 15623 9551 15629
rect 9493 15589 9505 15623
rect 9539 15620 9551 15623
rect 9539 15592 9674 15620
rect 9539 15589 9551 15592
rect 9493 15583 9551 15589
rect 8294 15552 8300 15564
rect 8255 15524 8300 15552
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 9646 15552 9674 15592
rect 9858 15580 9864 15632
rect 9916 15620 9922 15632
rect 10045 15623 10103 15629
rect 9916 15592 9961 15620
rect 9916 15580 9922 15592
rect 10045 15589 10057 15623
rect 10091 15589 10103 15623
rect 10045 15583 10103 15589
rect 10060 15552 10088 15583
rect 10134 15580 10140 15632
rect 10192 15620 10198 15632
rect 10413 15623 10471 15629
rect 10413 15620 10425 15623
rect 10192 15592 10425 15620
rect 10192 15580 10198 15592
rect 10413 15589 10425 15592
rect 10459 15589 10471 15623
rect 10413 15583 10471 15589
rect 10686 15552 10692 15564
rect 9646 15524 9904 15552
rect 7834 15444 7840 15496
rect 7892 15484 7898 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7892 15456 8033 15484
rect 7892 15444 7898 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15484 9735 15487
rect 9766 15484 9772 15496
rect 9723 15456 9772 15484
rect 9723 15453 9735 15456
rect 9677 15447 9735 15453
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8996 15320 9045 15348
rect 8996 15308 9002 15320
rect 9033 15317 9045 15320
rect 9079 15348 9091 15351
rect 9692 15348 9720 15447
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 9876 15484 9904 15524
rect 10060 15524 10692 15552
rect 10060 15484 10088 15524
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 9876 15456 10088 15484
rect 10686 15348 10692 15360
rect 9079 15320 9720 15348
rect 10647 15320 10692 15348
rect 9079 15317 9091 15320
rect 9033 15311 9091 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 1104 15258 12880 15280
rect 1104 15206 3315 15258
rect 3367 15206 3379 15258
rect 3431 15206 3443 15258
rect 3495 15206 3507 15258
rect 3559 15206 7982 15258
rect 8034 15206 8046 15258
rect 8098 15206 8110 15258
rect 8162 15206 8174 15258
rect 8226 15206 12880 15258
rect 1104 15184 12880 15206
rect 7374 15144 7380 15156
rect 7335 15116 7380 15144
rect 7374 15104 7380 15116
rect 7432 15104 7438 15156
rect 8113 15147 8171 15153
rect 8113 15113 8125 15147
rect 8159 15144 8171 15147
rect 8294 15144 8300 15156
rect 8159 15116 8300 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8294 15104 8300 15116
rect 8352 15144 8358 15156
rect 9214 15144 9220 15156
rect 8352 15116 9220 15144
rect 8352 15104 8358 15116
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 9950 15144 9956 15156
rect 9911 15116 9956 15144
rect 9950 15104 9956 15116
rect 10008 15144 10014 15156
rect 10321 15147 10379 15153
rect 10321 15144 10333 15147
rect 10008 15116 10333 15144
rect 10008 15104 10014 15116
rect 10321 15113 10333 15116
rect 10367 15144 10379 15147
rect 10367 15116 10548 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 8481 15011 8539 15017
rect 8481 14977 8493 15011
rect 8527 15008 8539 15011
rect 9306 15008 9312 15020
rect 8527 14980 9312 15008
rect 8527 14977 8539 14980
rect 8481 14971 8539 14977
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 9674 15008 9680 15020
rect 9635 14980 9680 15008
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 10520 15017 10548 15116
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 14977 10563 15011
rect 11238 15008 11244 15020
rect 11199 14980 11244 15008
rect 10505 14971 10563 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8895 14912 9137 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 9125 14909 9137 14912
rect 9171 14940 9183 14943
rect 9766 14940 9772 14952
rect 9171 14912 9772 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 7745 14875 7803 14881
rect 7745 14841 7757 14875
rect 7791 14872 7803 14875
rect 7834 14872 7840 14884
rect 7791 14844 7840 14872
rect 7791 14841 7803 14844
rect 7745 14835 7803 14841
rect 7834 14832 7840 14844
rect 7892 14872 7898 14884
rect 8938 14872 8944 14884
rect 7892 14844 8800 14872
rect 8899 14844 8944 14872
rect 7892 14832 7898 14844
rect 8772 14816 8800 14844
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 9306 14872 9312 14884
rect 9219 14844 9312 14872
rect 9306 14832 9312 14844
rect 9364 14872 9370 14884
rect 9582 14872 9588 14884
rect 9364 14844 9588 14872
rect 9364 14832 9370 14844
rect 9582 14832 9588 14844
rect 9640 14872 9646 14884
rect 10704 14872 10732 14900
rect 10870 14872 10876 14884
rect 9640 14844 10732 14872
rect 10831 14844 10876 14872
rect 9640 14832 9646 14844
rect 10870 14832 10876 14844
rect 10928 14872 10934 14884
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 10928 14844 11529 14872
rect 10928 14832 10934 14844
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 9217 14807 9275 14813
rect 9217 14804 9229 14807
rect 8812 14776 9229 14804
rect 8812 14764 8818 14776
rect 9217 14773 9229 14776
rect 9263 14773 9275 14807
rect 9217 14767 9275 14773
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 9950 14804 9956 14816
rect 9456 14776 9956 14804
rect 9456 14764 9462 14776
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 1104 14714 12880 14736
rect 1104 14662 5648 14714
rect 5700 14662 5712 14714
rect 5764 14662 5776 14714
rect 5828 14662 5840 14714
rect 5892 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 12880 14714
rect 1104 14640 12880 14662
rect 9125 14603 9183 14609
rect 9125 14569 9137 14603
rect 9171 14600 9183 14603
rect 9306 14600 9312 14612
rect 9171 14572 9312 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9214 14492 9220 14544
rect 9272 14532 9278 14544
rect 10689 14535 10747 14541
rect 10689 14532 10701 14535
rect 9272 14504 10701 14532
rect 9272 14492 9278 14504
rect 10689 14501 10701 14504
rect 10735 14532 10747 14535
rect 10778 14532 10784 14544
rect 10735 14504 10784 14532
rect 10735 14501 10747 14504
rect 10689 14495 10747 14501
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 8113 14467 8171 14473
rect 8113 14464 8125 14467
rect 7892 14436 8125 14464
rect 7892 14424 7898 14436
rect 8113 14433 8125 14436
rect 8159 14464 8171 14467
rect 8478 14464 8484 14476
rect 8159 14436 8484 14464
rect 8159 14433 8171 14436
rect 8113 14427 8171 14433
rect 8478 14424 8484 14436
rect 8536 14464 8542 14476
rect 9306 14464 9312 14476
rect 8536 14436 9312 14464
rect 8536 14424 8542 14436
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 9403 14436 9505 14464
rect 9493 14433 9505 14436
rect 9539 14464 9551 14467
rect 9766 14464 9772 14476
rect 9539 14436 9772 14464
rect 9539 14433 9551 14436
rect 9493 14427 9551 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 8754 14396 8760 14408
rect 8715 14368 8760 14396
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 10870 14396 10876 14408
rect 9723 14368 10876 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 8570 14288 8576 14340
rect 8628 14328 8634 14340
rect 9692 14328 9720 14359
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 8628 14300 9720 14328
rect 8628 14288 8634 14300
rect 1104 14170 12880 14192
rect 1104 14118 3315 14170
rect 3367 14118 3379 14170
rect 3431 14118 3443 14170
rect 3495 14118 3507 14170
rect 3559 14118 7982 14170
rect 8034 14118 8046 14170
rect 8098 14118 8110 14170
rect 8162 14118 8174 14170
rect 8226 14118 12880 14170
rect 1104 14096 12880 14118
rect 8938 13812 8944 13864
rect 8996 13852 9002 13864
rect 9398 13852 9404 13864
rect 8996 13824 9404 13852
rect 8996 13812 9002 13824
rect 9398 13812 9404 13824
rect 9456 13852 9462 13864
rect 10042 13852 10048 13864
rect 9456 13824 10048 13852
rect 9456 13812 9462 13824
rect 10042 13812 10048 13824
rect 10100 13812 10106 13864
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 8021 13719 8079 13725
rect 8021 13716 8033 13719
rect 7892 13688 8033 13716
rect 7892 13676 7898 13688
rect 8021 13685 8033 13688
rect 8067 13685 8079 13719
rect 8021 13679 8079 13685
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8812 13688 8953 13716
rect 8812 13676 8818 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 9766 13716 9772 13728
rect 9727 13688 9772 13716
rect 8941 13679 8999 13685
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 10042 13716 10048 13728
rect 10003 13688 10048 13716
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 1104 13626 12880 13648
rect 1104 13574 5648 13626
rect 5700 13574 5712 13626
rect 5764 13574 5776 13626
rect 5828 13574 5840 13626
rect 5892 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 12880 13626
rect 1104 13552 12880 13574
rect 11790 13512 11796 13524
rect 11751 13484 11796 13512
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 11146 13376 11152 13388
rect 11107 13348 11152 13376
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11296 13280 11345 13308
rect 11296 13268 11302 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 1104 13082 12880 13104
rect 1104 13030 3315 13082
rect 3367 13030 3379 13082
rect 3431 13030 3443 13082
rect 3495 13030 3507 13082
rect 3559 13030 7982 13082
rect 8034 13030 8046 13082
rect 8098 13030 8110 13082
rect 8162 13030 8174 13082
rect 8226 13030 12880 13082
rect 1104 13008 12880 13030
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 8205 12767 8263 12773
rect 8205 12733 8217 12767
rect 8251 12764 8263 12767
rect 9582 12764 9588 12776
rect 8251 12736 9588 12764
rect 8251 12733 8263 12736
rect 8205 12727 8263 12733
rect 1302 12588 1308 12640
rect 1360 12628 1366 12640
rect 7929 12631 7987 12637
rect 7929 12628 7941 12631
rect 1360 12600 7941 12628
rect 1360 12588 1366 12600
rect 7929 12597 7941 12600
rect 7975 12628 7987 12631
rect 8220 12628 8248 12727
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 8849 12699 8907 12705
rect 8849 12665 8861 12699
rect 8895 12696 8907 12699
rect 9030 12696 9036 12708
rect 8895 12668 9036 12696
rect 8895 12665 8907 12668
rect 8849 12659 8907 12665
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 7975 12600 8248 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11296 12600 11529 12628
rect 11296 12588 11302 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 11517 12591 11575 12597
rect 1104 12538 12880 12560
rect 1104 12486 5648 12538
rect 5700 12486 5712 12538
rect 5764 12486 5776 12538
rect 5828 12486 5840 12538
rect 5892 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 12880 12538
rect 1104 12464 12880 12486
rect 8754 12084 8760 12096
rect 8715 12056 8760 12084
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 1104 11994 12880 12016
rect 1104 11942 3315 11994
rect 3367 11942 3379 11994
rect 3431 11942 3443 11994
rect 3495 11942 3507 11994
rect 3559 11942 7982 11994
rect 8034 11942 8046 11994
rect 8098 11942 8110 11994
rect 8162 11942 8174 11994
rect 8226 11942 12880 11994
rect 1104 11920 12880 11942
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 9766 11744 9772 11756
rect 8711 11716 9772 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 9766 11704 9772 11716
rect 9824 11744 9830 11756
rect 9824 11716 9996 11744
rect 9824 11704 9830 11716
rect 8754 11676 8760 11688
rect 8715 11648 8760 11676
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9217 11679 9275 11685
rect 9217 11676 9229 11679
rect 9088 11648 9229 11676
rect 9088 11636 9094 11648
rect 9217 11645 9229 11648
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 9968 11685 9996 11716
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9456 11648 9597 11676
rect 9456 11636 9462 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11645 10011 11679
rect 9953 11639 10011 11645
rect 8297 11611 8355 11617
rect 8297 11577 8309 11611
rect 8343 11608 8355 11611
rect 9048 11608 9076 11636
rect 8343 11580 9076 11608
rect 8343 11577 8355 11580
rect 8297 11571 8355 11577
rect 10134 11540 10140 11552
rect 10095 11512 10140 11540
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 1104 11450 12880 11472
rect 1104 11398 5648 11450
rect 5700 11398 5712 11450
rect 5764 11398 5776 11450
rect 5828 11398 5840 11450
rect 5892 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 12880 11450
rect 1104 11376 12880 11398
rect 10686 11336 10692 11348
rect 10647 11308 10692 11336
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10192 11172 10333 11200
rect 10192 11160 10198 11172
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 8849 10999 8907 11005
rect 8849 10965 8861 10999
rect 8895 10996 8907 10999
rect 9398 10996 9404 11008
rect 8895 10968 9404 10996
rect 8895 10965 8907 10968
rect 8849 10959 8907 10965
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 1104 10906 12880 10928
rect 1104 10854 3315 10906
rect 3367 10854 3379 10906
rect 3431 10854 3443 10906
rect 3495 10854 3507 10906
rect 3559 10854 7982 10906
rect 8034 10854 8046 10906
rect 8098 10854 8110 10906
rect 8162 10854 8174 10906
rect 8226 10854 12880 10906
rect 1104 10832 12880 10854
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10689 10795 10747 10801
rect 10689 10792 10701 10795
rect 10192 10764 10701 10792
rect 10192 10752 10198 10764
rect 10689 10761 10701 10764
rect 10735 10761 10747 10795
rect 10689 10755 10747 10761
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9548 10424 10333 10452
rect 9548 10412 9554 10424
rect 10321 10421 10333 10424
rect 10367 10452 10379 10455
rect 10686 10452 10692 10464
rect 10367 10424 10692 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 1104 10362 12880 10384
rect 1104 10310 5648 10362
rect 5700 10310 5712 10362
rect 5764 10310 5776 10362
rect 5828 10310 5840 10362
rect 5892 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 12880 10362
rect 1104 10288 12880 10310
rect 1104 9818 12880 9840
rect 1104 9766 3315 9818
rect 3367 9766 3379 9818
rect 3431 9766 3443 9818
rect 3495 9766 3507 9818
rect 3559 9766 7982 9818
rect 8034 9766 8046 9818
rect 8098 9766 8110 9818
rect 8162 9766 8174 9818
rect 8226 9766 12880 9818
rect 1104 9744 12880 9766
rect 1104 9274 12880 9296
rect 1104 9222 5648 9274
rect 5700 9222 5712 9274
rect 5764 9222 5776 9274
rect 5828 9222 5840 9274
rect 5892 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 12880 9274
rect 1104 9200 12880 9222
rect 1104 8730 12880 8752
rect 1104 8678 3315 8730
rect 3367 8678 3379 8730
rect 3431 8678 3443 8730
rect 3495 8678 3507 8730
rect 3559 8678 7982 8730
rect 8034 8678 8046 8730
rect 8098 8678 8110 8730
rect 8162 8678 8174 8730
rect 8226 8678 12880 8730
rect 1104 8656 12880 8678
rect 1104 8186 12880 8208
rect 1104 8134 5648 8186
rect 5700 8134 5712 8186
rect 5764 8134 5776 8186
rect 5828 8134 5840 8186
rect 5892 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 12880 8186
rect 1104 8112 12880 8134
rect 1104 7642 12880 7664
rect 1104 7590 3315 7642
rect 3367 7590 3379 7642
rect 3431 7590 3443 7642
rect 3495 7590 3507 7642
rect 3559 7590 7982 7642
rect 8034 7590 8046 7642
rect 8098 7590 8110 7642
rect 8162 7590 8174 7642
rect 8226 7590 12880 7642
rect 1104 7568 12880 7590
rect 1104 7098 12880 7120
rect 1104 7046 5648 7098
rect 5700 7046 5712 7098
rect 5764 7046 5776 7098
rect 5828 7046 5840 7098
rect 5892 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 12880 7098
rect 1104 7024 12880 7046
rect 1104 6554 12880 6576
rect 1104 6502 3315 6554
rect 3367 6502 3379 6554
rect 3431 6502 3443 6554
rect 3495 6502 3507 6554
rect 3559 6502 7982 6554
rect 8034 6502 8046 6554
rect 8098 6502 8110 6554
rect 8162 6502 8174 6554
rect 8226 6502 12880 6554
rect 1104 6480 12880 6502
rect 1104 6010 12880 6032
rect 1104 5958 5648 6010
rect 5700 5958 5712 6010
rect 5764 5958 5776 6010
rect 5828 5958 5840 6010
rect 5892 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 12880 6010
rect 1104 5936 12880 5958
rect 1104 5466 12880 5488
rect 1104 5414 3315 5466
rect 3367 5414 3379 5466
rect 3431 5414 3443 5466
rect 3495 5414 3507 5466
rect 3559 5414 7982 5466
rect 8034 5414 8046 5466
rect 8098 5414 8110 5466
rect 8162 5414 8174 5466
rect 8226 5414 12880 5466
rect 1104 5392 12880 5414
rect 1104 4922 12880 4944
rect 1104 4870 5648 4922
rect 5700 4870 5712 4922
rect 5764 4870 5776 4922
rect 5828 4870 5840 4922
rect 5892 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 12880 4922
rect 1104 4848 12880 4870
rect 1104 4378 12880 4400
rect 1104 4326 3315 4378
rect 3367 4326 3379 4378
rect 3431 4326 3443 4378
rect 3495 4326 3507 4378
rect 3559 4326 7982 4378
rect 8034 4326 8046 4378
rect 8098 4326 8110 4378
rect 8162 4326 8174 4378
rect 8226 4326 12880 4378
rect 1104 4304 12880 4326
rect 11422 4264 11428 4276
rect 11383 4236 11428 4264
rect 11422 4224 11428 4236
rect 11480 4224 11486 4276
rect 9398 4196 9404 4208
rect 9359 4168 9404 4196
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 9214 4060 9220 4072
rect 9127 4032 9220 4060
rect 9214 4020 9220 4032
rect 9272 4060 9278 4072
rect 11238 4060 11244 4072
rect 9272 4032 9812 4060
rect 11151 4032 11244 4060
rect 9272 4020 9278 4032
rect 9784 3933 9812 4032
rect 11238 4020 11244 4032
rect 11296 4060 11302 4072
rect 11296 4032 11744 4060
rect 11296 4020 11302 4032
rect 11716 3936 11744 4032
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3924 9827 3927
rect 10042 3924 10048 3936
rect 9815 3896 10048 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11756 3896 11805 3924
rect 11756 3884 11762 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11793 3887 11851 3893
rect 1104 3834 12880 3856
rect 1104 3782 5648 3834
rect 5700 3782 5712 3834
rect 5764 3782 5776 3834
rect 5828 3782 5840 3834
rect 5892 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 12880 3834
rect 1104 3760 12880 3782
rect 8665 3723 8723 3729
rect 8665 3689 8677 3723
rect 8711 3720 8723 3723
rect 9398 3720 9404 3732
rect 8711 3692 9404 3720
rect 8711 3689 8723 3692
rect 8665 3683 8723 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 9548 3692 10517 3720
rect 9548 3680 9554 3692
rect 10505 3689 10517 3692
rect 10551 3720 10563 3723
rect 10686 3720 10692 3732
rect 10551 3692 10692 3720
rect 10551 3689 10563 3692
rect 10505 3683 10563 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 11057 3383 11115 3389
rect 11057 3349 11069 3383
rect 11103 3380 11115 3383
rect 11238 3380 11244 3392
rect 11103 3352 11244 3380
rect 11103 3349 11115 3352
rect 11057 3343 11115 3349
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 1104 3290 12880 3312
rect 1104 3238 3315 3290
rect 3367 3238 3379 3290
rect 3431 3238 3443 3290
rect 3495 3238 3507 3290
rect 3559 3238 7982 3290
rect 8034 3238 8046 3290
rect 8098 3238 8110 3290
rect 8162 3238 8174 3290
rect 8226 3238 12880 3290
rect 1104 3216 12880 3238
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 10045 3043 10103 3049
rect 8159 3012 9076 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 9048 2984 9076 3012
rect 10045 3009 10057 3043
rect 10091 3040 10103 3043
rect 10134 3040 10140 3052
rect 10091 3012 10140 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10134 3000 10140 3012
rect 10192 3040 10198 3052
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10192 3012 10701 3040
rect 10192 3000 10198 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2941 8631 2975
rect 9030 2972 9036 2984
rect 8991 2944 9036 2972
rect 8573 2935 8631 2941
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 7834 2836 7840 2848
rect 6052 2808 7840 2836
rect 6052 2796 6058 2808
rect 7834 2796 7840 2808
rect 7892 2836 7898 2848
rect 8389 2839 8447 2845
rect 8389 2836 8401 2839
rect 7892 2808 8401 2836
rect 7892 2796 7898 2808
rect 8389 2805 8401 2808
rect 8435 2836 8447 2839
rect 8588 2836 8616 2935
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9398 2972 9404 2984
rect 9359 2944 9404 2972
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 9766 2972 9772 2984
rect 9727 2944 9772 2972
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 8435 2808 8616 2836
rect 10413 2839 10471 2845
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 10413 2805 10425 2839
rect 10459 2836 10471 2839
rect 10686 2836 10692 2848
rect 10459 2808 10692 2836
rect 10459 2805 10471 2808
rect 10413 2799 10471 2805
rect 10686 2796 10692 2808
rect 10744 2836 10750 2848
rect 12342 2836 12348 2848
rect 10744 2808 12348 2836
rect 10744 2796 10750 2808
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 1104 2746 12880 2768
rect 1104 2694 5648 2746
rect 5700 2694 5712 2746
rect 5764 2694 5776 2746
rect 5828 2694 5840 2746
rect 5892 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 12880 2746
rect 1104 2672 12880 2694
rect 10962 2632 10968 2644
rect 10923 2604 10968 2632
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11698 2632 11704 2644
rect 11659 2604 11704 2632
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 11238 2496 11244 2508
rect 10643 2468 11244 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 11238 2456 11244 2468
rect 11296 2456 11302 2508
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 11020 2400 11069 2428
rect 11020 2388 11026 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8444 2264 8585 2292
rect 8444 2252 8450 2264
rect 8573 2261 8585 2264
rect 8619 2292 8631 2295
rect 9766 2292 9772 2304
rect 8619 2264 9772 2292
rect 8619 2261 8631 2264
rect 8573 2255 8631 2261
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 1104 2202 12880 2224
rect 1104 2150 3315 2202
rect 3367 2150 3379 2202
rect 3431 2150 3443 2202
rect 3495 2150 3507 2202
rect 3559 2150 7982 2202
rect 8034 2150 8046 2202
rect 8098 2150 8110 2202
rect 8162 2150 8174 2202
rect 8226 2150 12880 2202
rect 1104 2128 12880 2150
<< via1 >>
rect 3315 106598 3367 106650
rect 3379 106598 3431 106650
rect 3443 106598 3495 106650
rect 3507 106598 3559 106650
rect 7982 106598 8034 106650
rect 8046 106598 8098 106650
rect 8110 106598 8162 106650
rect 8174 106598 8226 106650
rect 5648 106054 5700 106106
rect 5712 106054 5764 106106
rect 5776 106054 5828 106106
rect 5840 106054 5892 106106
rect 10315 106054 10367 106106
rect 10379 106054 10431 106106
rect 10443 106054 10495 106106
rect 10507 106054 10559 106106
rect 3315 105510 3367 105562
rect 3379 105510 3431 105562
rect 3443 105510 3495 105562
rect 3507 105510 3559 105562
rect 7982 105510 8034 105562
rect 8046 105510 8098 105562
rect 8110 105510 8162 105562
rect 8174 105510 8226 105562
rect 5648 104966 5700 105018
rect 5712 104966 5764 105018
rect 5776 104966 5828 105018
rect 5840 104966 5892 105018
rect 10315 104966 10367 105018
rect 10379 104966 10431 105018
rect 10443 104966 10495 105018
rect 10507 104966 10559 105018
rect 3315 104422 3367 104474
rect 3379 104422 3431 104474
rect 3443 104422 3495 104474
rect 3507 104422 3559 104474
rect 7982 104422 8034 104474
rect 8046 104422 8098 104474
rect 8110 104422 8162 104474
rect 8174 104422 8226 104474
rect 5648 103878 5700 103930
rect 5712 103878 5764 103930
rect 5776 103878 5828 103930
rect 5840 103878 5892 103930
rect 10315 103878 10367 103930
rect 10379 103878 10431 103930
rect 10443 103878 10495 103930
rect 10507 103878 10559 103930
rect 3315 103334 3367 103386
rect 3379 103334 3431 103386
rect 3443 103334 3495 103386
rect 3507 103334 3559 103386
rect 7982 103334 8034 103386
rect 8046 103334 8098 103386
rect 8110 103334 8162 103386
rect 8174 103334 8226 103386
rect 5648 102790 5700 102842
rect 5712 102790 5764 102842
rect 5776 102790 5828 102842
rect 5840 102790 5892 102842
rect 10315 102790 10367 102842
rect 10379 102790 10431 102842
rect 10443 102790 10495 102842
rect 10507 102790 10559 102842
rect 3315 102246 3367 102298
rect 3379 102246 3431 102298
rect 3443 102246 3495 102298
rect 3507 102246 3559 102298
rect 7982 102246 8034 102298
rect 8046 102246 8098 102298
rect 8110 102246 8162 102298
rect 8174 102246 8226 102298
rect 5648 101702 5700 101754
rect 5712 101702 5764 101754
rect 5776 101702 5828 101754
rect 5840 101702 5892 101754
rect 10315 101702 10367 101754
rect 10379 101702 10431 101754
rect 10443 101702 10495 101754
rect 10507 101702 10559 101754
rect 3315 101158 3367 101210
rect 3379 101158 3431 101210
rect 3443 101158 3495 101210
rect 3507 101158 3559 101210
rect 7982 101158 8034 101210
rect 8046 101158 8098 101210
rect 8110 101158 8162 101210
rect 8174 101158 8226 101210
rect 5648 100614 5700 100666
rect 5712 100614 5764 100666
rect 5776 100614 5828 100666
rect 5840 100614 5892 100666
rect 10315 100614 10367 100666
rect 10379 100614 10431 100666
rect 10443 100614 10495 100666
rect 10507 100614 10559 100666
rect 3315 100070 3367 100122
rect 3379 100070 3431 100122
rect 3443 100070 3495 100122
rect 3507 100070 3559 100122
rect 7982 100070 8034 100122
rect 8046 100070 8098 100122
rect 8110 100070 8162 100122
rect 8174 100070 8226 100122
rect 5648 99526 5700 99578
rect 5712 99526 5764 99578
rect 5776 99526 5828 99578
rect 5840 99526 5892 99578
rect 10315 99526 10367 99578
rect 10379 99526 10431 99578
rect 10443 99526 10495 99578
rect 10507 99526 10559 99578
rect 3315 98982 3367 99034
rect 3379 98982 3431 99034
rect 3443 98982 3495 99034
rect 3507 98982 3559 99034
rect 7982 98982 8034 99034
rect 8046 98982 8098 99034
rect 8110 98982 8162 99034
rect 8174 98982 8226 99034
rect 5648 98438 5700 98490
rect 5712 98438 5764 98490
rect 5776 98438 5828 98490
rect 5840 98438 5892 98490
rect 10315 98438 10367 98490
rect 10379 98438 10431 98490
rect 10443 98438 10495 98490
rect 10507 98438 10559 98490
rect 3315 97894 3367 97946
rect 3379 97894 3431 97946
rect 3443 97894 3495 97946
rect 3507 97894 3559 97946
rect 7982 97894 8034 97946
rect 8046 97894 8098 97946
rect 8110 97894 8162 97946
rect 8174 97894 8226 97946
rect 11428 97835 11480 97844
rect 11428 97801 11437 97835
rect 11437 97801 11471 97835
rect 11471 97801 11480 97835
rect 11428 97792 11480 97801
rect 11244 97631 11296 97640
rect 11244 97597 11253 97631
rect 11253 97597 11287 97631
rect 11287 97597 11296 97631
rect 11244 97588 11296 97597
rect 5648 97350 5700 97402
rect 5712 97350 5764 97402
rect 5776 97350 5828 97402
rect 5840 97350 5892 97402
rect 10315 97350 10367 97402
rect 10379 97350 10431 97402
rect 10443 97350 10495 97402
rect 10507 97350 10559 97402
rect 3315 96806 3367 96858
rect 3379 96806 3431 96858
rect 3443 96806 3495 96858
rect 3507 96806 3559 96858
rect 7982 96806 8034 96858
rect 8046 96806 8098 96858
rect 8110 96806 8162 96858
rect 8174 96806 8226 96858
rect 5648 96262 5700 96314
rect 5712 96262 5764 96314
rect 5776 96262 5828 96314
rect 5840 96262 5892 96314
rect 10315 96262 10367 96314
rect 10379 96262 10431 96314
rect 10443 96262 10495 96314
rect 10507 96262 10559 96314
rect 3315 95718 3367 95770
rect 3379 95718 3431 95770
rect 3443 95718 3495 95770
rect 3507 95718 3559 95770
rect 7982 95718 8034 95770
rect 8046 95718 8098 95770
rect 8110 95718 8162 95770
rect 8174 95718 8226 95770
rect 5648 95174 5700 95226
rect 5712 95174 5764 95226
rect 5776 95174 5828 95226
rect 5840 95174 5892 95226
rect 10315 95174 10367 95226
rect 10379 95174 10431 95226
rect 10443 95174 10495 95226
rect 10507 95174 10559 95226
rect 11060 94936 11112 94988
rect 11152 94911 11204 94920
rect 11152 94877 11161 94911
rect 11161 94877 11195 94911
rect 11195 94877 11204 94911
rect 11152 94868 11204 94877
rect 11244 94800 11296 94852
rect 3315 94630 3367 94682
rect 3379 94630 3431 94682
rect 3443 94630 3495 94682
rect 3507 94630 3559 94682
rect 7982 94630 8034 94682
rect 8046 94630 8098 94682
rect 8110 94630 8162 94682
rect 8174 94630 8226 94682
rect 11152 94571 11204 94580
rect 11152 94537 11161 94571
rect 11161 94537 11195 94571
rect 11195 94537 11204 94571
rect 11152 94528 11204 94537
rect 11060 94256 11112 94308
rect 5648 94086 5700 94138
rect 5712 94086 5764 94138
rect 5776 94086 5828 94138
rect 5840 94086 5892 94138
rect 10315 94086 10367 94138
rect 10379 94086 10431 94138
rect 10443 94086 10495 94138
rect 10507 94086 10559 94138
rect 3315 93542 3367 93594
rect 3379 93542 3431 93594
rect 3443 93542 3495 93594
rect 3507 93542 3559 93594
rect 7982 93542 8034 93594
rect 8046 93542 8098 93594
rect 8110 93542 8162 93594
rect 8174 93542 8226 93594
rect 5648 92998 5700 93050
rect 5712 92998 5764 93050
rect 5776 92998 5828 93050
rect 5840 92998 5892 93050
rect 10315 92998 10367 93050
rect 10379 92998 10431 93050
rect 10443 92998 10495 93050
rect 10507 92998 10559 93050
rect 3315 92454 3367 92506
rect 3379 92454 3431 92506
rect 3443 92454 3495 92506
rect 3507 92454 3559 92506
rect 7982 92454 8034 92506
rect 8046 92454 8098 92506
rect 8110 92454 8162 92506
rect 8174 92454 8226 92506
rect 5648 91910 5700 91962
rect 5712 91910 5764 91962
rect 5776 91910 5828 91962
rect 5840 91910 5892 91962
rect 10315 91910 10367 91962
rect 10379 91910 10431 91962
rect 10443 91910 10495 91962
rect 10507 91910 10559 91962
rect 3315 91366 3367 91418
rect 3379 91366 3431 91418
rect 3443 91366 3495 91418
rect 3507 91366 3559 91418
rect 7982 91366 8034 91418
rect 8046 91366 8098 91418
rect 8110 91366 8162 91418
rect 8174 91366 8226 91418
rect 5648 90822 5700 90874
rect 5712 90822 5764 90874
rect 5776 90822 5828 90874
rect 5840 90822 5892 90874
rect 10315 90822 10367 90874
rect 10379 90822 10431 90874
rect 10443 90822 10495 90874
rect 10507 90822 10559 90874
rect 3315 90278 3367 90330
rect 3379 90278 3431 90330
rect 3443 90278 3495 90330
rect 3507 90278 3559 90330
rect 7982 90278 8034 90330
rect 8046 90278 8098 90330
rect 8110 90278 8162 90330
rect 8174 90278 8226 90330
rect 5648 89734 5700 89786
rect 5712 89734 5764 89786
rect 5776 89734 5828 89786
rect 5840 89734 5892 89786
rect 10315 89734 10367 89786
rect 10379 89734 10431 89786
rect 10443 89734 10495 89786
rect 10507 89734 10559 89786
rect 3315 89190 3367 89242
rect 3379 89190 3431 89242
rect 3443 89190 3495 89242
rect 3507 89190 3559 89242
rect 7982 89190 8034 89242
rect 8046 89190 8098 89242
rect 8110 89190 8162 89242
rect 8174 89190 8226 89242
rect 5648 88646 5700 88698
rect 5712 88646 5764 88698
rect 5776 88646 5828 88698
rect 5840 88646 5892 88698
rect 10315 88646 10367 88698
rect 10379 88646 10431 88698
rect 10443 88646 10495 88698
rect 10507 88646 10559 88698
rect 3315 88102 3367 88154
rect 3379 88102 3431 88154
rect 3443 88102 3495 88154
rect 3507 88102 3559 88154
rect 7982 88102 8034 88154
rect 8046 88102 8098 88154
rect 8110 88102 8162 88154
rect 8174 88102 8226 88154
rect 5648 87558 5700 87610
rect 5712 87558 5764 87610
rect 5776 87558 5828 87610
rect 5840 87558 5892 87610
rect 10315 87558 10367 87610
rect 10379 87558 10431 87610
rect 10443 87558 10495 87610
rect 10507 87558 10559 87610
rect 3315 87014 3367 87066
rect 3379 87014 3431 87066
rect 3443 87014 3495 87066
rect 3507 87014 3559 87066
rect 7982 87014 8034 87066
rect 8046 87014 8098 87066
rect 8110 87014 8162 87066
rect 8174 87014 8226 87066
rect 5648 86470 5700 86522
rect 5712 86470 5764 86522
rect 5776 86470 5828 86522
rect 5840 86470 5892 86522
rect 10315 86470 10367 86522
rect 10379 86470 10431 86522
rect 10443 86470 10495 86522
rect 10507 86470 10559 86522
rect 3315 85926 3367 85978
rect 3379 85926 3431 85978
rect 3443 85926 3495 85978
rect 3507 85926 3559 85978
rect 7982 85926 8034 85978
rect 8046 85926 8098 85978
rect 8110 85926 8162 85978
rect 8174 85926 8226 85978
rect 5648 85382 5700 85434
rect 5712 85382 5764 85434
rect 5776 85382 5828 85434
rect 5840 85382 5892 85434
rect 10315 85382 10367 85434
rect 10379 85382 10431 85434
rect 10443 85382 10495 85434
rect 10507 85382 10559 85434
rect 10692 85280 10744 85332
rect 11520 85187 11572 85196
rect 11520 85153 11529 85187
rect 11529 85153 11563 85187
rect 11563 85153 11572 85187
rect 11520 85144 11572 85153
rect 3315 84838 3367 84890
rect 3379 84838 3431 84890
rect 3443 84838 3495 84890
rect 3507 84838 3559 84890
rect 7982 84838 8034 84890
rect 8046 84838 8098 84890
rect 8110 84838 8162 84890
rect 8174 84838 8226 84890
rect 11520 84779 11572 84788
rect 11520 84745 11529 84779
rect 11529 84745 11563 84779
rect 11563 84745 11572 84779
rect 11520 84736 11572 84745
rect 11796 84736 11848 84788
rect 5648 84294 5700 84346
rect 5712 84294 5764 84346
rect 5776 84294 5828 84346
rect 5840 84294 5892 84346
rect 10315 84294 10367 84346
rect 10379 84294 10431 84346
rect 10443 84294 10495 84346
rect 10507 84294 10559 84346
rect 3315 83750 3367 83802
rect 3379 83750 3431 83802
rect 3443 83750 3495 83802
rect 3507 83750 3559 83802
rect 7982 83750 8034 83802
rect 8046 83750 8098 83802
rect 8110 83750 8162 83802
rect 8174 83750 8226 83802
rect 5648 83206 5700 83258
rect 5712 83206 5764 83258
rect 5776 83206 5828 83258
rect 5840 83206 5892 83258
rect 10315 83206 10367 83258
rect 10379 83206 10431 83258
rect 10443 83206 10495 83258
rect 10507 83206 10559 83258
rect 3315 82662 3367 82714
rect 3379 82662 3431 82714
rect 3443 82662 3495 82714
rect 3507 82662 3559 82714
rect 7982 82662 8034 82714
rect 8046 82662 8098 82714
rect 8110 82662 8162 82714
rect 8174 82662 8226 82714
rect 5648 82118 5700 82170
rect 5712 82118 5764 82170
rect 5776 82118 5828 82170
rect 5840 82118 5892 82170
rect 10315 82118 10367 82170
rect 10379 82118 10431 82170
rect 10443 82118 10495 82170
rect 10507 82118 10559 82170
rect 3315 81574 3367 81626
rect 3379 81574 3431 81626
rect 3443 81574 3495 81626
rect 3507 81574 3559 81626
rect 7982 81574 8034 81626
rect 8046 81574 8098 81626
rect 8110 81574 8162 81626
rect 8174 81574 8226 81626
rect 5648 81030 5700 81082
rect 5712 81030 5764 81082
rect 5776 81030 5828 81082
rect 5840 81030 5892 81082
rect 10315 81030 10367 81082
rect 10379 81030 10431 81082
rect 10443 81030 10495 81082
rect 10507 81030 10559 81082
rect 11796 80971 11848 80980
rect 11796 80937 11805 80971
rect 11805 80937 11839 80971
rect 11839 80937 11848 80971
rect 11796 80928 11848 80937
rect 11152 80835 11204 80844
rect 11152 80801 11161 80835
rect 11161 80801 11195 80835
rect 11195 80801 11204 80835
rect 11152 80792 11204 80801
rect 11336 80767 11388 80776
rect 11336 80733 11345 80767
rect 11345 80733 11379 80767
rect 11379 80733 11388 80767
rect 11336 80724 11388 80733
rect 3315 80486 3367 80538
rect 3379 80486 3431 80538
rect 3443 80486 3495 80538
rect 3507 80486 3559 80538
rect 7982 80486 8034 80538
rect 8046 80486 8098 80538
rect 8110 80486 8162 80538
rect 8174 80486 8226 80538
rect 11152 80427 11204 80436
rect 11152 80393 11161 80427
rect 11161 80393 11195 80427
rect 11195 80393 11204 80427
rect 11152 80384 11204 80393
rect 11152 80044 11204 80096
rect 11336 80044 11388 80096
rect 5648 79942 5700 79994
rect 5712 79942 5764 79994
rect 5776 79942 5828 79994
rect 5840 79942 5892 79994
rect 10315 79942 10367 79994
rect 10379 79942 10431 79994
rect 10443 79942 10495 79994
rect 10507 79942 10559 79994
rect 3315 79398 3367 79450
rect 3379 79398 3431 79450
rect 3443 79398 3495 79450
rect 3507 79398 3559 79450
rect 7982 79398 8034 79450
rect 8046 79398 8098 79450
rect 8110 79398 8162 79450
rect 8174 79398 8226 79450
rect 5648 78854 5700 78906
rect 5712 78854 5764 78906
rect 5776 78854 5828 78906
rect 5840 78854 5892 78906
rect 10315 78854 10367 78906
rect 10379 78854 10431 78906
rect 10443 78854 10495 78906
rect 10507 78854 10559 78906
rect 3315 78310 3367 78362
rect 3379 78310 3431 78362
rect 3443 78310 3495 78362
rect 3507 78310 3559 78362
rect 7982 78310 8034 78362
rect 8046 78310 8098 78362
rect 8110 78310 8162 78362
rect 8174 78310 8226 78362
rect 5648 77766 5700 77818
rect 5712 77766 5764 77818
rect 5776 77766 5828 77818
rect 5840 77766 5892 77818
rect 10315 77766 10367 77818
rect 10379 77766 10431 77818
rect 10443 77766 10495 77818
rect 10507 77766 10559 77818
rect 3315 77222 3367 77274
rect 3379 77222 3431 77274
rect 3443 77222 3495 77274
rect 3507 77222 3559 77274
rect 7982 77222 8034 77274
rect 8046 77222 8098 77274
rect 8110 77222 8162 77274
rect 8174 77222 8226 77274
rect 5648 76678 5700 76730
rect 5712 76678 5764 76730
rect 5776 76678 5828 76730
rect 5840 76678 5892 76730
rect 10315 76678 10367 76730
rect 10379 76678 10431 76730
rect 10443 76678 10495 76730
rect 10507 76678 10559 76730
rect 3315 76134 3367 76186
rect 3379 76134 3431 76186
rect 3443 76134 3495 76186
rect 3507 76134 3559 76186
rect 7982 76134 8034 76186
rect 8046 76134 8098 76186
rect 8110 76134 8162 76186
rect 8174 76134 8226 76186
rect 5648 75590 5700 75642
rect 5712 75590 5764 75642
rect 5776 75590 5828 75642
rect 5840 75590 5892 75642
rect 10315 75590 10367 75642
rect 10379 75590 10431 75642
rect 10443 75590 10495 75642
rect 10507 75590 10559 75642
rect 3315 75046 3367 75098
rect 3379 75046 3431 75098
rect 3443 75046 3495 75098
rect 3507 75046 3559 75098
rect 7982 75046 8034 75098
rect 8046 75046 8098 75098
rect 8110 75046 8162 75098
rect 8174 75046 8226 75098
rect 5648 74502 5700 74554
rect 5712 74502 5764 74554
rect 5776 74502 5828 74554
rect 5840 74502 5892 74554
rect 10315 74502 10367 74554
rect 10379 74502 10431 74554
rect 10443 74502 10495 74554
rect 10507 74502 10559 74554
rect 3315 73958 3367 74010
rect 3379 73958 3431 74010
rect 3443 73958 3495 74010
rect 3507 73958 3559 74010
rect 7982 73958 8034 74010
rect 8046 73958 8098 74010
rect 8110 73958 8162 74010
rect 8174 73958 8226 74010
rect 5648 73414 5700 73466
rect 5712 73414 5764 73466
rect 5776 73414 5828 73466
rect 5840 73414 5892 73466
rect 10315 73414 10367 73466
rect 10379 73414 10431 73466
rect 10443 73414 10495 73466
rect 10507 73414 10559 73466
rect 3315 72870 3367 72922
rect 3379 72870 3431 72922
rect 3443 72870 3495 72922
rect 3507 72870 3559 72922
rect 7982 72870 8034 72922
rect 8046 72870 8098 72922
rect 8110 72870 8162 72922
rect 8174 72870 8226 72922
rect 5648 72326 5700 72378
rect 5712 72326 5764 72378
rect 5776 72326 5828 72378
rect 5840 72326 5892 72378
rect 10315 72326 10367 72378
rect 10379 72326 10431 72378
rect 10443 72326 10495 72378
rect 10507 72326 10559 72378
rect 3315 71782 3367 71834
rect 3379 71782 3431 71834
rect 3443 71782 3495 71834
rect 3507 71782 3559 71834
rect 7982 71782 8034 71834
rect 8046 71782 8098 71834
rect 8110 71782 8162 71834
rect 8174 71782 8226 71834
rect 10968 71680 11020 71732
rect 11244 71519 11296 71528
rect 11244 71485 11253 71519
rect 11253 71485 11287 71519
rect 11287 71485 11296 71519
rect 11796 71519 11848 71528
rect 11244 71476 11296 71485
rect 11796 71485 11805 71519
rect 11805 71485 11839 71519
rect 11839 71485 11848 71519
rect 11796 71476 11848 71485
rect 5648 71238 5700 71290
rect 5712 71238 5764 71290
rect 5776 71238 5828 71290
rect 5840 71238 5892 71290
rect 10315 71238 10367 71290
rect 10379 71238 10431 71290
rect 10443 71238 10495 71290
rect 10507 71238 10559 71290
rect 3315 70694 3367 70746
rect 3379 70694 3431 70746
rect 3443 70694 3495 70746
rect 3507 70694 3559 70746
rect 7982 70694 8034 70746
rect 8046 70694 8098 70746
rect 8110 70694 8162 70746
rect 8174 70694 8226 70746
rect 5648 70150 5700 70202
rect 5712 70150 5764 70202
rect 5776 70150 5828 70202
rect 5840 70150 5892 70202
rect 10315 70150 10367 70202
rect 10379 70150 10431 70202
rect 10443 70150 10495 70202
rect 10507 70150 10559 70202
rect 3315 69606 3367 69658
rect 3379 69606 3431 69658
rect 3443 69606 3495 69658
rect 3507 69606 3559 69658
rect 7982 69606 8034 69658
rect 8046 69606 8098 69658
rect 8110 69606 8162 69658
rect 8174 69606 8226 69658
rect 5648 69062 5700 69114
rect 5712 69062 5764 69114
rect 5776 69062 5828 69114
rect 5840 69062 5892 69114
rect 10315 69062 10367 69114
rect 10379 69062 10431 69114
rect 10443 69062 10495 69114
rect 10507 69062 10559 69114
rect 3315 68518 3367 68570
rect 3379 68518 3431 68570
rect 3443 68518 3495 68570
rect 3507 68518 3559 68570
rect 7982 68518 8034 68570
rect 8046 68518 8098 68570
rect 8110 68518 8162 68570
rect 8174 68518 8226 68570
rect 5648 67974 5700 68026
rect 5712 67974 5764 68026
rect 5776 67974 5828 68026
rect 5840 67974 5892 68026
rect 10315 67974 10367 68026
rect 10379 67974 10431 68026
rect 10443 67974 10495 68026
rect 10507 67974 10559 68026
rect 3315 67430 3367 67482
rect 3379 67430 3431 67482
rect 3443 67430 3495 67482
rect 3507 67430 3559 67482
rect 7982 67430 8034 67482
rect 8046 67430 8098 67482
rect 8110 67430 8162 67482
rect 8174 67430 8226 67482
rect 5648 66886 5700 66938
rect 5712 66886 5764 66938
rect 5776 66886 5828 66938
rect 5840 66886 5892 66938
rect 10315 66886 10367 66938
rect 10379 66886 10431 66938
rect 10443 66886 10495 66938
rect 10507 66886 10559 66938
rect 11796 66827 11848 66836
rect 11796 66793 11805 66827
rect 11805 66793 11839 66827
rect 11839 66793 11848 66827
rect 11796 66784 11848 66793
rect 11428 66648 11480 66700
rect 11336 66623 11388 66632
rect 11336 66589 11345 66623
rect 11345 66589 11379 66623
rect 11379 66589 11388 66623
rect 11336 66580 11388 66589
rect 3315 66342 3367 66394
rect 3379 66342 3431 66394
rect 3443 66342 3495 66394
rect 3507 66342 3559 66394
rect 7982 66342 8034 66394
rect 8046 66342 8098 66394
rect 8110 66342 8162 66394
rect 8174 66342 8226 66394
rect 11428 66240 11480 66292
rect 10140 65968 10192 66020
rect 11336 65968 11388 66020
rect 5648 65798 5700 65850
rect 5712 65798 5764 65850
rect 5776 65798 5828 65850
rect 5840 65798 5892 65850
rect 10315 65798 10367 65850
rect 10379 65798 10431 65850
rect 10443 65798 10495 65850
rect 10507 65798 10559 65850
rect 3315 65254 3367 65306
rect 3379 65254 3431 65306
rect 3443 65254 3495 65306
rect 3507 65254 3559 65306
rect 7982 65254 8034 65306
rect 8046 65254 8098 65306
rect 8110 65254 8162 65306
rect 8174 65254 8226 65306
rect 5648 64710 5700 64762
rect 5712 64710 5764 64762
rect 5776 64710 5828 64762
rect 5840 64710 5892 64762
rect 10315 64710 10367 64762
rect 10379 64710 10431 64762
rect 10443 64710 10495 64762
rect 10507 64710 10559 64762
rect 3315 64166 3367 64218
rect 3379 64166 3431 64218
rect 3443 64166 3495 64218
rect 3507 64166 3559 64218
rect 7982 64166 8034 64218
rect 8046 64166 8098 64218
rect 8110 64166 8162 64218
rect 8174 64166 8226 64218
rect 5648 63622 5700 63674
rect 5712 63622 5764 63674
rect 5776 63622 5828 63674
rect 5840 63622 5892 63674
rect 10315 63622 10367 63674
rect 10379 63622 10431 63674
rect 10443 63622 10495 63674
rect 10507 63622 10559 63674
rect 3315 63078 3367 63130
rect 3379 63078 3431 63130
rect 3443 63078 3495 63130
rect 3507 63078 3559 63130
rect 7982 63078 8034 63130
rect 8046 63078 8098 63130
rect 8110 63078 8162 63130
rect 8174 63078 8226 63130
rect 5648 62534 5700 62586
rect 5712 62534 5764 62586
rect 5776 62534 5828 62586
rect 5840 62534 5892 62586
rect 10315 62534 10367 62586
rect 10379 62534 10431 62586
rect 10443 62534 10495 62586
rect 10507 62534 10559 62586
rect 3315 61990 3367 62042
rect 3379 61990 3431 62042
rect 3443 61990 3495 62042
rect 3507 61990 3559 62042
rect 7982 61990 8034 62042
rect 8046 61990 8098 62042
rect 8110 61990 8162 62042
rect 8174 61990 8226 62042
rect 5648 61446 5700 61498
rect 5712 61446 5764 61498
rect 5776 61446 5828 61498
rect 5840 61446 5892 61498
rect 10315 61446 10367 61498
rect 10379 61446 10431 61498
rect 10443 61446 10495 61498
rect 10507 61446 10559 61498
rect 3315 60902 3367 60954
rect 3379 60902 3431 60954
rect 3443 60902 3495 60954
rect 3507 60902 3559 60954
rect 7982 60902 8034 60954
rect 8046 60902 8098 60954
rect 8110 60902 8162 60954
rect 8174 60902 8226 60954
rect 5648 60358 5700 60410
rect 5712 60358 5764 60410
rect 5776 60358 5828 60410
rect 5840 60358 5892 60410
rect 10315 60358 10367 60410
rect 10379 60358 10431 60410
rect 10443 60358 10495 60410
rect 10507 60358 10559 60410
rect 3315 59814 3367 59866
rect 3379 59814 3431 59866
rect 3443 59814 3495 59866
rect 3507 59814 3559 59866
rect 7982 59814 8034 59866
rect 8046 59814 8098 59866
rect 8110 59814 8162 59866
rect 8174 59814 8226 59866
rect 5648 59270 5700 59322
rect 5712 59270 5764 59322
rect 5776 59270 5828 59322
rect 5840 59270 5892 59322
rect 10315 59270 10367 59322
rect 10379 59270 10431 59322
rect 10443 59270 10495 59322
rect 10507 59270 10559 59322
rect 3315 58726 3367 58778
rect 3379 58726 3431 58778
rect 3443 58726 3495 58778
rect 3507 58726 3559 58778
rect 7982 58726 8034 58778
rect 8046 58726 8098 58778
rect 8110 58726 8162 58778
rect 8174 58726 8226 58778
rect 11428 58667 11480 58676
rect 11428 58633 11437 58667
rect 11437 58633 11471 58667
rect 11471 58633 11480 58667
rect 11428 58624 11480 58633
rect 11244 58463 11296 58472
rect 11244 58429 11253 58463
rect 11253 58429 11287 58463
rect 11287 58429 11296 58463
rect 11796 58463 11848 58472
rect 11244 58420 11296 58429
rect 11796 58429 11805 58463
rect 11805 58429 11839 58463
rect 11839 58429 11848 58463
rect 11796 58420 11848 58429
rect 5648 58182 5700 58234
rect 5712 58182 5764 58234
rect 5776 58182 5828 58234
rect 5840 58182 5892 58234
rect 10315 58182 10367 58234
rect 10379 58182 10431 58234
rect 10443 58182 10495 58234
rect 10507 58182 10559 58234
rect 3315 57638 3367 57690
rect 3379 57638 3431 57690
rect 3443 57638 3495 57690
rect 3507 57638 3559 57690
rect 7982 57638 8034 57690
rect 8046 57638 8098 57690
rect 8110 57638 8162 57690
rect 8174 57638 8226 57690
rect 5648 57094 5700 57146
rect 5712 57094 5764 57146
rect 5776 57094 5828 57146
rect 5840 57094 5892 57146
rect 10315 57094 10367 57146
rect 10379 57094 10431 57146
rect 10443 57094 10495 57146
rect 10507 57094 10559 57146
rect 3315 56550 3367 56602
rect 3379 56550 3431 56602
rect 3443 56550 3495 56602
rect 3507 56550 3559 56602
rect 7982 56550 8034 56602
rect 8046 56550 8098 56602
rect 8110 56550 8162 56602
rect 8174 56550 8226 56602
rect 5648 56006 5700 56058
rect 5712 56006 5764 56058
rect 5776 56006 5828 56058
rect 5840 56006 5892 56058
rect 10315 56006 10367 56058
rect 10379 56006 10431 56058
rect 10443 56006 10495 56058
rect 10507 56006 10559 56058
rect 3315 55462 3367 55514
rect 3379 55462 3431 55514
rect 3443 55462 3495 55514
rect 3507 55462 3559 55514
rect 7982 55462 8034 55514
rect 8046 55462 8098 55514
rect 8110 55462 8162 55514
rect 8174 55462 8226 55514
rect 5648 54918 5700 54970
rect 5712 54918 5764 54970
rect 5776 54918 5828 54970
rect 5840 54918 5892 54970
rect 10315 54918 10367 54970
rect 10379 54918 10431 54970
rect 10443 54918 10495 54970
rect 10507 54918 10559 54970
rect 3315 54374 3367 54426
rect 3379 54374 3431 54426
rect 3443 54374 3495 54426
rect 3507 54374 3559 54426
rect 7982 54374 8034 54426
rect 8046 54374 8098 54426
rect 8110 54374 8162 54426
rect 8174 54374 8226 54426
rect 5648 53830 5700 53882
rect 5712 53830 5764 53882
rect 5776 53830 5828 53882
rect 5840 53830 5892 53882
rect 10315 53830 10367 53882
rect 10379 53830 10431 53882
rect 10443 53830 10495 53882
rect 10507 53830 10559 53882
rect 11796 53771 11848 53780
rect 11796 53737 11805 53771
rect 11805 53737 11839 53771
rect 11839 53737 11848 53771
rect 11796 53728 11848 53737
rect 11428 53592 11480 53644
rect 11612 53524 11664 53576
rect 3315 53286 3367 53338
rect 3379 53286 3431 53338
rect 3443 53286 3495 53338
rect 3507 53286 3559 53338
rect 7982 53286 8034 53338
rect 8046 53286 8098 53338
rect 8110 53286 8162 53338
rect 8174 53286 8226 53338
rect 11428 53184 11480 53236
rect 11612 52887 11664 52896
rect 11612 52853 11621 52887
rect 11621 52853 11655 52887
rect 11655 52853 11664 52887
rect 11612 52844 11664 52853
rect 5648 52742 5700 52794
rect 5712 52742 5764 52794
rect 5776 52742 5828 52794
rect 5840 52742 5892 52794
rect 10315 52742 10367 52794
rect 10379 52742 10431 52794
rect 10443 52742 10495 52794
rect 10507 52742 10559 52794
rect 3315 52198 3367 52250
rect 3379 52198 3431 52250
rect 3443 52198 3495 52250
rect 3507 52198 3559 52250
rect 7982 52198 8034 52250
rect 8046 52198 8098 52250
rect 8110 52198 8162 52250
rect 8174 52198 8226 52250
rect 5648 51654 5700 51706
rect 5712 51654 5764 51706
rect 5776 51654 5828 51706
rect 5840 51654 5892 51706
rect 10315 51654 10367 51706
rect 10379 51654 10431 51706
rect 10443 51654 10495 51706
rect 10507 51654 10559 51706
rect 3315 51110 3367 51162
rect 3379 51110 3431 51162
rect 3443 51110 3495 51162
rect 3507 51110 3559 51162
rect 7982 51110 8034 51162
rect 8046 51110 8098 51162
rect 8110 51110 8162 51162
rect 8174 51110 8226 51162
rect 5648 50566 5700 50618
rect 5712 50566 5764 50618
rect 5776 50566 5828 50618
rect 5840 50566 5892 50618
rect 10315 50566 10367 50618
rect 10379 50566 10431 50618
rect 10443 50566 10495 50618
rect 10507 50566 10559 50618
rect 3315 50022 3367 50074
rect 3379 50022 3431 50074
rect 3443 50022 3495 50074
rect 3507 50022 3559 50074
rect 7982 50022 8034 50074
rect 8046 50022 8098 50074
rect 8110 50022 8162 50074
rect 8174 50022 8226 50074
rect 5648 49478 5700 49530
rect 5712 49478 5764 49530
rect 5776 49478 5828 49530
rect 5840 49478 5892 49530
rect 10315 49478 10367 49530
rect 10379 49478 10431 49530
rect 10443 49478 10495 49530
rect 10507 49478 10559 49530
rect 3315 48934 3367 48986
rect 3379 48934 3431 48986
rect 3443 48934 3495 48986
rect 3507 48934 3559 48986
rect 7982 48934 8034 48986
rect 8046 48934 8098 48986
rect 8110 48934 8162 48986
rect 8174 48934 8226 48986
rect 5648 48390 5700 48442
rect 5712 48390 5764 48442
rect 5776 48390 5828 48442
rect 5840 48390 5892 48442
rect 10315 48390 10367 48442
rect 10379 48390 10431 48442
rect 10443 48390 10495 48442
rect 10507 48390 10559 48442
rect 3315 47846 3367 47898
rect 3379 47846 3431 47898
rect 3443 47846 3495 47898
rect 3507 47846 3559 47898
rect 7982 47846 8034 47898
rect 8046 47846 8098 47898
rect 8110 47846 8162 47898
rect 8174 47846 8226 47898
rect 5648 47302 5700 47354
rect 5712 47302 5764 47354
rect 5776 47302 5828 47354
rect 5840 47302 5892 47354
rect 10315 47302 10367 47354
rect 10379 47302 10431 47354
rect 10443 47302 10495 47354
rect 10507 47302 10559 47354
rect 3315 46758 3367 46810
rect 3379 46758 3431 46810
rect 3443 46758 3495 46810
rect 3507 46758 3559 46810
rect 7982 46758 8034 46810
rect 8046 46758 8098 46810
rect 8110 46758 8162 46810
rect 8174 46758 8226 46810
rect 5648 46214 5700 46266
rect 5712 46214 5764 46266
rect 5776 46214 5828 46266
rect 5840 46214 5892 46266
rect 10315 46214 10367 46266
rect 10379 46214 10431 46266
rect 10443 46214 10495 46266
rect 10507 46214 10559 46266
rect 3315 45670 3367 45722
rect 3379 45670 3431 45722
rect 3443 45670 3495 45722
rect 3507 45670 3559 45722
rect 7982 45670 8034 45722
rect 8046 45670 8098 45722
rect 8110 45670 8162 45722
rect 8174 45670 8226 45722
rect 5648 45126 5700 45178
rect 5712 45126 5764 45178
rect 5776 45126 5828 45178
rect 5840 45126 5892 45178
rect 10315 45126 10367 45178
rect 10379 45126 10431 45178
rect 10443 45126 10495 45178
rect 10507 45126 10559 45178
rect 11704 45067 11756 45076
rect 11704 45033 11713 45067
rect 11713 45033 11747 45067
rect 11747 45033 11756 45067
rect 11704 45024 11756 45033
rect 11520 44931 11572 44940
rect 11520 44897 11529 44931
rect 11529 44897 11563 44931
rect 11563 44897 11572 44931
rect 11520 44888 11572 44897
rect 3315 44582 3367 44634
rect 3379 44582 3431 44634
rect 3443 44582 3495 44634
rect 3507 44582 3559 44634
rect 7982 44582 8034 44634
rect 8046 44582 8098 44634
rect 8110 44582 8162 44634
rect 8174 44582 8226 44634
rect 11520 44523 11572 44532
rect 11520 44489 11529 44523
rect 11529 44489 11563 44523
rect 11563 44489 11572 44523
rect 11520 44480 11572 44489
rect 5648 44038 5700 44090
rect 5712 44038 5764 44090
rect 5776 44038 5828 44090
rect 5840 44038 5892 44090
rect 10315 44038 10367 44090
rect 10379 44038 10431 44090
rect 10443 44038 10495 44090
rect 10507 44038 10559 44090
rect 3315 43494 3367 43546
rect 3379 43494 3431 43546
rect 3443 43494 3495 43546
rect 3507 43494 3559 43546
rect 7982 43494 8034 43546
rect 8046 43494 8098 43546
rect 8110 43494 8162 43546
rect 8174 43494 8226 43546
rect 5648 42950 5700 43002
rect 5712 42950 5764 43002
rect 5776 42950 5828 43002
rect 5840 42950 5892 43002
rect 10315 42950 10367 43002
rect 10379 42950 10431 43002
rect 10443 42950 10495 43002
rect 10507 42950 10559 43002
rect 3315 42406 3367 42458
rect 3379 42406 3431 42458
rect 3443 42406 3495 42458
rect 3507 42406 3559 42458
rect 7982 42406 8034 42458
rect 8046 42406 8098 42458
rect 8110 42406 8162 42458
rect 8174 42406 8226 42458
rect 5648 41862 5700 41914
rect 5712 41862 5764 41914
rect 5776 41862 5828 41914
rect 5840 41862 5892 41914
rect 10315 41862 10367 41914
rect 10379 41862 10431 41914
rect 10443 41862 10495 41914
rect 10507 41862 10559 41914
rect 3315 41318 3367 41370
rect 3379 41318 3431 41370
rect 3443 41318 3495 41370
rect 3507 41318 3559 41370
rect 7982 41318 8034 41370
rect 8046 41318 8098 41370
rect 8110 41318 8162 41370
rect 8174 41318 8226 41370
rect 5648 40774 5700 40826
rect 5712 40774 5764 40826
rect 5776 40774 5828 40826
rect 5840 40774 5892 40826
rect 10315 40774 10367 40826
rect 10379 40774 10431 40826
rect 10443 40774 10495 40826
rect 10507 40774 10559 40826
rect 3315 40230 3367 40282
rect 3379 40230 3431 40282
rect 3443 40230 3495 40282
rect 3507 40230 3559 40282
rect 7982 40230 8034 40282
rect 8046 40230 8098 40282
rect 8110 40230 8162 40282
rect 8174 40230 8226 40282
rect 10784 40171 10836 40180
rect 10784 40137 10793 40171
rect 10793 40137 10827 40171
rect 10827 40137 10836 40171
rect 11520 40171 11572 40180
rect 10784 40128 10836 40137
rect 11520 40137 11529 40171
rect 11529 40137 11563 40171
rect 11563 40137 11572 40171
rect 11520 40128 11572 40137
rect 11244 39924 11296 39976
rect 5648 39686 5700 39738
rect 5712 39686 5764 39738
rect 5776 39686 5828 39738
rect 5840 39686 5892 39738
rect 10315 39686 10367 39738
rect 10379 39686 10431 39738
rect 10443 39686 10495 39738
rect 10507 39686 10559 39738
rect 11244 39244 11296 39296
rect 3315 39142 3367 39194
rect 3379 39142 3431 39194
rect 3443 39142 3495 39194
rect 3507 39142 3559 39194
rect 7982 39142 8034 39194
rect 8046 39142 8098 39194
rect 8110 39142 8162 39194
rect 8174 39142 8226 39194
rect 5648 38598 5700 38650
rect 5712 38598 5764 38650
rect 5776 38598 5828 38650
rect 5840 38598 5892 38650
rect 10315 38598 10367 38650
rect 10379 38598 10431 38650
rect 10443 38598 10495 38650
rect 10507 38598 10559 38650
rect 3315 38054 3367 38106
rect 3379 38054 3431 38106
rect 3443 38054 3495 38106
rect 3507 38054 3559 38106
rect 7982 38054 8034 38106
rect 8046 38054 8098 38106
rect 8110 38054 8162 38106
rect 8174 38054 8226 38106
rect 5648 37510 5700 37562
rect 5712 37510 5764 37562
rect 5776 37510 5828 37562
rect 5840 37510 5892 37562
rect 10315 37510 10367 37562
rect 10379 37510 10431 37562
rect 10443 37510 10495 37562
rect 10507 37510 10559 37562
rect 3315 36966 3367 37018
rect 3379 36966 3431 37018
rect 3443 36966 3495 37018
rect 3507 36966 3559 37018
rect 7982 36966 8034 37018
rect 8046 36966 8098 37018
rect 8110 36966 8162 37018
rect 8174 36966 8226 37018
rect 5648 36422 5700 36474
rect 5712 36422 5764 36474
rect 5776 36422 5828 36474
rect 5840 36422 5892 36474
rect 10315 36422 10367 36474
rect 10379 36422 10431 36474
rect 10443 36422 10495 36474
rect 10507 36422 10559 36474
rect 3315 35878 3367 35930
rect 3379 35878 3431 35930
rect 3443 35878 3495 35930
rect 3507 35878 3559 35930
rect 7982 35878 8034 35930
rect 8046 35878 8098 35930
rect 8110 35878 8162 35930
rect 8174 35878 8226 35930
rect 5648 35334 5700 35386
rect 5712 35334 5764 35386
rect 5776 35334 5828 35386
rect 5840 35334 5892 35386
rect 10315 35334 10367 35386
rect 10379 35334 10431 35386
rect 10443 35334 10495 35386
rect 10507 35334 10559 35386
rect 3315 34790 3367 34842
rect 3379 34790 3431 34842
rect 3443 34790 3495 34842
rect 3507 34790 3559 34842
rect 7982 34790 8034 34842
rect 8046 34790 8098 34842
rect 8110 34790 8162 34842
rect 8174 34790 8226 34842
rect 5648 34246 5700 34298
rect 5712 34246 5764 34298
rect 5776 34246 5828 34298
rect 5840 34246 5892 34298
rect 10315 34246 10367 34298
rect 10379 34246 10431 34298
rect 10443 34246 10495 34298
rect 10507 34246 10559 34298
rect 3315 33702 3367 33754
rect 3379 33702 3431 33754
rect 3443 33702 3495 33754
rect 3507 33702 3559 33754
rect 7982 33702 8034 33754
rect 8046 33702 8098 33754
rect 8110 33702 8162 33754
rect 8174 33702 8226 33754
rect 5648 33158 5700 33210
rect 5712 33158 5764 33210
rect 5776 33158 5828 33210
rect 5840 33158 5892 33210
rect 10315 33158 10367 33210
rect 10379 33158 10431 33210
rect 10443 33158 10495 33210
rect 10507 33158 10559 33210
rect 3315 32614 3367 32666
rect 3379 32614 3431 32666
rect 3443 32614 3495 32666
rect 3507 32614 3559 32666
rect 7982 32614 8034 32666
rect 8046 32614 8098 32666
rect 8110 32614 8162 32666
rect 8174 32614 8226 32666
rect 5648 32070 5700 32122
rect 5712 32070 5764 32122
rect 5776 32070 5828 32122
rect 5840 32070 5892 32122
rect 10315 32070 10367 32122
rect 10379 32070 10431 32122
rect 10443 32070 10495 32122
rect 10507 32070 10559 32122
rect 3315 31526 3367 31578
rect 3379 31526 3431 31578
rect 3443 31526 3495 31578
rect 3507 31526 3559 31578
rect 7982 31526 8034 31578
rect 8046 31526 8098 31578
rect 8110 31526 8162 31578
rect 8174 31526 8226 31578
rect 11428 31467 11480 31476
rect 11428 31433 11437 31467
rect 11437 31433 11471 31467
rect 11471 31433 11480 31467
rect 11428 31424 11480 31433
rect 10968 31288 11020 31340
rect 5648 30982 5700 31034
rect 5712 30982 5764 31034
rect 5776 30982 5828 31034
rect 5840 30982 5892 31034
rect 10315 30982 10367 31034
rect 10379 30982 10431 31034
rect 10443 30982 10495 31034
rect 10507 30982 10559 31034
rect 3315 30438 3367 30490
rect 3379 30438 3431 30490
rect 3443 30438 3495 30490
rect 3507 30438 3559 30490
rect 7982 30438 8034 30490
rect 8046 30438 8098 30490
rect 8110 30438 8162 30490
rect 8174 30438 8226 30490
rect 5648 29894 5700 29946
rect 5712 29894 5764 29946
rect 5776 29894 5828 29946
rect 5840 29894 5892 29946
rect 10315 29894 10367 29946
rect 10379 29894 10431 29946
rect 10443 29894 10495 29946
rect 10507 29894 10559 29946
rect 3315 29350 3367 29402
rect 3379 29350 3431 29402
rect 3443 29350 3495 29402
rect 3507 29350 3559 29402
rect 7982 29350 8034 29402
rect 8046 29350 8098 29402
rect 8110 29350 8162 29402
rect 8174 29350 8226 29402
rect 5648 28806 5700 28858
rect 5712 28806 5764 28858
rect 5776 28806 5828 28858
rect 5840 28806 5892 28858
rect 10315 28806 10367 28858
rect 10379 28806 10431 28858
rect 10443 28806 10495 28858
rect 10507 28806 10559 28858
rect 3315 28262 3367 28314
rect 3379 28262 3431 28314
rect 3443 28262 3495 28314
rect 3507 28262 3559 28314
rect 7982 28262 8034 28314
rect 8046 28262 8098 28314
rect 8110 28262 8162 28314
rect 8174 28262 8226 28314
rect 5648 27718 5700 27770
rect 5712 27718 5764 27770
rect 5776 27718 5828 27770
rect 5840 27718 5892 27770
rect 10315 27718 10367 27770
rect 10379 27718 10431 27770
rect 10443 27718 10495 27770
rect 10507 27718 10559 27770
rect 3315 27174 3367 27226
rect 3379 27174 3431 27226
rect 3443 27174 3495 27226
rect 3507 27174 3559 27226
rect 7982 27174 8034 27226
rect 8046 27174 8098 27226
rect 8110 27174 8162 27226
rect 8174 27174 8226 27226
rect 10784 27115 10836 27124
rect 10784 27081 10793 27115
rect 10793 27081 10827 27115
rect 10827 27081 10836 27115
rect 10784 27072 10836 27081
rect 10968 27072 11020 27124
rect 10968 26868 11020 26920
rect 5648 26630 5700 26682
rect 5712 26630 5764 26682
rect 5776 26630 5828 26682
rect 5840 26630 5892 26682
rect 10315 26630 10367 26682
rect 10379 26630 10431 26682
rect 10443 26630 10495 26682
rect 10507 26630 10559 26682
rect 9404 26188 9456 26240
rect 10968 26188 11020 26240
rect 3315 26086 3367 26138
rect 3379 26086 3431 26138
rect 3443 26086 3495 26138
rect 3507 26086 3559 26138
rect 7982 26086 8034 26138
rect 8046 26086 8098 26138
rect 8110 26086 8162 26138
rect 8174 26086 8226 26138
rect 5648 25542 5700 25594
rect 5712 25542 5764 25594
rect 5776 25542 5828 25594
rect 5840 25542 5892 25594
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 3315 24998 3367 25050
rect 3379 24998 3431 25050
rect 3443 24998 3495 25050
rect 3507 24998 3559 25050
rect 7982 24998 8034 25050
rect 8046 24998 8098 25050
rect 8110 24998 8162 25050
rect 8174 24998 8226 25050
rect 5648 24454 5700 24506
rect 5712 24454 5764 24506
rect 5776 24454 5828 24506
rect 5840 24454 5892 24506
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 3315 23910 3367 23962
rect 3379 23910 3431 23962
rect 3443 23910 3495 23962
rect 3507 23910 3559 23962
rect 7982 23910 8034 23962
rect 8046 23910 8098 23962
rect 8110 23910 8162 23962
rect 8174 23910 8226 23962
rect 5648 23366 5700 23418
rect 5712 23366 5764 23418
rect 5776 23366 5828 23418
rect 5840 23366 5892 23418
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 3315 22822 3367 22874
rect 3379 22822 3431 22874
rect 3443 22822 3495 22874
rect 3507 22822 3559 22874
rect 7982 22822 8034 22874
rect 8046 22822 8098 22874
rect 8110 22822 8162 22874
rect 8174 22822 8226 22874
rect 5648 22278 5700 22330
rect 5712 22278 5764 22330
rect 5776 22278 5828 22330
rect 5840 22278 5892 22330
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 3315 21734 3367 21786
rect 3379 21734 3431 21786
rect 3443 21734 3495 21786
rect 3507 21734 3559 21786
rect 7982 21734 8034 21786
rect 8046 21734 8098 21786
rect 8110 21734 8162 21786
rect 8174 21734 8226 21786
rect 5648 21190 5700 21242
rect 5712 21190 5764 21242
rect 5776 21190 5828 21242
rect 5840 21190 5892 21242
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 3315 20646 3367 20698
rect 3379 20646 3431 20698
rect 3443 20646 3495 20698
rect 3507 20646 3559 20698
rect 7982 20646 8034 20698
rect 8046 20646 8098 20698
rect 8110 20646 8162 20698
rect 8174 20646 8226 20698
rect 5648 20102 5700 20154
rect 5712 20102 5764 20154
rect 5776 20102 5828 20154
rect 5840 20102 5892 20154
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 3315 19558 3367 19610
rect 3379 19558 3431 19610
rect 3443 19558 3495 19610
rect 3507 19558 3559 19610
rect 7982 19558 8034 19610
rect 8046 19558 8098 19610
rect 8110 19558 8162 19610
rect 8174 19558 8226 19610
rect 11244 19499 11296 19508
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 10048 19252 10100 19304
rect 10784 19116 10836 19168
rect 5648 19014 5700 19066
rect 5712 19014 5764 19066
rect 5776 19014 5828 19066
rect 5840 19014 5892 19066
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 11612 18955 11664 18964
rect 11612 18921 11621 18955
rect 11621 18921 11655 18955
rect 11655 18921 11664 18955
rect 11612 18912 11664 18921
rect 10784 18844 10836 18896
rect 8760 18708 8812 18760
rect 11796 18708 11848 18760
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 10048 18572 10100 18624
rect 3315 18470 3367 18522
rect 3379 18470 3431 18522
rect 3443 18470 3495 18522
rect 3507 18470 3559 18522
rect 7982 18470 8034 18522
rect 8046 18470 8098 18522
rect 8110 18470 8162 18522
rect 8174 18470 8226 18522
rect 9404 18411 9456 18420
rect 9404 18377 9413 18411
rect 9413 18377 9447 18411
rect 9447 18377 9456 18411
rect 9404 18368 9456 18377
rect 11152 18411 11204 18420
rect 11152 18377 11161 18411
rect 11161 18377 11195 18411
rect 11195 18377 11204 18411
rect 11152 18368 11204 18377
rect 11796 18411 11848 18420
rect 11796 18377 11805 18411
rect 11805 18377 11839 18411
rect 11839 18377 11848 18411
rect 11796 18368 11848 18377
rect 8576 18164 8628 18216
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 10784 18028 10836 18080
rect 5648 17926 5700 17978
rect 5712 17926 5764 17978
rect 5776 17926 5828 17978
rect 5840 17926 5892 17978
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 10784 17756 10836 17808
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 8668 17527 8720 17536
rect 8668 17493 8677 17527
rect 8677 17493 8711 17527
rect 8711 17493 8720 17527
rect 8668 17484 8720 17493
rect 3315 17382 3367 17434
rect 3379 17382 3431 17434
rect 3443 17382 3495 17434
rect 3507 17382 3559 17434
rect 7982 17382 8034 17434
rect 8046 17382 8098 17434
rect 8110 17382 8162 17434
rect 8174 17382 8226 17434
rect 10140 17280 10192 17332
rect 10692 17212 10744 17264
rect 8484 17076 8536 17128
rect 9772 17076 9824 17128
rect 9864 17119 9916 17128
rect 9864 17085 9873 17119
rect 9873 17085 9907 17119
rect 9907 17085 9916 17119
rect 11244 17119 11296 17128
rect 9864 17076 9916 17085
rect 11244 17085 11253 17119
rect 11253 17085 11287 17119
rect 11287 17085 11296 17119
rect 11796 17119 11848 17128
rect 11244 17076 11296 17085
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 8300 16940 8352 16992
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 8576 16940 8628 16992
rect 10784 16940 10836 16992
rect 5648 16838 5700 16890
rect 5712 16838 5764 16890
rect 5776 16838 5828 16890
rect 5840 16838 5892 16890
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 9956 16736 10008 16788
rect 10784 16668 10836 16720
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 8576 16464 8628 16516
rect 9956 16464 10008 16516
rect 8944 16396 8996 16448
rect 3315 16294 3367 16346
rect 3379 16294 3431 16346
rect 3443 16294 3495 16346
rect 3507 16294 3559 16346
rect 7982 16294 8034 16346
rect 8046 16294 8098 16346
rect 8110 16294 8162 16346
rect 8174 16294 8226 16346
rect 10692 16192 10744 16244
rect 11244 16192 11296 16244
rect 10048 16124 10100 16176
rect 8300 16056 8352 16108
rect 7840 15920 7892 15972
rect 9036 15988 9088 16040
rect 9772 16031 9824 16040
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 9956 15988 10008 16040
rect 8944 15852 8996 15904
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 5648 15750 5700 15802
rect 5712 15750 5764 15802
rect 5776 15750 5828 15802
rect 5840 15750 5892 15802
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 9956 15691 10008 15700
rect 7380 15580 7432 15632
rect 8576 15580 8628 15632
rect 8760 15623 8812 15632
rect 8760 15589 8769 15623
rect 8769 15589 8803 15623
rect 8803 15589 8812 15623
rect 8760 15580 8812 15589
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 10140 15580 10192 15632
rect 7840 15444 7892 15496
rect 8944 15308 8996 15360
rect 9772 15444 9824 15496
rect 10692 15512 10744 15564
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 3315 15206 3367 15258
rect 3379 15206 3431 15258
rect 3443 15206 3495 15258
rect 3507 15206 3559 15258
rect 7982 15206 8034 15258
rect 8046 15206 8098 15258
rect 8110 15206 8162 15258
rect 8174 15206 8226 15258
rect 7380 15147 7432 15156
rect 7380 15113 7389 15147
rect 7389 15113 7423 15147
rect 7423 15113 7432 15147
rect 7380 15104 7432 15113
rect 8300 15104 8352 15156
rect 9220 15104 9272 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 9312 14968 9364 15020
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 11244 15011 11296 15020
rect 11244 14977 11253 15011
rect 11253 14977 11287 15011
rect 11287 14977 11296 15011
rect 11244 14968 11296 14977
rect 9772 14900 9824 14952
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 7840 14832 7892 14884
rect 8944 14875 8996 14884
rect 8944 14841 8953 14875
rect 8953 14841 8987 14875
rect 8987 14841 8996 14875
rect 8944 14832 8996 14841
rect 9312 14875 9364 14884
rect 9312 14841 9321 14875
rect 9321 14841 9355 14875
rect 9355 14841 9364 14875
rect 9312 14832 9364 14841
rect 9588 14832 9640 14884
rect 10876 14875 10928 14884
rect 10876 14841 10885 14875
rect 10885 14841 10919 14875
rect 10919 14841 10928 14875
rect 10876 14832 10928 14841
rect 8760 14764 8812 14816
rect 9404 14764 9456 14816
rect 9956 14764 10008 14816
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 5648 14662 5700 14714
rect 5712 14662 5764 14714
rect 5776 14662 5828 14714
rect 5840 14662 5892 14714
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 9312 14560 9364 14612
rect 9220 14492 9272 14544
rect 10784 14492 10836 14544
rect 7840 14424 7892 14476
rect 8484 14424 8536 14476
rect 9312 14424 9364 14476
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 8760 14399 8812 14408
rect 8760 14365 8769 14399
rect 8769 14365 8803 14399
rect 8803 14365 8812 14399
rect 8760 14356 8812 14365
rect 8576 14288 8628 14340
rect 10876 14356 10928 14408
rect 3315 14118 3367 14170
rect 3379 14118 3431 14170
rect 3443 14118 3495 14170
rect 3507 14118 3559 14170
rect 7982 14118 8034 14170
rect 8046 14118 8098 14170
rect 8110 14118 8162 14170
rect 8174 14118 8226 14170
rect 8944 13812 8996 13864
rect 9404 13812 9456 13864
rect 10048 13812 10100 13864
rect 7840 13676 7892 13728
rect 8760 13676 8812 13728
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 5648 13574 5700 13626
rect 5712 13574 5764 13626
rect 5776 13574 5828 13626
rect 5840 13574 5892 13626
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 11796 13515 11848 13524
rect 11796 13481 11805 13515
rect 11805 13481 11839 13515
rect 11839 13481 11848 13515
rect 11796 13472 11848 13481
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 11244 13268 11296 13320
rect 3315 13030 3367 13082
rect 3379 13030 3431 13082
rect 3443 13030 3495 13082
rect 3507 13030 3559 13082
rect 7982 13030 8034 13082
rect 8046 13030 8098 13082
rect 8110 13030 8162 13082
rect 8174 13030 8226 13082
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 1308 12588 1360 12640
rect 9588 12724 9640 12776
rect 9036 12656 9088 12708
rect 11244 12588 11296 12640
rect 5648 12486 5700 12538
rect 5712 12486 5764 12538
rect 5776 12486 5828 12538
rect 5840 12486 5892 12538
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 8760 12087 8812 12096
rect 8760 12053 8769 12087
rect 8769 12053 8803 12087
rect 8803 12053 8812 12087
rect 8760 12044 8812 12053
rect 3315 11942 3367 11994
rect 3379 11942 3431 11994
rect 3443 11942 3495 11994
rect 3507 11942 3559 11994
rect 7982 11942 8034 11994
rect 8046 11942 8098 11994
rect 8110 11942 8162 11994
rect 8174 11942 8226 11994
rect 9772 11704 9824 11756
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 9036 11636 9088 11688
rect 9404 11636 9456 11688
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 5648 11398 5700 11450
rect 5712 11398 5764 11450
rect 5776 11398 5828 11450
rect 5840 11398 5892 11450
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 10692 11339 10744 11348
rect 10692 11305 10701 11339
rect 10701 11305 10735 11339
rect 10735 11305 10744 11339
rect 10692 11296 10744 11305
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 10140 11160 10192 11212
rect 9404 10956 9456 11008
rect 3315 10854 3367 10906
rect 3379 10854 3431 10906
rect 3443 10854 3495 10906
rect 3507 10854 3559 10906
rect 7982 10854 8034 10906
rect 8046 10854 8098 10906
rect 8110 10854 8162 10906
rect 8174 10854 8226 10906
rect 10140 10752 10192 10804
rect 9496 10412 9548 10464
rect 10692 10412 10744 10464
rect 5648 10310 5700 10362
rect 5712 10310 5764 10362
rect 5776 10310 5828 10362
rect 5840 10310 5892 10362
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 3315 9766 3367 9818
rect 3379 9766 3431 9818
rect 3443 9766 3495 9818
rect 3507 9766 3559 9818
rect 7982 9766 8034 9818
rect 8046 9766 8098 9818
rect 8110 9766 8162 9818
rect 8174 9766 8226 9818
rect 5648 9222 5700 9274
rect 5712 9222 5764 9274
rect 5776 9222 5828 9274
rect 5840 9222 5892 9274
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 3315 8678 3367 8730
rect 3379 8678 3431 8730
rect 3443 8678 3495 8730
rect 3507 8678 3559 8730
rect 7982 8678 8034 8730
rect 8046 8678 8098 8730
rect 8110 8678 8162 8730
rect 8174 8678 8226 8730
rect 5648 8134 5700 8186
rect 5712 8134 5764 8186
rect 5776 8134 5828 8186
rect 5840 8134 5892 8186
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 3315 7590 3367 7642
rect 3379 7590 3431 7642
rect 3443 7590 3495 7642
rect 3507 7590 3559 7642
rect 7982 7590 8034 7642
rect 8046 7590 8098 7642
rect 8110 7590 8162 7642
rect 8174 7590 8226 7642
rect 5648 7046 5700 7098
rect 5712 7046 5764 7098
rect 5776 7046 5828 7098
rect 5840 7046 5892 7098
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 3315 6502 3367 6554
rect 3379 6502 3431 6554
rect 3443 6502 3495 6554
rect 3507 6502 3559 6554
rect 7982 6502 8034 6554
rect 8046 6502 8098 6554
rect 8110 6502 8162 6554
rect 8174 6502 8226 6554
rect 5648 5958 5700 6010
rect 5712 5958 5764 6010
rect 5776 5958 5828 6010
rect 5840 5958 5892 6010
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 3315 5414 3367 5466
rect 3379 5414 3431 5466
rect 3443 5414 3495 5466
rect 3507 5414 3559 5466
rect 7982 5414 8034 5466
rect 8046 5414 8098 5466
rect 8110 5414 8162 5466
rect 8174 5414 8226 5466
rect 5648 4870 5700 4922
rect 5712 4870 5764 4922
rect 5776 4870 5828 4922
rect 5840 4870 5892 4922
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 3315 4326 3367 4378
rect 3379 4326 3431 4378
rect 3443 4326 3495 4378
rect 3507 4326 3559 4378
rect 7982 4326 8034 4378
rect 8046 4326 8098 4378
rect 8110 4326 8162 4378
rect 8174 4326 8226 4378
rect 11428 4267 11480 4276
rect 11428 4233 11437 4267
rect 11437 4233 11471 4267
rect 11471 4233 11480 4267
rect 11428 4224 11480 4233
rect 9404 4199 9456 4208
rect 9404 4165 9413 4199
rect 9413 4165 9447 4199
rect 9447 4165 9456 4199
rect 9404 4156 9456 4165
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 11244 4063 11296 4072
rect 9220 4020 9272 4029
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 10048 3884 10100 3936
rect 11704 3884 11756 3936
rect 5648 3782 5700 3834
rect 5712 3782 5764 3834
rect 5776 3782 5828 3834
rect 5840 3782 5892 3834
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 9404 3680 9456 3732
rect 9496 3680 9548 3732
rect 10692 3680 10744 3732
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 11244 3340 11296 3392
rect 3315 3238 3367 3290
rect 3379 3238 3431 3290
rect 3443 3238 3495 3290
rect 3507 3238 3559 3290
rect 7982 3238 8034 3290
rect 8046 3238 8098 3290
rect 8110 3238 8162 3290
rect 8174 3238 8226 3290
rect 10140 3000 10192 3052
rect 9036 2975 9088 2984
rect 6000 2796 6052 2848
rect 7840 2796 7892 2848
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 10692 2796 10744 2848
rect 12348 2796 12400 2848
rect 5648 2694 5700 2746
rect 5712 2694 5764 2746
rect 5776 2694 5828 2746
rect 5840 2694 5892 2746
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 10968 2635 11020 2644
rect 10968 2601 10977 2635
rect 10977 2601 11011 2635
rect 11011 2601 11020 2635
rect 10968 2592 11020 2601
rect 11704 2635 11756 2644
rect 11704 2601 11713 2635
rect 11713 2601 11747 2635
rect 11747 2601 11756 2635
rect 11704 2592 11756 2601
rect 11244 2499 11296 2508
rect 11244 2465 11253 2499
rect 11253 2465 11287 2499
rect 11287 2465 11296 2499
rect 11244 2456 11296 2465
rect 10968 2388 11020 2440
rect 8392 2252 8444 2304
rect 9772 2252 9824 2304
rect 3315 2150 3367 2202
rect 3379 2150 3431 2202
rect 3443 2150 3495 2202
rect 3507 2150 3559 2202
rect 7982 2150 8034 2202
rect 8046 2150 8098 2202
rect 8110 2150 8162 2202
rect 8174 2150 8226 2202
<< metal2 >>
rect 3289 106652 3585 106672
rect 3345 106650 3369 106652
rect 3425 106650 3449 106652
rect 3505 106650 3529 106652
rect 3367 106598 3369 106650
rect 3431 106598 3443 106650
rect 3505 106598 3507 106650
rect 3345 106596 3369 106598
rect 3425 106596 3449 106598
rect 3505 106596 3529 106598
rect 3289 106576 3585 106596
rect 7956 106652 8252 106672
rect 8012 106650 8036 106652
rect 8092 106650 8116 106652
rect 8172 106650 8196 106652
rect 8034 106598 8036 106650
rect 8098 106598 8110 106650
rect 8172 106598 8174 106650
rect 8012 106596 8036 106598
rect 8092 106596 8116 106598
rect 8172 106596 8196 106598
rect 7956 106576 8252 106596
rect 5622 106108 5918 106128
rect 5678 106106 5702 106108
rect 5758 106106 5782 106108
rect 5838 106106 5862 106108
rect 5700 106054 5702 106106
rect 5764 106054 5776 106106
rect 5838 106054 5840 106106
rect 5678 106052 5702 106054
rect 5758 106052 5782 106054
rect 5838 106052 5862 106054
rect 5622 106032 5918 106052
rect 10289 106108 10585 106128
rect 10345 106106 10369 106108
rect 10425 106106 10449 106108
rect 10505 106106 10529 106108
rect 10367 106054 10369 106106
rect 10431 106054 10443 106106
rect 10505 106054 10507 106106
rect 10345 106052 10369 106054
rect 10425 106052 10449 106054
rect 10505 106052 10529 106054
rect 10289 106032 10585 106052
rect 3289 105564 3585 105584
rect 3345 105562 3369 105564
rect 3425 105562 3449 105564
rect 3505 105562 3529 105564
rect 3367 105510 3369 105562
rect 3431 105510 3443 105562
rect 3505 105510 3507 105562
rect 3345 105508 3369 105510
rect 3425 105508 3449 105510
rect 3505 105508 3529 105510
rect 3289 105488 3585 105508
rect 7956 105564 8252 105584
rect 8012 105562 8036 105564
rect 8092 105562 8116 105564
rect 8172 105562 8196 105564
rect 8034 105510 8036 105562
rect 8098 105510 8110 105562
rect 8172 105510 8174 105562
rect 8012 105508 8036 105510
rect 8092 105508 8116 105510
rect 8172 105508 8196 105510
rect 7956 105488 8252 105508
rect 11426 105496 11482 105505
rect 11426 105431 11482 105440
rect 5622 105020 5918 105040
rect 5678 105018 5702 105020
rect 5758 105018 5782 105020
rect 5838 105018 5862 105020
rect 5700 104966 5702 105018
rect 5764 104966 5776 105018
rect 5838 104966 5840 105018
rect 5678 104964 5702 104966
rect 5758 104964 5782 104966
rect 5838 104964 5862 104966
rect 5622 104944 5918 104964
rect 10289 105020 10585 105040
rect 10345 105018 10369 105020
rect 10425 105018 10449 105020
rect 10505 105018 10529 105020
rect 10367 104966 10369 105018
rect 10431 104966 10443 105018
rect 10505 104966 10507 105018
rect 10345 104964 10369 104966
rect 10425 104964 10449 104966
rect 10505 104964 10529 104966
rect 10289 104944 10585 104964
rect 3289 104476 3585 104496
rect 3345 104474 3369 104476
rect 3425 104474 3449 104476
rect 3505 104474 3529 104476
rect 3367 104422 3369 104474
rect 3431 104422 3443 104474
rect 3505 104422 3507 104474
rect 3345 104420 3369 104422
rect 3425 104420 3449 104422
rect 3505 104420 3529 104422
rect 3289 104400 3585 104420
rect 7956 104476 8252 104496
rect 8012 104474 8036 104476
rect 8092 104474 8116 104476
rect 8172 104474 8196 104476
rect 8034 104422 8036 104474
rect 8098 104422 8110 104474
rect 8172 104422 8174 104474
rect 8012 104420 8036 104422
rect 8092 104420 8116 104422
rect 8172 104420 8196 104422
rect 7956 104400 8252 104420
rect 5622 103932 5918 103952
rect 5678 103930 5702 103932
rect 5758 103930 5782 103932
rect 5838 103930 5862 103932
rect 5700 103878 5702 103930
rect 5764 103878 5776 103930
rect 5838 103878 5840 103930
rect 5678 103876 5702 103878
rect 5758 103876 5782 103878
rect 5838 103876 5862 103878
rect 5622 103856 5918 103876
rect 10289 103932 10585 103952
rect 10345 103930 10369 103932
rect 10425 103930 10449 103932
rect 10505 103930 10529 103932
rect 10367 103878 10369 103930
rect 10431 103878 10443 103930
rect 10505 103878 10507 103930
rect 10345 103876 10369 103878
rect 10425 103876 10449 103878
rect 10505 103876 10529 103878
rect 10289 103856 10585 103876
rect 3289 103388 3585 103408
rect 3345 103386 3369 103388
rect 3425 103386 3449 103388
rect 3505 103386 3529 103388
rect 3367 103334 3369 103386
rect 3431 103334 3443 103386
rect 3505 103334 3507 103386
rect 3345 103332 3369 103334
rect 3425 103332 3449 103334
rect 3505 103332 3529 103334
rect 3289 103312 3585 103332
rect 7956 103388 8252 103408
rect 8012 103386 8036 103388
rect 8092 103386 8116 103388
rect 8172 103386 8196 103388
rect 8034 103334 8036 103386
rect 8098 103334 8110 103386
rect 8172 103334 8174 103386
rect 8012 103332 8036 103334
rect 8092 103332 8116 103334
rect 8172 103332 8196 103334
rect 7956 103312 8252 103332
rect 5622 102844 5918 102864
rect 5678 102842 5702 102844
rect 5758 102842 5782 102844
rect 5838 102842 5862 102844
rect 5700 102790 5702 102842
rect 5764 102790 5776 102842
rect 5838 102790 5840 102842
rect 5678 102788 5702 102790
rect 5758 102788 5782 102790
rect 5838 102788 5862 102790
rect 5622 102768 5918 102788
rect 10289 102844 10585 102864
rect 10345 102842 10369 102844
rect 10425 102842 10449 102844
rect 10505 102842 10529 102844
rect 10367 102790 10369 102842
rect 10431 102790 10443 102842
rect 10505 102790 10507 102842
rect 10345 102788 10369 102790
rect 10425 102788 10449 102790
rect 10505 102788 10529 102790
rect 10289 102768 10585 102788
rect 3289 102300 3585 102320
rect 3345 102298 3369 102300
rect 3425 102298 3449 102300
rect 3505 102298 3529 102300
rect 3367 102246 3369 102298
rect 3431 102246 3443 102298
rect 3505 102246 3507 102298
rect 3345 102244 3369 102246
rect 3425 102244 3449 102246
rect 3505 102244 3529 102246
rect 3289 102224 3585 102244
rect 7956 102300 8252 102320
rect 8012 102298 8036 102300
rect 8092 102298 8116 102300
rect 8172 102298 8196 102300
rect 8034 102246 8036 102298
rect 8098 102246 8110 102298
rect 8172 102246 8174 102298
rect 8012 102244 8036 102246
rect 8092 102244 8116 102246
rect 8172 102244 8196 102246
rect 7956 102224 8252 102244
rect 110 102096 166 102105
rect 110 102031 166 102040
rect 124 97209 152 102031
rect 5622 101756 5918 101776
rect 5678 101754 5702 101756
rect 5758 101754 5782 101756
rect 5838 101754 5862 101756
rect 5700 101702 5702 101754
rect 5764 101702 5776 101754
rect 5838 101702 5840 101754
rect 5678 101700 5702 101702
rect 5758 101700 5782 101702
rect 5838 101700 5862 101702
rect 5622 101680 5918 101700
rect 10289 101756 10585 101776
rect 10345 101754 10369 101756
rect 10425 101754 10449 101756
rect 10505 101754 10529 101756
rect 10367 101702 10369 101754
rect 10431 101702 10443 101754
rect 10505 101702 10507 101754
rect 10345 101700 10369 101702
rect 10425 101700 10449 101702
rect 10505 101700 10529 101702
rect 10289 101680 10585 101700
rect 3289 101212 3585 101232
rect 3345 101210 3369 101212
rect 3425 101210 3449 101212
rect 3505 101210 3529 101212
rect 3367 101158 3369 101210
rect 3431 101158 3443 101210
rect 3505 101158 3507 101210
rect 3345 101156 3369 101158
rect 3425 101156 3449 101158
rect 3505 101156 3529 101158
rect 3289 101136 3585 101156
rect 7956 101212 8252 101232
rect 8012 101210 8036 101212
rect 8092 101210 8116 101212
rect 8172 101210 8196 101212
rect 8034 101158 8036 101210
rect 8098 101158 8110 101210
rect 8172 101158 8174 101210
rect 8012 101156 8036 101158
rect 8092 101156 8116 101158
rect 8172 101156 8196 101158
rect 7956 101136 8252 101156
rect 5622 100668 5918 100688
rect 5678 100666 5702 100668
rect 5758 100666 5782 100668
rect 5838 100666 5862 100668
rect 5700 100614 5702 100666
rect 5764 100614 5776 100666
rect 5838 100614 5840 100666
rect 5678 100612 5702 100614
rect 5758 100612 5782 100614
rect 5838 100612 5862 100614
rect 5622 100592 5918 100612
rect 10289 100668 10585 100688
rect 10345 100666 10369 100668
rect 10425 100666 10449 100668
rect 10505 100666 10529 100668
rect 10367 100614 10369 100666
rect 10431 100614 10443 100666
rect 10505 100614 10507 100666
rect 10345 100612 10369 100614
rect 10425 100612 10449 100614
rect 10505 100612 10529 100614
rect 10289 100592 10585 100612
rect 3289 100124 3585 100144
rect 3345 100122 3369 100124
rect 3425 100122 3449 100124
rect 3505 100122 3529 100124
rect 3367 100070 3369 100122
rect 3431 100070 3443 100122
rect 3505 100070 3507 100122
rect 3345 100068 3369 100070
rect 3425 100068 3449 100070
rect 3505 100068 3529 100070
rect 3289 100048 3585 100068
rect 7956 100124 8252 100144
rect 8012 100122 8036 100124
rect 8092 100122 8116 100124
rect 8172 100122 8196 100124
rect 8034 100070 8036 100122
rect 8098 100070 8110 100122
rect 8172 100070 8174 100122
rect 8012 100068 8036 100070
rect 8092 100068 8116 100070
rect 8172 100068 8196 100070
rect 7956 100048 8252 100068
rect 5622 99580 5918 99600
rect 5678 99578 5702 99580
rect 5758 99578 5782 99580
rect 5838 99578 5862 99580
rect 5700 99526 5702 99578
rect 5764 99526 5776 99578
rect 5838 99526 5840 99578
rect 5678 99524 5702 99526
rect 5758 99524 5782 99526
rect 5838 99524 5862 99526
rect 5622 99504 5918 99524
rect 10289 99580 10585 99600
rect 10345 99578 10369 99580
rect 10425 99578 10449 99580
rect 10505 99578 10529 99580
rect 10367 99526 10369 99578
rect 10431 99526 10443 99578
rect 10505 99526 10507 99578
rect 10345 99524 10369 99526
rect 10425 99524 10449 99526
rect 10505 99524 10529 99526
rect 10289 99504 10585 99524
rect 3289 99036 3585 99056
rect 3345 99034 3369 99036
rect 3425 99034 3449 99036
rect 3505 99034 3529 99036
rect 3367 98982 3369 99034
rect 3431 98982 3443 99034
rect 3505 98982 3507 99034
rect 3345 98980 3369 98982
rect 3425 98980 3449 98982
rect 3505 98980 3529 98982
rect 3289 98960 3585 98980
rect 7956 99036 8252 99056
rect 8012 99034 8036 99036
rect 8092 99034 8116 99036
rect 8172 99034 8196 99036
rect 8034 98982 8036 99034
rect 8098 98982 8110 99034
rect 8172 98982 8174 99034
rect 8012 98980 8036 98982
rect 8092 98980 8116 98982
rect 8172 98980 8196 98982
rect 7956 98960 8252 98980
rect 11150 98696 11206 98705
rect 11150 98631 11206 98640
rect 5622 98492 5918 98512
rect 5678 98490 5702 98492
rect 5758 98490 5782 98492
rect 5838 98490 5862 98492
rect 5700 98438 5702 98490
rect 5764 98438 5776 98490
rect 5838 98438 5840 98490
rect 5678 98436 5702 98438
rect 5758 98436 5782 98438
rect 5838 98436 5862 98438
rect 5622 98416 5918 98436
rect 10289 98492 10585 98512
rect 10345 98490 10369 98492
rect 10425 98490 10449 98492
rect 10505 98490 10529 98492
rect 10367 98438 10369 98490
rect 10431 98438 10443 98490
rect 10505 98438 10507 98490
rect 10345 98436 10369 98438
rect 10425 98436 10449 98438
rect 10505 98436 10529 98438
rect 10289 98416 10585 98436
rect 3289 97948 3585 97968
rect 3345 97946 3369 97948
rect 3425 97946 3449 97948
rect 3505 97946 3529 97948
rect 3367 97894 3369 97946
rect 3431 97894 3443 97946
rect 3505 97894 3507 97946
rect 3345 97892 3369 97894
rect 3425 97892 3449 97894
rect 3505 97892 3529 97894
rect 3289 97872 3585 97892
rect 7956 97948 8252 97968
rect 8012 97946 8036 97948
rect 8092 97946 8116 97948
rect 8172 97946 8196 97948
rect 8034 97894 8036 97946
rect 8098 97894 8110 97946
rect 8172 97894 8174 97946
rect 8012 97892 8036 97894
rect 8092 97892 8116 97894
rect 8172 97892 8196 97894
rect 7956 97872 8252 97892
rect 5622 97404 5918 97424
rect 5678 97402 5702 97404
rect 5758 97402 5782 97404
rect 5838 97402 5862 97404
rect 5700 97350 5702 97402
rect 5764 97350 5776 97402
rect 5838 97350 5840 97402
rect 5678 97348 5702 97350
rect 5758 97348 5782 97350
rect 5838 97348 5862 97350
rect 5622 97328 5918 97348
rect 10289 97404 10585 97424
rect 10345 97402 10369 97404
rect 10425 97402 10449 97404
rect 10505 97402 10529 97404
rect 10367 97350 10369 97402
rect 10431 97350 10443 97402
rect 10505 97350 10507 97402
rect 10345 97348 10369 97350
rect 10425 97348 10449 97350
rect 10505 97348 10529 97350
rect 10289 97328 10585 97348
rect 110 97200 166 97209
rect 110 97135 166 97144
rect 3289 96860 3585 96880
rect 3345 96858 3369 96860
rect 3425 96858 3449 96860
rect 3505 96858 3529 96860
rect 3367 96806 3369 96858
rect 3431 96806 3443 96858
rect 3505 96806 3507 96858
rect 3345 96804 3369 96806
rect 3425 96804 3449 96806
rect 3505 96804 3529 96806
rect 3289 96784 3585 96804
rect 7956 96860 8252 96880
rect 8012 96858 8036 96860
rect 8092 96858 8116 96860
rect 8172 96858 8196 96860
rect 8034 96806 8036 96858
rect 8098 96806 8110 96858
rect 8172 96806 8174 96858
rect 8012 96804 8036 96806
rect 8092 96804 8116 96806
rect 8172 96804 8196 96806
rect 7956 96784 8252 96804
rect 5622 96316 5918 96336
rect 5678 96314 5702 96316
rect 5758 96314 5782 96316
rect 5838 96314 5862 96316
rect 5700 96262 5702 96314
rect 5764 96262 5776 96314
rect 5838 96262 5840 96314
rect 5678 96260 5702 96262
rect 5758 96260 5782 96262
rect 5838 96260 5862 96262
rect 5622 96240 5918 96260
rect 10289 96316 10585 96336
rect 10345 96314 10369 96316
rect 10425 96314 10449 96316
rect 10505 96314 10529 96316
rect 10367 96262 10369 96314
rect 10431 96262 10443 96314
rect 10505 96262 10507 96314
rect 10345 96260 10369 96262
rect 10425 96260 10449 96262
rect 10505 96260 10529 96262
rect 10289 96240 10585 96260
rect 3289 95772 3585 95792
rect 3345 95770 3369 95772
rect 3425 95770 3449 95772
rect 3505 95770 3529 95772
rect 3367 95718 3369 95770
rect 3431 95718 3443 95770
rect 3505 95718 3507 95770
rect 3345 95716 3369 95718
rect 3425 95716 3449 95718
rect 3505 95716 3529 95718
rect 3289 95696 3585 95716
rect 7956 95772 8252 95792
rect 8012 95770 8036 95772
rect 8092 95770 8116 95772
rect 8172 95770 8196 95772
rect 8034 95718 8036 95770
rect 8098 95718 8110 95770
rect 8172 95718 8174 95770
rect 8012 95716 8036 95718
rect 8092 95716 8116 95718
rect 8172 95716 8196 95718
rect 7956 95696 8252 95716
rect 5622 95228 5918 95248
rect 5678 95226 5702 95228
rect 5758 95226 5782 95228
rect 5838 95226 5862 95228
rect 5700 95174 5702 95226
rect 5764 95174 5776 95226
rect 5838 95174 5840 95226
rect 5678 95172 5702 95174
rect 5758 95172 5782 95174
rect 5838 95172 5862 95174
rect 5622 95152 5918 95172
rect 10289 95228 10585 95248
rect 10345 95226 10369 95228
rect 10425 95226 10449 95228
rect 10505 95226 10529 95228
rect 10367 95174 10369 95226
rect 10431 95174 10443 95226
rect 10505 95174 10507 95226
rect 10345 95172 10369 95174
rect 10425 95172 10449 95174
rect 10505 95172 10529 95174
rect 10289 95152 10585 95172
rect 11060 94988 11112 94994
rect 11060 94930 11112 94936
rect 3289 94684 3585 94704
rect 3345 94682 3369 94684
rect 3425 94682 3449 94684
rect 3505 94682 3529 94684
rect 3367 94630 3369 94682
rect 3431 94630 3443 94682
rect 3505 94630 3507 94682
rect 3345 94628 3369 94630
rect 3425 94628 3449 94630
rect 3505 94628 3529 94630
rect 3289 94608 3585 94628
rect 7956 94684 8252 94704
rect 8012 94682 8036 94684
rect 8092 94682 8116 94684
rect 8172 94682 8196 94684
rect 8034 94630 8036 94682
rect 8098 94630 8110 94682
rect 8172 94630 8174 94682
rect 8012 94628 8036 94630
rect 8092 94628 8116 94630
rect 8172 94628 8196 94630
rect 7956 94608 8252 94628
rect 11072 94314 11100 94930
rect 11164 94926 11192 98631
rect 11440 97850 11468 105431
rect 11428 97844 11480 97850
rect 11428 97786 11480 97792
rect 11244 97640 11296 97646
rect 11244 97582 11296 97588
rect 11256 97209 11284 97582
rect 11242 97200 11298 97209
rect 11242 97135 11298 97144
rect 11152 94920 11204 94926
rect 11152 94862 11204 94868
rect 11164 94586 11192 94862
rect 11256 94858 11284 97135
rect 11244 94852 11296 94858
rect 11244 94794 11296 94800
rect 11152 94580 11204 94586
rect 11152 94522 11204 94528
rect 11060 94308 11112 94314
rect 11060 94250 11112 94256
rect 5622 94140 5918 94160
rect 5678 94138 5702 94140
rect 5758 94138 5782 94140
rect 5838 94138 5862 94140
rect 5700 94086 5702 94138
rect 5764 94086 5776 94138
rect 5838 94086 5840 94138
rect 5678 94084 5702 94086
rect 5758 94084 5782 94086
rect 5838 94084 5862 94086
rect 5622 94064 5918 94084
rect 10289 94140 10585 94160
rect 10345 94138 10369 94140
rect 10425 94138 10449 94140
rect 10505 94138 10529 94140
rect 10367 94086 10369 94138
rect 10431 94086 10443 94138
rect 10505 94086 10507 94138
rect 10345 94084 10369 94086
rect 10425 94084 10449 94086
rect 10505 94084 10529 94086
rect 10289 94064 10585 94084
rect 3289 93596 3585 93616
rect 3345 93594 3369 93596
rect 3425 93594 3449 93596
rect 3505 93594 3529 93596
rect 3367 93542 3369 93594
rect 3431 93542 3443 93594
rect 3505 93542 3507 93594
rect 3345 93540 3369 93542
rect 3425 93540 3449 93542
rect 3505 93540 3529 93542
rect 3289 93520 3585 93540
rect 7956 93596 8252 93616
rect 8012 93594 8036 93596
rect 8092 93594 8116 93596
rect 8172 93594 8196 93596
rect 8034 93542 8036 93594
rect 8098 93542 8110 93594
rect 8172 93542 8174 93594
rect 8012 93540 8036 93542
rect 8092 93540 8116 93542
rect 8172 93540 8196 93542
rect 7956 93520 8252 93540
rect 5622 93052 5918 93072
rect 5678 93050 5702 93052
rect 5758 93050 5782 93052
rect 5838 93050 5862 93052
rect 5700 92998 5702 93050
rect 5764 92998 5776 93050
rect 5838 92998 5840 93050
rect 5678 92996 5702 92998
rect 5758 92996 5782 92998
rect 5838 92996 5862 92998
rect 5622 92976 5918 92996
rect 10289 93052 10585 93072
rect 10345 93050 10369 93052
rect 10425 93050 10449 93052
rect 10505 93050 10529 93052
rect 10367 92998 10369 93050
rect 10431 92998 10443 93050
rect 10505 92998 10507 93050
rect 10345 92996 10369 92998
rect 10425 92996 10449 92998
rect 10505 92996 10529 92998
rect 10289 92976 10585 92996
rect 3289 92508 3585 92528
rect 3345 92506 3369 92508
rect 3425 92506 3449 92508
rect 3505 92506 3529 92508
rect 3367 92454 3369 92506
rect 3431 92454 3443 92506
rect 3505 92454 3507 92506
rect 3345 92452 3369 92454
rect 3425 92452 3449 92454
rect 3505 92452 3529 92454
rect 3289 92432 3585 92452
rect 7956 92508 8252 92528
rect 8012 92506 8036 92508
rect 8092 92506 8116 92508
rect 8172 92506 8196 92508
rect 8034 92454 8036 92506
rect 8098 92454 8110 92506
rect 8172 92454 8174 92506
rect 8012 92452 8036 92454
rect 8092 92452 8116 92454
rect 8172 92452 8196 92454
rect 7956 92432 8252 92452
rect 5622 91964 5918 91984
rect 5678 91962 5702 91964
rect 5758 91962 5782 91964
rect 5838 91962 5862 91964
rect 5700 91910 5702 91962
rect 5764 91910 5776 91962
rect 5838 91910 5840 91962
rect 5678 91908 5702 91910
rect 5758 91908 5782 91910
rect 5838 91908 5862 91910
rect 5622 91888 5918 91908
rect 10289 91964 10585 91984
rect 10345 91962 10369 91964
rect 10425 91962 10449 91964
rect 10505 91962 10529 91964
rect 10367 91910 10369 91962
rect 10431 91910 10443 91962
rect 10505 91910 10507 91962
rect 10345 91908 10369 91910
rect 10425 91908 10449 91910
rect 10505 91908 10529 91910
rect 10289 91888 10585 91908
rect 10690 91896 10746 91905
rect 10690 91831 10746 91840
rect 3289 91420 3585 91440
rect 3345 91418 3369 91420
rect 3425 91418 3449 91420
rect 3505 91418 3529 91420
rect 3367 91366 3369 91418
rect 3431 91366 3443 91418
rect 3505 91366 3507 91418
rect 3345 91364 3369 91366
rect 3425 91364 3449 91366
rect 3505 91364 3529 91366
rect 3289 91344 3585 91364
rect 7956 91420 8252 91440
rect 8012 91418 8036 91420
rect 8092 91418 8116 91420
rect 8172 91418 8196 91420
rect 8034 91366 8036 91418
rect 8098 91366 8110 91418
rect 8172 91366 8174 91418
rect 8012 91364 8036 91366
rect 8092 91364 8116 91366
rect 8172 91364 8196 91366
rect 7956 91344 8252 91364
rect 5622 90876 5918 90896
rect 5678 90874 5702 90876
rect 5758 90874 5782 90876
rect 5838 90874 5862 90876
rect 5700 90822 5702 90874
rect 5764 90822 5776 90874
rect 5838 90822 5840 90874
rect 5678 90820 5702 90822
rect 5758 90820 5782 90822
rect 5838 90820 5862 90822
rect 5622 90800 5918 90820
rect 10289 90876 10585 90896
rect 10345 90874 10369 90876
rect 10425 90874 10449 90876
rect 10505 90874 10529 90876
rect 10367 90822 10369 90874
rect 10431 90822 10443 90874
rect 10505 90822 10507 90874
rect 10345 90820 10369 90822
rect 10425 90820 10449 90822
rect 10505 90820 10529 90822
rect 10289 90800 10585 90820
rect 3289 90332 3585 90352
rect 3345 90330 3369 90332
rect 3425 90330 3449 90332
rect 3505 90330 3529 90332
rect 3367 90278 3369 90330
rect 3431 90278 3443 90330
rect 3505 90278 3507 90330
rect 3345 90276 3369 90278
rect 3425 90276 3449 90278
rect 3505 90276 3529 90278
rect 3289 90256 3585 90276
rect 7956 90332 8252 90352
rect 8012 90330 8036 90332
rect 8092 90330 8116 90332
rect 8172 90330 8196 90332
rect 8034 90278 8036 90330
rect 8098 90278 8110 90330
rect 8172 90278 8174 90330
rect 8012 90276 8036 90278
rect 8092 90276 8116 90278
rect 8172 90276 8196 90278
rect 7956 90256 8252 90276
rect 5622 89788 5918 89808
rect 5678 89786 5702 89788
rect 5758 89786 5782 89788
rect 5838 89786 5862 89788
rect 5700 89734 5702 89786
rect 5764 89734 5776 89786
rect 5838 89734 5840 89786
rect 5678 89732 5702 89734
rect 5758 89732 5782 89734
rect 5838 89732 5862 89734
rect 5622 89712 5918 89732
rect 10289 89788 10585 89808
rect 10345 89786 10369 89788
rect 10425 89786 10449 89788
rect 10505 89786 10529 89788
rect 10367 89734 10369 89786
rect 10431 89734 10443 89786
rect 10505 89734 10507 89786
rect 10345 89732 10369 89734
rect 10425 89732 10449 89734
rect 10505 89732 10529 89734
rect 10289 89712 10585 89732
rect 3289 89244 3585 89264
rect 3345 89242 3369 89244
rect 3425 89242 3449 89244
rect 3505 89242 3529 89244
rect 3367 89190 3369 89242
rect 3431 89190 3443 89242
rect 3505 89190 3507 89242
rect 3345 89188 3369 89190
rect 3425 89188 3449 89190
rect 3505 89188 3529 89190
rect 3289 89168 3585 89188
rect 7956 89244 8252 89264
rect 8012 89242 8036 89244
rect 8092 89242 8116 89244
rect 8172 89242 8196 89244
rect 8034 89190 8036 89242
rect 8098 89190 8110 89242
rect 8172 89190 8174 89242
rect 8012 89188 8036 89190
rect 8092 89188 8116 89190
rect 8172 89188 8196 89190
rect 7956 89168 8252 89188
rect 5622 88700 5918 88720
rect 5678 88698 5702 88700
rect 5758 88698 5782 88700
rect 5838 88698 5862 88700
rect 5700 88646 5702 88698
rect 5764 88646 5776 88698
rect 5838 88646 5840 88698
rect 5678 88644 5702 88646
rect 5758 88644 5782 88646
rect 5838 88644 5862 88646
rect 5622 88624 5918 88644
rect 10289 88700 10585 88720
rect 10345 88698 10369 88700
rect 10425 88698 10449 88700
rect 10505 88698 10529 88700
rect 10367 88646 10369 88698
rect 10431 88646 10443 88698
rect 10505 88646 10507 88698
rect 10345 88644 10369 88646
rect 10425 88644 10449 88646
rect 10505 88644 10529 88646
rect 10289 88624 10585 88644
rect 110 88496 166 88505
rect 110 88431 166 88440
rect 124 85241 152 88431
rect 3289 88156 3585 88176
rect 3345 88154 3369 88156
rect 3425 88154 3449 88156
rect 3505 88154 3529 88156
rect 3367 88102 3369 88154
rect 3431 88102 3443 88154
rect 3505 88102 3507 88154
rect 3345 88100 3369 88102
rect 3425 88100 3449 88102
rect 3505 88100 3529 88102
rect 3289 88080 3585 88100
rect 7956 88156 8252 88176
rect 8012 88154 8036 88156
rect 8092 88154 8116 88156
rect 8172 88154 8196 88156
rect 8034 88102 8036 88154
rect 8098 88102 8110 88154
rect 8172 88102 8174 88154
rect 8012 88100 8036 88102
rect 8092 88100 8116 88102
rect 8172 88100 8196 88102
rect 7956 88080 8252 88100
rect 5622 87612 5918 87632
rect 5678 87610 5702 87612
rect 5758 87610 5782 87612
rect 5838 87610 5862 87612
rect 5700 87558 5702 87610
rect 5764 87558 5776 87610
rect 5838 87558 5840 87610
rect 5678 87556 5702 87558
rect 5758 87556 5782 87558
rect 5838 87556 5862 87558
rect 5622 87536 5918 87556
rect 10289 87612 10585 87632
rect 10345 87610 10369 87612
rect 10425 87610 10449 87612
rect 10505 87610 10529 87612
rect 10367 87558 10369 87610
rect 10431 87558 10443 87610
rect 10505 87558 10507 87610
rect 10345 87556 10369 87558
rect 10425 87556 10449 87558
rect 10505 87556 10529 87558
rect 10289 87536 10585 87556
rect 3289 87068 3585 87088
rect 3345 87066 3369 87068
rect 3425 87066 3449 87068
rect 3505 87066 3529 87068
rect 3367 87014 3369 87066
rect 3431 87014 3443 87066
rect 3505 87014 3507 87066
rect 3345 87012 3369 87014
rect 3425 87012 3449 87014
rect 3505 87012 3529 87014
rect 3289 86992 3585 87012
rect 7956 87068 8252 87088
rect 8012 87066 8036 87068
rect 8092 87066 8116 87068
rect 8172 87066 8196 87068
rect 8034 87014 8036 87066
rect 8098 87014 8110 87066
rect 8172 87014 8174 87066
rect 8012 87012 8036 87014
rect 8092 87012 8116 87014
rect 8172 87012 8196 87014
rect 7956 86992 8252 87012
rect 5622 86524 5918 86544
rect 5678 86522 5702 86524
rect 5758 86522 5782 86524
rect 5838 86522 5862 86524
rect 5700 86470 5702 86522
rect 5764 86470 5776 86522
rect 5838 86470 5840 86522
rect 5678 86468 5702 86470
rect 5758 86468 5782 86470
rect 5838 86468 5862 86470
rect 5622 86448 5918 86468
rect 10289 86524 10585 86544
rect 10345 86522 10369 86524
rect 10425 86522 10449 86524
rect 10505 86522 10529 86524
rect 10367 86470 10369 86522
rect 10431 86470 10443 86522
rect 10505 86470 10507 86522
rect 10345 86468 10369 86470
rect 10425 86468 10449 86470
rect 10505 86468 10529 86470
rect 10289 86448 10585 86468
rect 3289 85980 3585 86000
rect 3345 85978 3369 85980
rect 3425 85978 3449 85980
rect 3505 85978 3529 85980
rect 3367 85926 3369 85978
rect 3431 85926 3443 85978
rect 3505 85926 3507 85978
rect 3345 85924 3369 85926
rect 3425 85924 3449 85926
rect 3505 85924 3529 85926
rect 3289 85904 3585 85924
rect 7956 85980 8252 86000
rect 8012 85978 8036 85980
rect 8092 85978 8116 85980
rect 8172 85978 8196 85980
rect 8034 85926 8036 85978
rect 8098 85926 8110 85978
rect 8172 85926 8174 85978
rect 8012 85924 8036 85926
rect 8092 85924 8116 85926
rect 8172 85924 8196 85926
rect 7956 85904 8252 85924
rect 5622 85436 5918 85456
rect 5678 85434 5702 85436
rect 5758 85434 5782 85436
rect 5838 85434 5862 85436
rect 5700 85382 5702 85434
rect 5764 85382 5776 85434
rect 5838 85382 5840 85434
rect 5678 85380 5702 85382
rect 5758 85380 5782 85382
rect 5838 85380 5862 85382
rect 5622 85360 5918 85380
rect 10289 85436 10585 85456
rect 10345 85434 10369 85436
rect 10425 85434 10449 85436
rect 10505 85434 10529 85436
rect 10367 85382 10369 85434
rect 10431 85382 10443 85434
rect 10505 85382 10507 85434
rect 10345 85380 10369 85382
rect 10425 85380 10449 85382
rect 10505 85380 10529 85382
rect 10289 85360 10585 85380
rect 10704 85338 10732 91831
rect 10692 85332 10744 85338
rect 10692 85274 10744 85280
rect 110 85232 166 85241
rect 110 85167 166 85176
rect 3289 84892 3585 84912
rect 3345 84890 3369 84892
rect 3425 84890 3449 84892
rect 3505 84890 3529 84892
rect 3367 84838 3369 84890
rect 3431 84838 3443 84890
rect 3505 84838 3507 84890
rect 3345 84836 3369 84838
rect 3425 84836 3449 84838
rect 3505 84836 3529 84838
rect 3289 84816 3585 84836
rect 7956 84892 8252 84912
rect 8012 84890 8036 84892
rect 8092 84890 8116 84892
rect 8172 84890 8196 84892
rect 8034 84838 8036 84890
rect 8098 84838 8110 84890
rect 8172 84838 8174 84890
rect 8012 84836 8036 84838
rect 8092 84836 8116 84838
rect 8172 84836 8196 84838
rect 7956 84816 8252 84836
rect 5622 84348 5918 84368
rect 5678 84346 5702 84348
rect 5758 84346 5782 84348
rect 5838 84346 5862 84348
rect 5700 84294 5702 84346
rect 5764 84294 5776 84346
rect 5838 84294 5840 84346
rect 5678 84292 5702 84294
rect 5758 84292 5782 84294
rect 5838 84292 5862 84294
rect 5622 84272 5918 84292
rect 10289 84348 10585 84368
rect 10345 84346 10369 84348
rect 10425 84346 10449 84348
rect 10505 84346 10529 84348
rect 10367 84294 10369 84346
rect 10431 84294 10443 84346
rect 10505 84294 10507 84346
rect 10345 84292 10369 84294
rect 10425 84292 10449 84294
rect 10505 84292 10529 84294
rect 10289 84272 10585 84292
rect 3289 83804 3585 83824
rect 3345 83802 3369 83804
rect 3425 83802 3449 83804
rect 3505 83802 3529 83804
rect 3367 83750 3369 83802
rect 3431 83750 3443 83802
rect 3505 83750 3507 83802
rect 3345 83748 3369 83750
rect 3425 83748 3449 83750
rect 3505 83748 3529 83750
rect 3289 83728 3585 83748
rect 7956 83804 8252 83824
rect 8012 83802 8036 83804
rect 8092 83802 8116 83804
rect 8172 83802 8196 83804
rect 8034 83750 8036 83802
rect 8098 83750 8110 83802
rect 8172 83750 8174 83802
rect 8012 83748 8036 83750
rect 8092 83748 8116 83750
rect 8172 83748 8196 83750
rect 7956 83728 8252 83748
rect 5622 83260 5918 83280
rect 5678 83258 5702 83260
rect 5758 83258 5782 83260
rect 5838 83258 5862 83260
rect 5700 83206 5702 83258
rect 5764 83206 5776 83258
rect 5838 83206 5840 83258
rect 5678 83204 5702 83206
rect 5758 83204 5782 83206
rect 5838 83204 5862 83206
rect 5622 83184 5918 83204
rect 10289 83260 10585 83280
rect 10345 83258 10369 83260
rect 10425 83258 10449 83260
rect 10505 83258 10529 83260
rect 10367 83206 10369 83258
rect 10431 83206 10443 83258
rect 10505 83206 10507 83258
rect 10345 83204 10369 83206
rect 10425 83204 10449 83206
rect 10505 83204 10529 83206
rect 10289 83184 10585 83204
rect 3289 82716 3585 82736
rect 3345 82714 3369 82716
rect 3425 82714 3449 82716
rect 3505 82714 3529 82716
rect 3367 82662 3369 82714
rect 3431 82662 3443 82714
rect 3505 82662 3507 82714
rect 3345 82660 3369 82662
rect 3425 82660 3449 82662
rect 3505 82660 3529 82662
rect 3289 82640 3585 82660
rect 7956 82716 8252 82736
rect 8012 82714 8036 82716
rect 8092 82714 8116 82716
rect 8172 82714 8196 82716
rect 8034 82662 8036 82714
rect 8098 82662 8110 82714
rect 8172 82662 8174 82714
rect 8012 82660 8036 82662
rect 8092 82660 8116 82662
rect 8172 82660 8196 82662
rect 7956 82640 8252 82660
rect 5622 82172 5918 82192
rect 5678 82170 5702 82172
rect 5758 82170 5782 82172
rect 5838 82170 5862 82172
rect 5700 82118 5702 82170
rect 5764 82118 5776 82170
rect 5838 82118 5840 82170
rect 5678 82116 5702 82118
rect 5758 82116 5782 82118
rect 5838 82116 5862 82118
rect 5622 82096 5918 82116
rect 10289 82172 10585 82192
rect 10345 82170 10369 82172
rect 10425 82170 10449 82172
rect 10505 82170 10529 82172
rect 10367 82118 10369 82170
rect 10431 82118 10443 82170
rect 10505 82118 10507 82170
rect 10345 82116 10369 82118
rect 10425 82116 10449 82118
rect 10505 82116 10529 82118
rect 10289 82096 10585 82116
rect 3289 81628 3585 81648
rect 3345 81626 3369 81628
rect 3425 81626 3449 81628
rect 3505 81626 3529 81628
rect 3367 81574 3369 81626
rect 3431 81574 3443 81626
rect 3505 81574 3507 81626
rect 3345 81572 3369 81574
rect 3425 81572 3449 81574
rect 3505 81572 3529 81574
rect 3289 81552 3585 81572
rect 7956 81628 8252 81648
rect 8012 81626 8036 81628
rect 8092 81626 8116 81628
rect 8172 81626 8196 81628
rect 8034 81574 8036 81626
rect 8098 81574 8110 81626
rect 8172 81574 8174 81626
rect 8012 81572 8036 81574
rect 8092 81572 8116 81574
rect 8172 81572 8196 81574
rect 7956 81552 8252 81572
rect 5622 81084 5918 81104
rect 5678 81082 5702 81084
rect 5758 81082 5782 81084
rect 5838 81082 5862 81084
rect 5700 81030 5702 81082
rect 5764 81030 5776 81082
rect 5838 81030 5840 81082
rect 5678 81028 5702 81030
rect 5758 81028 5782 81030
rect 5838 81028 5862 81030
rect 5622 81008 5918 81028
rect 10289 81084 10585 81104
rect 10345 81082 10369 81084
rect 10425 81082 10449 81084
rect 10505 81082 10529 81084
rect 10367 81030 10369 81082
rect 10431 81030 10443 81082
rect 10505 81030 10507 81082
rect 10345 81028 10369 81030
rect 10425 81028 10449 81030
rect 10505 81028 10529 81030
rect 10289 81008 10585 81028
rect 3289 80540 3585 80560
rect 3345 80538 3369 80540
rect 3425 80538 3449 80540
rect 3505 80538 3529 80540
rect 3367 80486 3369 80538
rect 3431 80486 3443 80538
rect 3505 80486 3507 80538
rect 3345 80484 3369 80486
rect 3425 80484 3449 80486
rect 3505 80484 3529 80486
rect 3289 80464 3585 80484
rect 7956 80540 8252 80560
rect 8012 80538 8036 80540
rect 8092 80538 8116 80540
rect 8172 80538 8196 80540
rect 8034 80486 8036 80538
rect 8098 80486 8110 80538
rect 8172 80486 8174 80538
rect 8012 80484 8036 80486
rect 8092 80484 8116 80486
rect 8172 80484 8196 80486
rect 7956 80464 8252 80484
rect 5622 79996 5918 80016
rect 5678 79994 5702 79996
rect 5758 79994 5782 79996
rect 5838 79994 5862 79996
rect 5700 79942 5702 79994
rect 5764 79942 5776 79994
rect 5838 79942 5840 79994
rect 5678 79940 5702 79942
rect 5758 79940 5782 79942
rect 5838 79940 5862 79942
rect 5622 79920 5918 79940
rect 10289 79996 10585 80016
rect 10345 79994 10369 79996
rect 10425 79994 10449 79996
rect 10505 79994 10529 79996
rect 10367 79942 10369 79994
rect 10431 79942 10443 79994
rect 10505 79942 10507 79994
rect 10345 79940 10369 79942
rect 10425 79940 10449 79942
rect 10505 79940 10529 79942
rect 10289 79920 10585 79940
rect 3289 79452 3585 79472
rect 3345 79450 3369 79452
rect 3425 79450 3449 79452
rect 3505 79450 3529 79452
rect 3367 79398 3369 79450
rect 3431 79398 3443 79450
rect 3505 79398 3507 79450
rect 3345 79396 3369 79398
rect 3425 79396 3449 79398
rect 3505 79396 3529 79398
rect 3289 79376 3585 79396
rect 7956 79452 8252 79472
rect 8012 79450 8036 79452
rect 8092 79450 8116 79452
rect 8172 79450 8196 79452
rect 8034 79398 8036 79450
rect 8098 79398 8110 79450
rect 8172 79398 8174 79450
rect 8012 79396 8036 79398
rect 8092 79396 8116 79398
rect 8172 79396 8196 79398
rect 7956 79376 8252 79396
rect 5622 78908 5918 78928
rect 5678 78906 5702 78908
rect 5758 78906 5782 78908
rect 5838 78906 5862 78908
rect 5700 78854 5702 78906
rect 5764 78854 5776 78906
rect 5838 78854 5840 78906
rect 5678 78852 5702 78854
rect 5758 78852 5782 78854
rect 5838 78852 5862 78854
rect 5622 78832 5918 78852
rect 10289 78908 10585 78928
rect 10345 78906 10369 78908
rect 10425 78906 10449 78908
rect 10505 78906 10529 78908
rect 10367 78854 10369 78906
rect 10431 78854 10443 78906
rect 10505 78854 10507 78906
rect 10345 78852 10369 78854
rect 10425 78852 10449 78854
rect 10505 78852 10529 78854
rect 10289 78832 10585 78852
rect 3289 78364 3585 78384
rect 3345 78362 3369 78364
rect 3425 78362 3449 78364
rect 3505 78362 3529 78364
rect 3367 78310 3369 78362
rect 3431 78310 3443 78362
rect 3505 78310 3507 78362
rect 3345 78308 3369 78310
rect 3425 78308 3449 78310
rect 3505 78308 3529 78310
rect 3289 78288 3585 78308
rect 7956 78364 8252 78384
rect 8012 78362 8036 78364
rect 8092 78362 8116 78364
rect 8172 78362 8196 78364
rect 8034 78310 8036 78362
rect 8098 78310 8110 78362
rect 8172 78310 8174 78362
rect 8012 78308 8036 78310
rect 8092 78308 8116 78310
rect 8172 78308 8196 78310
rect 7956 78288 8252 78308
rect 10966 78296 11022 78305
rect 10966 78231 11022 78240
rect 5622 77820 5918 77840
rect 5678 77818 5702 77820
rect 5758 77818 5782 77820
rect 5838 77818 5862 77820
rect 5700 77766 5702 77818
rect 5764 77766 5776 77818
rect 5838 77766 5840 77818
rect 5678 77764 5702 77766
rect 5758 77764 5782 77766
rect 5838 77764 5862 77766
rect 5622 77744 5918 77764
rect 10289 77820 10585 77840
rect 10345 77818 10369 77820
rect 10425 77818 10449 77820
rect 10505 77818 10529 77820
rect 10367 77766 10369 77818
rect 10431 77766 10443 77818
rect 10505 77766 10507 77818
rect 10345 77764 10369 77766
rect 10425 77764 10449 77766
rect 10505 77764 10529 77766
rect 10289 77744 10585 77764
rect 3289 77276 3585 77296
rect 3345 77274 3369 77276
rect 3425 77274 3449 77276
rect 3505 77274 3529 77276
rect 3367 77222 3369 77274
rect 3431 77222 3443 77274
rect 3505 77222 3507 77274
rect 3345 77220 3369 77222
rect 3425 77220 3449 77222
rect 3505 77220 3529 77222
rect 3289 77200 3585 77220
rect 7956 77276 8252 77296
rect 8012 77274 8036 77276
rect 8092 77274 8116 77276
rect 8172 77274 8196 77276
rect 8034 77222 8036 77274
rect 8098 77222 8110 77274
rect 8172 77222 8174 77274
rect 8012 77220 8036 77222
rect 8092 77220 8116 77222
rect 8172 77220 8196 77222
rect 7956 77200 8252 77220
rect 5622 76732 5918 76752
rect 5678 76730 5702 76732
rect 5758 76730 5782 76732
rect 5838 76730 5862 76732
rect 5700 76678 5702 76730
rect 5764 76678 5776 76730
rect 5838 76678 5840 76730
rect 5678 76676 5702 76678
rect 5758 76676 5782 76678
rect 5838 76676 5862 76678
rect 5622 76656 5918 76676
rect 10289 76732 10585 76752
rect 10345 76730 10369 76732
rect 10425 76730 10449 76732
rect 10505 76730 10529 76732
rect 10367 76678 10369 76730
rect 10431 76678 10443 76730
rect 10505 76678 10507 76730
rect 10345 76676 10369 76678
rect 10425 76676 10449 76678
rect 10505 76676 10529 76678
rect 10289 76656 10585 76676
rect 3289 76188 3585 76208
rect 3345 76186 3369 76188
rect 3425 76186 3449 76188
rect 3505 76186 3529 76188
rect 3367 76134 3369 76186
rect 3431 76134 3443 76186
rect 3505 76134 3507 76186
rect 3345 76132 3369 76134
rect 3425 76132 3449 76134
rect 3505 76132 3529 76134
rect 3289 76112 3585 76132
rect 7956 76188 8252 76208
rect 8012 76186 8036 76188
rect 8092 76186 8116 76188
rect 8172 76186 8196 76188
rect 8034 76134 8036 76186
rect 8098 76134 8110 76186
rect 8172 76134 8174 76186
rect 8012 76132 8036 76134
rect 8092 76132 8116 76134
rect 8172 76132 8196 76134
rect 7956 76112 8252 76132
rect 5622 75644 5918 75664
rect 5678 75642 5702 75644
rect 5758 75642 5782 75644
rect 5838 75642 5862 75644
rect 5700 75590 5702 75642
rect 5764 75590 5776 75642
rect 5838 75590 5840 75642
rect 5678 75588 5702 75590
rect 5758 75588 5782 75590
rect 5838 75588 5862 75590
rect 5622 75568 5918 75588
rect 10289 75644 10585 75664
rect 10345 75642 10369 75644
rect 10425 75642 10449 75644
rect 10505 75642 10529 75644
rect 10367 75590 10369 75642
rect 10431 75590 10443 75642
rect 10505 75590 10507 75642
rect 10345 75588 10369 75590
rect 10425 75588 10449 75590
rect 10505 75588 10529 75590
rect 10289 75568 10585 75588
rect 3289 75100 3585 75120
rect 3345 75098 3369 75100
rect 3425 75098 3449 75100
rect 3505 75098 3529 75100
rect 3367 75046 3369 75098
rect 3431 75046 3443 75098
rect 3505 75046 3507 75098
rect 3345 75044 3369 75046
rect 3425 75044 3449 75046
rect 3505 75044 3529 75046
rect 3289 75024 3585 75044
rect 7956 75100 8252 75120
rect 8012 75098 8036 75100
rect 8092 75098 8116 75100
rect 8172 75098 8196 75100
rect 8034 75046 8036 75098
rect 8098 75046 8110 75098
rect 8172 75046 8174 75098
rect 8012 75044 8036 75046
rect 8092 75044 8116 75046
rect 8172 75044 8196 75046
rect 7956 75024 8252 75044
rect 110 74896 166 74905
rect 110 74831 166 74840
rect 124 71641 152 74831
rect 5622 74556 5918 74576
rect 5678 74554 5702 74556
rect 5758 74554 5782 74556
rect 5838 74554 5862 74556
rect 5700 74502 5702 74554
rect 5764 74502 5776 74554
rect 5838 74502 5840 74554
rect 5678 74500 5702 74502
rect 5758 74500 5782 74502
rect 5838 74500 5862 74502
rect 5622 74480 5918 74500
rect 10289 74556 10585 74576
rect 10345 74554 10369 74556
rect 10425 74554 10449 74556
rect 10505 74554 10529 74556
rect 10367 74502 10369 74554
rect 10431 74502 10443 74554
rect 10505 74502 10507 74554
rect 10345 74500 10369 74502
rect 10425 74500 10449 74502
rect 10505 74500 10529 74502
rect 10289 74480 10585 74500
rect 3289 74012 3585 74032
rect 3345 74010 3369 74012
rect 3425 74010 3449 74012
rect 3505 74010 3529 74012
rect 3367 73958 3369 74010
rect 3431 73958 3443 74010
rect 3505 73958 3507 74010
rect 3345 73956 3369 73958
rect 3425 73956 3449 73958
rect 3505 73956 3529 73958
rect 3289 73936 3585 73956
rect 7956 74012 8252 74032
rect 8012 74010 8036 74012
rect 8092 74010 8116 74012
rect 8172 74010 8196 74012
rect 8034 73958 8036 74010
rect 8098 73958 8110 74010
rect 8172 73958 8174 74010
rect 8012 73956 8036 73958
rect 8092 73956 8116 73958
rect 8172 73956 8196 73958
rect 7956 73936 8252 73956
rect 5622 73468 5918 73488
rect 5678 73466 5702 73468
rect 5758 73466 5782 73468
rect 5838 73466 5862 73468
rect 5700 73414 5702 73466
rect 5764 73414 5776 73466
rect 5838 73414 5840 73466
rect 5678 73412 5702 73414
rect 5758 73412 5782 73414
rect 5838 73412 5862 73414
rect 5622 73392 5918 73412
rect 10289 73468 10585 73488
rect 10345 73466 10369 73468
rect 10425 73466 10449 73468
rect 10505 73466 10529 73468
rect 10367 73414 10369 73466
rect 10431 73414 10443 73466
rect 10505 73414 10507 73466
rect 10345 73412 10369 73414
rect 10425 73412 10449 73414
rect 10505 73412 10529 73414
rect 10289 73392 10585 73412
rect 3289 72924 3585 72944
rect 3345 72922 3369 72924
rect 3425 72922 3449 72924
rect 3505 72922 3529 72924
rect 3367 72870 3369 72922
rect 3431 72870 3443 72922
rect 3505 72870 3507 72922
rect 3345 72868 3369 72870
rect 3425 72868 3449 72870
rect 3505 72868 3529 72870
rect 3289 72848 3585 72868
rect 7956 72924 8252 72944
rect 8012 72922 8036 72924
rect 8092 72922 8116 72924
rect 8172 72922 8196 72924
rect 8034 72870 8036 72922
rect 8098 72870 8110 72922
rect 8172 72870 8174 72922
rect 8012 72868 8036 72870
rect 8092 72868 8116 72870
rect 8172 72868 8196 72870
rect 7956 72848 8252 72868
rect 5622 72380 5918 72400
rect 5678 72378 5702 72380
rect 5758 72378 5782 72380
rect 5838 72378 5862 72380
rect 5700 72326 5702 72378
rect 5764 72326 5776 72378
rect 5838 72326 5840 72378
rect 5678 72324 5702 72326
rect 5758 72324 5782 72326
rect 5838 72324 5862 72326
rect 5622 72304 5918 72324
rect 10289 72380 10585 72400
rect 10345 72378 10369 72380
rect 10425 72378 10449 72380
rect 10505 72378 10529 72380
rect 10367 72326 10369 72378
rect 10431 72326 10443 72378
rect 10505 72326 10507 72378
rect 10345 72324 10369 72326
rect 10425 72324 10449 72326
rect 10505 72324 10529 72326
rect 10289 72304 10585 72324
rect 3289 71836 3585 71856
rect 3345 71834 3369 71836
rect 3425 71834 3449 71836
rect 3505 71834 3529 71836
rect 3367 71782 3369 71834
rect 3431 71782 3443 71834
rect 3505 71782 3507 71834
rect 3345 71780 3369 71782
rect 3425 71780 3449 71782
rect 3505 71780 3529 71782
rect 3289 71760 3585 71780
rect 7956 71836 8252 71856
rect 8012 71834 8036 71836
rect 8092 71834 8116 71836
rect 8172 71834 8196 71836
rect 8034 71782 8036 71834
rect 8098 71782 8110 71834
rect 8172 71782 8174 71834
rect 8012 71780 8036 71782
rect 8092 71780 8116 71782
rect 8172 71780 8196 71782
rect 7956 71760 8252 71780
rect 10980 71738 11008 78231
rect 10968 71732 11020 71738
rect 10968 71674 11020 71680
rect 110 71632 166 71641
rect 110 71567 166 71576
rect 5622 71292 5918 71312
rect 5678 71290 5702 71292
rect 5758 71290 5782 71292
rect 5838 71290 5862 71292
rect 5700 71238 5702 71290
rect 5764 71238 5776 71290
rect 5838 71238 5840 71290
rect 5678 71236 5702 71238
rect 5758 71236 5782 71238
rect 5838 71236 5862 71238
rect 5622 71216 5918 71236
rect 10289 71292 10585 71312
rect 10345 71290 10369 71292
rect 10425 71290 10449 71292
rect 10505 71290 10529 71292
rect 10367 71238 10369 71290
rect 10431 71238 10443 71290
rect 10505 71238 10507 71290
rect 10345 71236 10369 71238
rect 10425 71236 10449 71238
rect 10505 71236 10529 71238
rect 10289 71216 10585 71236
rect 3289 70748 3585 70768
rect 3345 70746 3369 70748
rect 3425 70746 3449 70748
rect 3505 70746 3529 70748
rect 3367 70694 3369 70746
rect 3431 70694 3443 70746
rect 3505 70694 3507 70746
rect 3345 70692 3369 70694
rect 3425 70692 3449 70694
rect 3505 70692 3529 70694
rect 3289 70672 3585 70692
rect 7956 70748 8252 70768
rect 8012 70746 8036 70748
rect 8092 70746 8116 70748
rect 8172 70746 8196 70748
rect 8034 70694 8036 70746
rect 8098 70694 8110 70746
rect 8172 70694 8174 70746
rect 8012 70692 8036 70694
rect 8092 70692 8116 70694
rect 8172 70692 8196 70694
rect 7956 70672 8252 70692
rect 5622 70204 5918 70224
rect 5678 70202 5702 70204
rect 5758 70202 5782 70204
rect 5838 70202 5862 70204
rect 5700 70150 5702 70202
rect 5764 70150 5776 70202
rect 5838 70150 5840 70202
rect 5678 70148 5702 70150
rect 5758 70148 5782 70150
rect 5838 70148 5862 70150
rect 5622 70128 5918 70148
rect 10289 70204 10585 70224
rect 10345 70202 10369 70204
rect 10425 70202 10449 70204
rect 10505 70202 10529 70204
rect 10367 70150 10369 70202
rect 10431 70150 10443 70202
rect 10505 70150 10507 70202
rect 10345 70148 10369 70150
rect 10425 70148 10449 70150
rect 10505 70148 10529 70150
rect 10289 70128 10585 70148
rect 3289 69660 3585 69680
rect 3345 69658 3369 69660
rect 3425 69658 3449 69660
rect 3505 69658 3529 69660
rect 3367 69606 3369 69658
rect 3431 69606 3443 69658
rect 3505 69606 3507 69658
rect 3345 69604 3369 69606
rect 3425 69604 3449 69606
rect 3505 69604 3529 69606
rect 3289 69584 3585 69604
rect 7956 69660 8252 69680
rect 8012 69658 8036 69660
rect 8092 69658 8116 69660
rect 8172 69658 8196 69660
rect 8034 69606 8036 69658
rect 8098 69606 8110 69658
rect 8172 69606 8174 69658
rect 8012 69604 8036 69606
rect 8092 69604 8116 69606
rect 8172 69604 8196 69606
rect 7956 69584 8252 69604
rect 5622 69116 5918 69136
rect 5678 69114 5702 69116
rect 5758 69114 5782 69116
rect 5838 69114 5862 69116
rect 5700 69062 5702 69114
rect 5764 69062 5776 69114
rect 5838 69062 5840 69114
rect 5678 69060 5702 69062
rect 5758 69060 5782 69062
rect 5838 69060 5862 69062
rect 5622 69040 5918 69060
rect 10289 69116 10585 69136
rect 10345 69114 10369 69116
rect 10425 69114 10449 69116
rect 10505 69114 10529 69116
rect 10367 69062 10369 69114
rect 10431 69062 10443 69114
rect 10505 69062 10507 69114
rect 10345 69060 10369 69062
rect 10425 69060 10449 69062
rect 10505 69060 10529 69062
rect 10289 69040 10585 69060
rect 3289 68572 3585 68592
rect 3345 68570 3369 68572
rect 3425 68570 3449 68572
rect 3505 68570 3529 68572
rect 3367 68518 3369 68570
rect 3431 68518 3443 68570
rect 3505 68518 3507 68570
rect 3345 68516 3369 68518
rect 3425 68516 3449 68518
rect 3505 68516 3529 68518
rect 3289 68496 3585 68516
rect 7956 68572 8252 68592
rect 8012 68570 8036 68572
rect 8092 68570 8116 68572
rect 8172 68570 8196 68572
rect 8034 68518 8036 68570
rect 8098 68518 8110 68570
rect 8172 68518 8174 68570
rect 8012 68516 8036 68518
rect 8092 68516 8116 68518
rect 8172 68516 8196 68518
rect 7956 68496 8252 68516
rect 5622 68028 5918 68048
rect 5678 68026 5702 68028
rect 5758 68026 5782 68028
rect 5838 68026 5862 68028
rect 5700 67974 5702 68026
rect 5764 67974 5776 68026
rect 5838 67974 5840 68026
rect 5678 67972 5702 67974
rect 5758 67972 5782 67974
rect 5838 67972 5862 67974
rect 5622 67952 5918 67972
rect 10289 68028 10585 68048
rect 10345 68026 10369 68028
rect 10425 68026 10449 68028
rect 10505 68026 10529 68028
rect 10367 67974 10369 68026
rect 10431 67974 10443 68026
rect 10505 67974 10507 68026
rect 10345 67972 10369 67974
rect 10425 67972 10449 67974
rect 10505 67972 10529 67974
rect 10289 67952 10585 67972
rect 3289 67484 3585 67504
rect 3345 67482 3369 67484
rect 3425 67482 3449 67484
rect 3505 67482 3529 67484
rect 3367 67430 3369 67482
rect 3431 67430 3443 67482
rect 3505 67430 3507 67482
rect 3345 67428 3369 67430
rect 3425 67428 3449 67430
rect 3505 67428 3529 67430
rect 3289 67408 3585 67428
rect 7956 67484 8252 67504
rect 8012 67482 8036 67484
rect 8092 67482 8116 67484
rect 8172 67482 8196 67484
rect 8034 67430 8036 67482
rect 8098 67430 8110 67482
rect 8172 67430 8174 67482
rect 8012 67428 8036 67430
rect 8092 67428 8116 67430
rect 8172 67428 8196 67430
rect 7956 67408 8252 67428
rect 5622 66940 5918 66960
rect 5678 66938 5702 66940
rect 5758 66938 5782 66940
rect 5838 66938 5862 66940
rect 5700 66886 5702 66938
rect 5764 66886 5776 66938
rect 5838 66886 5840 66938
rect 5678 66884 5702 66886
rect 5758 66884 5782 66886
rect 5838 66884 5862 66886
rect 5622 66864 5918 66884
rect 10289 66940 10585 66960
rect 10345 66938 10369 66940
rect 10425 66938 10449 66940
rect 10505 66938 10529 66940
rect 10367 66886 10369 66938
rect 10431 66886 10443 66938
rect 10505 66886 10507 66938
rect 10345 66884 10369 66886
rect 10425 66884 10449 66886
rect 10505 66884 10529 66886
rect 10289 66864 10585 66884
rect 3289 66396 3585 66416
rect 3345 66394 3369 66396
rect 3425 66394 3449 66396
rect 3505 66394 3529 66396
rect 3367 66342 3369 66394
rect 3431 66342 3443 66394
rect 3505 66342 3507 66394
rect 3345 66340 3369 66342
rect 3425 66340 3449 66342
rect 3505 66340 3529 66342
rect 3289 66320 3585 66340
rect 7956 66396 8252 66416
rect 8012 66394 8036 66396
rect 8092 66394 8116 66396
rect 8172 66394 8196 66396
rect 8034 66342 8036 66394
rect 8098 66342 8110 66394
rect 8172 66342 8174 66394
rect 8012 66340 8036 66342
rect 8092 66340 8116 66342
rect 8172 66340 8196 66342
rect 7956 66320 8252 66340
rect 10140 66020 10192 66026
rect 10140 65962 10192 65968
rect 5622 65852 5918 65872
rect 5678 65850 5702 65852
rect 5758 65850 5782 65852
rect 5838 65850 5862 65852
rect 5700 65798 5702 65850
rect 5764 65798 5776 65850
rect 5838 65798 5840 65850
rect 5678 65796 5702 65798
rect 5758 65796 5782 65798
rect 5838 65796 5862 65798
rect 5622 65776 5918 65796
rect 3289 65308 3585 65328
rect 3345 65306 3369 65308
rect 3425 65306 3449 65308
rect 3505 65306 3529 65308
rect 3367 65254 3369 65306
rect 3431 65254 3443 65306
rect 3505 65254 3507 65306
rect 3345 65252 3369 65254
rect 3425 65252 3449 65254
rect 3505 65252 3529 65254
rect 3289 65232 3585 65252
rect 7956 65308 8252 65328
rect 8012 65306 8036 65308
rect 8092 65306 8116 65308
rect 8172 65306 8196 65308
rect 8034 65254 8036 65306
rect 8098 65254 8110 65306
rect 8172 65254 8174 65306
rect 8012 65252 8036 65254
rect 8092 65252 8116 65254
rect 8172 65252 8196 65254
rect 7956 65232 8252 65252
rect 5622 64764 5918 64784
rect 5678 64762 5702 64764
rect 5758 64762 5782 64764
rect 5838 64762 5862 64764
rect 5700 64710 5702 64762
rect 5764 64710 5776 64762
rect 5838 64710 5840 64762
rect 5678 64708 5702 64710
rect 5758 64708 5782 64710
rect 5838 64708 5862 64710
rect 5622 64688 5918 64708
rect 3289 64220 3585 64240
rect 3345 64218 3369 64220
rect 3425 64218 3449 64220
rect 3505 64218 3529 64220
rect 3367 64166 3369 64218
rect 3431 64166 3443 64218
rect 3505 64166 3507 64218
rect 3345 64164 3369 64166
rect 3425 64164 3449 64166
rect 3505 64164 3529 64166
rect 3289 64144 3585 64164
rect 7956 64220 8252 64240
rect 8012 64218 8036 64220
rect 8092 64218 8116 64220
rect 8172 64218 8196 64220
rect 8034 64166 8036 64218
rect 8098 64166 8110 64218
rect 8172 64166 8174 64218
rect 8012 64164 8036 64166
rect 8092 64164 8116 64166
rect 8172 64164 8196 64166
rect 7956 64144 8252 64164
rect 5622 63676 5918 63696
rect 5678 63674 5702 63676
rect 5758 63674 5782 63676
rect 5838 63674 5862 63676
rect 5700 63622 5702 63674
rect 5764 63622 5776 63674
rect 5838 63622 5840 63674
rect 5678 63620 5702 63622
rect 5758 63620 5782 63622
rect 5838 63620 5862 63622
rect 5622 63600 5918 63620
rect 3289 63132 3585 63152
rect 3345 63130 3369 63132
rect 3425 63130 3449 63132
rect 3505 63130 3529 63132
rect 3367 63078 3369 63130
rect 3431 63078 3443 63130
rect 3505 63078 3507 63130
rect 3345 63076 3369 63078
rect 3425 63076 3449 63078
rect 3505 63076 3529 63078
rect 3289 63056 3585 63076
rect 7956 63132 8252 63152
rect 8012 63130 8036 63132
rect 8092 63130 8116 63132
rect 8172 63130 8196 63132
rect 8034 63078 8036 63130
rect 8098 63078 8110 63130
rect 8172 63078 8174 63130
rect 8012 63076 8036 63078
rect 8092 63076 8116 63078
rect 8172 63076 8196 63078
rect 7956 63056 8252 63076
rect 5622 62588 5918 62608
rect 5678 62586 5702 62588
rect 5758 62586 5782 62588
rect 5838 62586 5862 62588
rect 5700 62534 5702 62586
rect 5764 62534 5776 62586
rect 5838 62534 5840 62586
rect 5678 62532 5702 62534
rect 5758 62532 5782 62534
rect 5838 62532 5862 62534
rect 5622 62512 5918 62532
rect 3289 62044 3585 62064
rect 3345 62042 3369 62044
rect 3425 62042 3449 62044
rect 3505 62042 3529 62044
rect 3367 61990 3369 62042
rect 3431 61990 3443 62042
rect 3505 61990 3507 62042
rect 3345 61988 3369 61990
rect 3425 61988 3449 61990
rect 3505 61988 3529 61990
rect 3289 61968 3585 61988
rect 7956 62044 8252 62064
rect 8012 62042 8036 62044
rect 8092 62042 8116 62044
rect 8172 62042 8196 62044
rect 8034 61990 8036 62042
rect 8098 61990 8110 62042
rect 8172 61990 8174 62042
rect 8012 61988 8036 61990
rect 8092 61988 8116 61990
rect 8172 61988 8196 61990
rect 7956 61968 8252 61988
rect 5622 61500 5918 61520
rect 5678 61498 5702 61500
rect 5758 61498 5782 61500
rect 5838 61498 5862 61500
rect 5700 61446 5702 61498
rect 5764 61446 5776 61498
rect 5838 61446 5840 61498
rect 5678 61444 5702 61446
rect 5758 61444 5782 61446
rect 5838 61444 5862 61446
rect 5622 61424 5918 61444
rect 110 61296 166 61305
rect 110 61231 166 61240
rect 124 58585 152 61231
rect 3289 60956 3585 60976
rect 3345 60954 3369 60956
rect 3425 60954 3449 60956
rect 3505 60954 3529 60956
rect 3367 60902 3369 60954
rect 3431 60902 3443 60954
rect 3505 60902 3507 60954
rect 3345 60900 3369 60902
rect 3425 60900 3449 60902
rect 3505 60900 3529 60902
rect 3289 60880 3585 60900
rect 7956 60956 8252 60976
rect 8012 60954 8036 60956
rect 8092 60954 8116 60956
rect 8172 60954 8196 60956
rect 8034 60902 8036 60954
rect 8098 60902 8110 60954
rect 8172 60902 8174 60954
rect 8012 60900 8036 60902
rect 8092 60900 8116 60902
rect 8172 60900 8196 60902
rect 7956 60880 8252 60900
rect 5622 60412 5918 60432
rect 5678 60410 5702 60412
rect 5758 60410 5782 60412
rect 5838 60410 5862 60412
rect 5700 60358 5702 60410
rect 5764 60358 5776 60410
rect 5838 60358 5840 60410
rect 5678 60356 5702 60358
rect 5758 60356 5782 60358
rect 5838 60356 5862 60358
rect 5622 60336 5918 60356
rect 3289 59868 3585 59888
rect 3345 59866 3369 59868
rect 3425 59866 3449 59868
rect 3505 59866 3529 59868
rect 3367 59814 3369 59866
rect 3431 59814 3443 59866
rect 3505 59814 3507 59866
rect 3345 59812 3369 59814
rect 3425 59812 3449 59814
rect 3505 59812 3529 59814
rect 3289 59792 3585 59812
rect 7956 59868 8252 59888
rect 8012 59866 8036 59868
rect 8092 59866 8116 59868
rect 8172 59866 8196 59868
rect 8034 59814 8036 59866
rect 8098 59814 8110 59866
rect 8172 59814 8174 59866
rect 8012 59812 8036 59814
rect 8092 59812 8116 59814
rect 8172 59812 8196 59814
rect 7956 59792 8252 59812
rect 5622 59324 5918 59344
rect 5678 59322 5702 59324
rect 5758 59322 5782 59324
rect 5838 59322 5862 59324
rect 5700 59270 5702 59322
rect 5764 59270 5776 59322
rect 5838 59270 5840 59322
rect 5678 59268 5702 59270
rect 5758 59268 5782 59270
rect 5838 59268 5862 59270
rect 5622 59248 5918 59268
rect 3289 58780 3585 58800
rect 3345 58778 3369 58780
rect 3425 58778 3449 58780
rect 3505 58778 3529 58780
rect 3367 58726 3369 58778
rect 3431 58726 3443 58778
rect 3505 58726 3507 58778
rect 3345 58724 3369 58726
rect 3425 58724 3449 58726
rect 3505 58724 3529 58726
rect 3289 58704 3585 58724
rect 7956 58780 8252 58800
rect 8012 58778 8036 58780
rect 8092 58778 8116 58780
rect 8172 58778 8196 58780
rect 8034 58726 8036 58778
rect 8098 58726 8110 58778
rect 8172 58726 8174 58778
rect 8012 58724 8036 58726
rect 8092 58724 8116 58726
rect 8172 58724 8196 58726
rect 7956 58704 8252 58724
rect 110 58576 166 58585
rect 110 58511 166 58520
rect 5622 58236 5918 58256
rect 5678 58234 5702 58236
rect 5758 58234 5782 58236
rect 5838 58234 5862 58236
rect 5700 58182 5702 58234
rect 5764 58182 5776 58234
rect 5838 58182 5840 58234
rect 5678 58180 5702 58182
rect 5758 58180 5782 58182
rect 5838 58180 5862 58182
rect 5622 58160 5918 58180
rect 3289 57692 3585 57712
rect 3345 57690 3369 57692
rect 3425 57690 3449 57692
rect 3505 57690 3529 57692
rect 3367 57638 3369 57690
rect 3431 57638 3443 57690
rect 3505 57638 3507 57690
rect 3345 57636 3369 57638
rect 3425 57636 3449 57638
rect 3505 57636 3529 57638
rect 3289 57616 3585 57636
rect 7956 57692 8252 57712
rect 8012 57690 8036 57692
rect 8092 57690 8116 57692
rect 8172 57690 8196 57692
rect 8034 57638 8036 57690
rect 8098 57638 8110 57690
rect 8172 57638 8174 57690
rect 8012 57636 8036 57638
rect 8092 57636 8116 57638
rect 8172 57636 8196 57638
rect 7956 57616 8252 57636
rect 5622 57148 5918 57168
rect 5678 57146 5702 57148
rect 5758 57146 5782 57148
rect 5838 57146 5862 57148
rect 5700 57094 5702 57146
rect 5764 57094 5776 57146
rect 5838 57094 5840 57146
rect 5678 57092 5702 57094
rect 5758 57092 5782 57094
rect 5838 57092 5862 57094
rect 5622 57072 5918 57092
rect 3289 56604 3585 56624
rect 3345 56602 3369 56604
rect 3425 56602 3449 56604
rect 3505 56602 3529 56604
rect 3367 56550 3369 56602
rect 3431 56550 3443 56602
rect 3505 56550 3507 56602
rect 3345 56548 3369 56550
rect 3425 56548 3449 56550
rect 3505 56548 3529 56550
rect 3289 56528 3585 56548
rect 7956 56604 8252 56624
rect 8012 56602 8036 56604
rect 8092 56602 8116 56604
rect 8172 56602 8196 56604
rect 8034 56550 8036 56602
rect 8098 56550 8110 56602
rect 8172 56550 8174 56602
rect 8012 56548 8036 56550
rect 8092 56548 8116 56550
rect 8172 56548 8196 56550
rect 7956 56528 8252 56548
rect 5622 56060 5918 56080
rect 5678 56058 5702 56060
rect 5758 56058 5782 56060
rect 5838 56058 5862 56060
rect 5700 56006 5702 56058
rect 5764 56006 5776 56058
rect 5838 56006 5840 56058
rect 5678 56004 5702 56006
rect 5758 56004 5782 56006
rect 5838 56004 5862 56006
rect 5622 55984 5918 56004
rect 3289 55516 3585 55536
rect 3345 55514 3369 55516
rect 3425 55514 3449 55516
rect 3505 55514 3529 55516
rect 3367 55462 3369 55514
rect 3431 55462 3443 55514
rect 3505 55462 3507 55514
rect 3345 55460 3369 55462
rect 3425 55460 3449 55462
rect 3505 55460 3529 55462
rect 3289 55440 3585 55460
rect 7956 55516 8252 55536
rect 8012 55514 8036 55516
rect 8092 55514 8116 55516
rect 8172 55514 8196 55516
rect 8034 55462 8036 55514
rect 8098 55462 8110 55514
rect 8172 55462 8174 55514
rect 8012 55460 8036 55462
rect 8092 55460 8116 55462
rect 8172 55460 8196 55462
rect 7956 55440 8252 55460
rect 5622 54972 5918 54992
rect 5678 54970 5702 54972
rect 5758 54970 5782 54972
rect 5838 54970 5862 54972
rect 5700 54918 5702 54970
rect 5764 54918 5776 54970
rect 5838 54918 5840 54970
rect 5678 54916 5702 54918
rect 5758 54916 5782 54918
rect 5838 54916 5862 54918
rect 5622 54896 5918 54916
rect 3289 54428 3585 54448
rect 3345 54426 3369 54428
rect 3425 54426 3449 54428
rect 3505 54426 3529 54428
rect 3367 54374 3369 54426
rect 3431 54374 3443 54426
rect 3505 54374 3507 54426
rect 3345 54372 3369 54374
rect 3425 54372 3449 54374
rect 3505 54372 3529 54374
rect 3289 54352 3585 54372
rect 7956 54428 8252 54448
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8034 54374 8036 54426
rect 8098 54374 8110 54426
rect 8172 54374 8174 54426
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 7956 54352 8252 54372
rect 5622 53884 5918 53904
rect 5678 53882 5702 53884
rect 5758 53882 5782 53884
rect 5838 53882 5862 53884
rect 5700 53830 5702 53882
rect 5764 53830 5776 53882
rect 5838 53830 5840 53882
rect 5678 53828 5702 53830
rect 5758 53828 5782 53830
rect 5838 53828 5862 53830
rect 5622 53808 5918 53828
rect 3289 53340 3585 53360
rect 3345 53338 3369 53340
rect 3425 53338 3449 53340
rect 3505 53338 3529 53340
rect 3367 53286 3369 53338
rect 3431 53286 3443 53338
rect 3505 53286 3507 53338
rect 3345 53284 3369 53286
rect 3425 53284 3449 53286
rect 3505 53284 3529 53286
rect 3289 53264 3585 53284
rect 7956 53340 8252 53360
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8034 53286 8036 53338
rect 8098 53286 8110 53338
rect 8172 53286 8174 53338
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 7956 53264 8252 53284
rect 5622 52796 5918 52816
rect 5678 52794 5702 52796
rect 5758 52794 5782 52796
rect 5838 52794 5862 52796
rect 5700 52742 5702 52794
rect 5764 52742 5776 52794
rect 5838 52742 5840 52794
rect 5678 52740 5702 52742
rect 5758 52740 5782 52742
rect 5838 52740 5862 52742
rect 5622 52720 5918 52740
rect 3289 52252 3585 52272
rect 3345 52250 3369 52252
rect 3425 52250 3449 52252
rect 3505 52250 3529 52252
rect 3367 52198 3369 52250
rect 3431 52198 3443 52250
rect 3505 52198 3507 52250
rect 3345 52196 3369 52198
rect 3425 52196 3449 52198
rect 3505 52196 3529 52198
rect 3289 52176 3585 52196
rect 7956 52252 8252 52272
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8034 52198 8036 52250
rect 8098 52198 8110 52250
rect 8172 52198 8174 52250
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 7956 52176 8252 52196
rect 5622 51708 5918 51728
rect 5678 51706 5702 51708
rect 5758 51706 5782 51708
rect 5838 51706 5862 51708
rect 5700 51654 5702 51706
rect 5764 51654 5776 51706
rect 5838 51654 5840 51706
rect 5678 51652 5702 51654
rect 5758 51652 5782 51654
rect 5838 51652 5862 51654
rect 5622 51632 5918 51652
rect 3289 51164 3585 51184
rect 3345 51162 3369 51164
rect 3425 51162 3449 51164
rect 3505 51162 3529 51164
rect 3367 51110 3369 51162
rect 3431 51110 3443 51162
rect 3505 51110 3507 51162
rect 3345 51108 3369 51110
rect 3425 51108 3449 51110
rect 3505 51108 3529 51110
rect 3289 51088 3585 51108
rect 7956 51164 8252 51184
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8034 51110 8036 51162
rect 8098 51110 8110 51162
rect 8172 51110 8174 51162
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 7956 51088 8252 51108
rect 5622 50620 5918 50640
rect 5678 50618 5702 50620
rect 5758 50618 5782 50620
rect 5838 50618 5862 50620
rect 5700 50566 5702 50618
rect 5764 50566 5776 50618
rect 5838 50566 5840 50618
rect 5678 50564 5702 50566
rect 5758 50564 5782 50566
rect 5838 50564 5862 50566
rect 5622 50544 5918 50564
rect 3289 50076 3585 50096
rect 3345 50074 3369 50076
rect 3425 50074 3449 50076
rect 3505 50074 3529 50076
rect 3367 50022 3369 50074
rect 3431 50022 3443 50074
rect 3505 50022 3507 50074
rect 3345 50020 3369 50022
rect 3425 50020 3449 50022
rect 3505 50020 3529 50022
rect 3289 50000 3585 50020
rect 7956 50076 8252 50096
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8034 50022 8036 50074
rect 8098 50022 8110 50074
rect 8172 50022 8174 50074
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 7956 50000 8252 50020
rect 5622 49532 5918 49552
rect 5678 49530 5702 49532
rect 5758 49530 5782 49532
rect 5838 49530 5862 49532
rect 5700 49478 5702 49530
rect 5764 49478 5776 49530
rect 5838 49478 5840 49530
rect 5678 49476 5702 49478
rect 5758 49476 5782 49478
rect 5838 49476 5862 49478
rect 5622 49456 5918 49476
rect 3289 48988 3585 49008
rect 3345 48986 3369 48988
rect 3425 48986 3449 48988
rect 3505 48986 3529 48988
rect 3367 48934 3369 48986
rect 3431 48934 3443 48986
rect 3505 48934 3507 48986
rect 3345 48932 3369 48934
rect 3425 48932 3449 48934
rect 3505 48932 3529 48934
rect 3289 48912 3585 48932
rect 7956 48988 8252 49008
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8034 48934 8036 48986
rect 8098 48934 8110 48986
rect 8172 48934 8174 48986
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 7956 48912 8252 48932
rect 5622 48444 5918 48464
rect 5678 48442 5702 48444
rect 5758 48442 5782 48444
rect 5838 48442 5862 48444
rect 5700 48390 5702 48442
rect 5764 48390 5776 48442
rect 5838 48390 5840 48442
rect 5678 48388 5702 48390
rect 5758 48388 5782 48390
rect 5838 48388 5862 48390
rect 5622 48368 5918 48388
rect 3289 47900 3585 47920
rect 3345 47898 3369 47900
rect 3425 47898 3449 47900
rect 3505 47898 3529 47900
rect 3367 47846 3369 47898
rect 3431 47846 3443 47898
rect 3505 47846 3507 47898
rect 3345 47844 3369 47846
rect 3425 47844 3449 47846
rect 3505 47844 3529 47846
rect 3289 47824 3585 47844
rect 7956 47900 8252 47920
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8034 47846 8036 47898
rect 8098 47846 8110 47898
rect 8172 47846 8174 47898
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 7956 47824 8252 47844
rect 110 47696 166 47705
rect 110 47631 166 47640
rect 124 44849 152 47631
rect 5622 47356 5918 47376
rect 5678 47354 5702 47356
rect 5758 47354 5782 47356
rect 5838 47354 5862 47356
rect 5700 47302 5702 47354
rect 5764 47302 5776 47354
rect 5838 47302 5840 47354
rect 5678 47300 5702 47302
rect 5758 47300 5782 47302
rect 5838 47300 5862 47302
rect 5622 47280 5918 47300
rect 3289 46812 3585 46832
rect 3345 46810 3369 46812
rect 3425 46810 3449 46812
rect 3505 46810 3529 46812
rect 3367 46758 3369 46810
rect 3431 46758 3443 46810
rect 3505 46758 3507 46810
rect 3345 46756 3369 46758
rect 3425 46756 3449 46758
rect 3505 46756 3529 46758
rect 3289 46736 3585 46756
rect 7956 46812 8252 46832
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8034 46758 8036 46810
rect 8098 46758 8110 46810
rect 8172 46758 8174 46810
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 7956 46736 8252 46756
rect 5622 46268 5918 46288
rect 5678 46266 5702 46268
rect 5758 46266 5782 46268
rect 5838 46266 5862 46268
rect 5700 46214 5702 46266
rect 5764 46214 5776 46266
rect 5838 46214 5840 46266
rect 5678 46212 5702 46214
rect 5758 46212 5782 46214
rect 5838 46212 5862 46214
rect 5622 46192 5918 46212
rect 3289 45724 3585 45744
rect 3345 45722 3369 45724
rect 3425 45722 3449 45724
rect 3505 45722 3529 45724
rect 3367 45670 3369 45722
rect 3431 45670 3443 45722
rect 3505 45670 3507 45722
rect 3345 45668 3369 45670
rect 3425 45668 3449 45670
rect 3505 45668 3529 45670
rect 3289 45648 3585 45668
rect 7956 45724 8252 45744
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8034 45670 8036 45722
rect 8098 45670 8110 45722
rect 8172 45670 8174 45722
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 7956 45648 8252 45668
rect 5622 45180 5918 45200
rect 5678 45178 5702 45180
rect 5758 45178 5782 45180
rect 5838 45178 5862 45180
rect 5700 45126 5702 45178
rect 5764 45126 5776 45178
rect 5838 45126 5840 45178
rect 5678 45124 5702 45126
rect 5758 45124 5782 45126
rect 5838 45124 5862 45126
rect 5622 45104 5918 45124
rect 110 44840 166 44849
rect 110 44775 166 44784
rect 3289 44636 3585 44656
rect 3345 44634 3369 44636
rect 3425 44634 3449 44636
rect 3505 44634 3529 44636
rect 3367 44582 3369 44634
rect 3431 44582 3443 44634
rect 3505 44582 3507 44634
rect 3345 44580 3369 44582
rect 3425 44580 3449 44582
rect 3505 44580 3529 44582
rect 3289 44560 3585 44580
rect 7956 44636 8252 44656
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8034 44582 8036 44634
rect 8098 44582 8110 44634
rect 8172 44582 8174 44634
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 7956 44560 8252 44580
rect 5622 44092 5918 44112
rect 5678 44090 5702 44092
rect 5758 44090 5782 44092
rect 5838 44090 5862 44092
rect 5700 44038 5702 44090
rect 5764 44038 5776 44090
rect 5838 44038 5840 44090
rect 5678 44036 5702 44038
rect 5758 44036 5782 44038
rect 5838 44036 5862 44038
rect 5622 44016 5918 44036
rect 3289 43548 3585 43568
rect 3345 43546 3369 43548
rect 3425 43546 3449 43548
rect 3505 43546 3529 43548
rect 3367 43494 3369 43546
rect 3431 43494 3443 43546
rect 3505 43494 3507 43546
rect 3345 43492 3369 43494
rect 3425 43492 3449 43494
rect 3505 43492 3529 43494
rect 3289 43472 3585 43492
rect 7956 43548 8252 43568
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8034 43494 8036 43546
rect 8098 43494 8110 43546
rect 8172 43494 8174 43546
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 7956 43472 8252 43492
rect 5622 43004 5918 43024
rect 5678 43002 5702 43004
rect 5758 43002 5782 43004
rect 5838 43002 5862 43004
rect 5700 42950 5702 43002
rect 5764 42950 5776 43002
rect 5838 42950 5840 43002
rect 5678 42948 5702 42950
rect 5758 42948 5782 42950
rect 5838 42948 5862 42950
rect 5622 42928 5918 42948
rect 3289 42460 3585 42480
rect 3345 42458 3369 42460
rect 3425 42458 3449 42460
rect 3505 42458 3529 42460
rect 3367 42406 3369 42458
rect 3431 42406 3443 42458
rect 3505 42406 3507 42458
rect 3345 42404 3369 42406
rect 3425 42404 3449 42406
rect 3505 42404 3529 42406
rect 3289 42384 3585 42404
rect 7956 42460 8252 42480
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8034 42406 8036 42458
rect 8098 42406 8110 42458
rect 8172 42406 8174 42458
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 7956 42384 8252 42404
rect 5622 41916 5918 41936
rect 5678 41914 5702 41916
rect 5758 41914 5782 41916
rect 5838 41914 5862 41916
rect 5700 41862 5702 41914
rect 5764 41862 5776 41914
rect 5838 41862 5840 41914
rect 5678 41860 5702 41862
rect 5758 41860 5782 41862
rect 5838 41860 5862 41862
rect 5622 41840 5918 41860
rect 3289 41372 3585 41392
rect 3345 41370 3369 41372
rect 3425 41370 3449 41372
rect 3505 41370 3529 41372
rect 3367 41318 3369 41370
rect 3431 41318 3443 41370
rect 3505 41318 3507 41370
rect 3345 41316 3369 41318
rect 3425 41316 3449 41318
rect 3505 41316 3529 41318
rect 3289 41296 3585 41316
rect 7956 41372 8252 41392
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8034 41318 8036 41370
rect 8098 41318 8110 41370
rect 8172 41318 8174 41370
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 7956 41296 8252 41316
rect 5622 40828 5918 40848
rect 5678 40826 5702 40828
rect 5758 40826 5782 40828
rect 5838 40826 5862 40828
rect 5700 40774 5702 40826
rect 5764 40774 5776 40826
rect 5838 40774 5840 40826
rect 5678 40772 5702 40774
rect 5758 40772 5782 40774
rect 5838 40772 5862 40774
rect 5622 40752 5918 40772
rect 3289 40284 3585 40304
rect 3345 40282 3369 40284
rect 3425 40282 3449 40284
rect 3505 40282 3529 40284
rect 3367 40230 3369 40282
rect 3431 40230 3443 40282
rect 3505 40230 3507 40282
rect 3345 40228 3369 40230
rect 3425 40228 3449 40230
rect 3505 40228 3529 40230
rect 3289 40208 3585 40228
rect 7956 40284 8252 40304
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8034 40230 8036 40282
rect 8098 40230 8110 40282
rect 8172 40230 8174 40282
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 7956 40208 8252 40228
rect 5622 39740 5918 39760
rect 5678 39738 5702 39740
rect 5758 39738 5782 39740
rect 5838 39738 5862 39740
rect 5700 39686 5702 39738
rect 5764 39686 5776 39738
rect 5838 39686 5840 39738
rect 5678 39684 5702 39686
rect 5758 39684 5782 39686
rect 5838 39684 5862 39686
rect 5622 39664 5918 39684
rect 3289 39196 3585 39216
rect 3345 39194 3369 39196
rect 3425 39194 3449 39196
rect 3505 39194 3529 39196
rect 3367 39142 3369 39194
rect 3431 39142 3443 39194
rect 3505 39142 3507 39194
rect 3345 39140 3369 39142
rect 3425 39140 3449 39142
rect 3505 39140 3529 39142
rect 3289 39120 3585 39140
rect 7956 39196 8252 39216
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8034 39142 8036 39194
rect 8098 39142 8110 39194
rect 8172 39142 8174 39194
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 7956 39120 8252 39140
rect 5622 38652 5918 38672
rect 5678 38650 5702 38652
rect 5758 38650 5782 38652
rect 5838 38650 5862 38652
rect 5700 38598 5702 38650
rect 5764 38598 5776 38650
rect 5838 38598 5840 38650
rect 5678 38596 5702 38598
rect 5758 38596 5782 38598
rect 5838 38596 5862 38598
rect 5622 38576 5918 38596
rect 3289 38108 3585 38128
rect 3345 38106 3369 38108
rect 3425 38106 3449 38108
rect 3505 38106 3529 38108
rect 3367 38054 3369 38106
rect 3431 38054 3443 38106
rect 3505 38054 3507 38106
rect 3345 38052 3369 38054
rect 3425 38052 3449 38054
rect 3505 38052 3529 38054
rect 3289 38032 3585 38052
rect 7956 38108 8252 38128
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8034 38054 8036 38106
rect 8098 38054 8110 38106
rect 8172 38054 8174 38106
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 7956 38032 8252 38052
rect 5622 37564 5918 37584
rect 5678 37562 5702 37564
rect 5758 37562 5782 37564
rect 5838 37562 5862 37564
rect 5700 37510 5702 37562
rect 5764 37510 5776 37562
rect 5838 37510 5840 37562
rect 5678 37508 5702 37510
rect 5758 37508 5782 37510
rect 5838 37508 5862 37510
rect 5622 37488 5918 37508
rect 3289 37020 3585 37040
rect 3345 37018 3369 37020
rect 3425 37018 3449 37020
rect 3505 37018 3529 37020
rect 3367 36966 3369 37018
rect 3431 36966 3443 37018
rect 3505 36966 3507 37018
rect 3345 36964 3369 36966
rect 3425 36964 3449 36966
rect 3505 36964 3529 36966
rect 3289 36944 3585 36964
rect 7956 37020 8252 37040
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8034 36966 8036 37018
rect 8098 36966 8110 37018
rect 8172 36966 8174 37018
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 7956 36944 8252 36964
rect 5622 36476 5918 36496
rect 5678 36474 5702 36476
rect 5758 36474 5782 36476
rect 5838 36474 5862 36476
rect 5700 36422 5702 36474
rect 5764 36422 5776 36474
rect 5838 36422 5840 36474
rect 5678 36420 5702 36422
rect 5758 36420 5782 36422
rect 5838 36420 5862 36422
rect 5622 36400 5918 36420
rect 3289 35932 3585 35952
rect 3345 35930 3369 35932
rect 3425 35930 3449 35932
rect 3505 35930 3529 35932
rect 3367 35878 3369 35930
rect 3431 35878 3443 35930
rect 3505 35878 3507 35930
rect 3345 35876 3369 35878
rect 3425 35876 3449 35878
rect 3505 35876 3529 35878
rect 3289 35856 3585 35876
rect 7956 35932 8252 35952
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8034 35878 8036 35930
rect 8098 35878 8110 35930
rect 8172 35878 8174 35930
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 7956 35856 8252 35876
rect 5622 35388 5918 35408
rect 5678 35386 5702 35388
rect 5758 35386 5782 35388
rect 5838 35386 5862 35388
rect 5700 35334 5702 35386
rect 5764 35334 5776 35386
rect 5838 35334 5840 35386
rect 5678 35332 5702 35334
rect 5758 35332 5782 35334
rect 5838 35332 5862 35334
rect 5622 35312 5918 35332
rect 3289 34844 3585 34864
rect 3345 34842 3369 34844
rect 3425 34842 3449 34844
rect 3505 34842 3529 34844
rect 3367 34790 3369 34842
rect 3431 34790 3443 34842
rect 3505 34790 3507 34842
rect 3345 34788 3369 34790
rect 3425 34788 3449 34790
rect 3505 34788 3529 34790
rect 3289 34768 3585 34788
rect 7956 34844 8252 34864
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8034 34790 8036 34842
rect 8098 34790 8110 34842
rect 8172 34790 8174 34842
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 7956 34768 8252 34788
rect 5622 34300 5918 34320
rect 5678 34298 5702 34300
rect 5758 34298 5782 34300
rect 5838 34298 5862 34300
rect 5700 34246 5702 34298
rect 5764 34246 5776 34298
rect 5838 34246 5840 34298
rect 5678 34244 5702 34246
rect 5758 34244 5782 34246
rect 5838 34244 5862 34246
rect 5622 34224 5918 34244
rect 110 34096 166 34105
rect 110 34031 166 34040
rect 124 31249 152 34031
rect 3289 33756 3585 33776
rect 3345 33754 3369 33756
rect 3425 33754 3449 33756
rect 3505 33754 3529 33756
rect 3367 33702 3369 33754
rect 3431 33702 3443 33754
rect 3505 33702 3507 33754
rect 3345 33700 3369 33702
rect 3425 33700 3449 33702
rect 3505 33700 3529 33702
rect 3289 33680 3585 33700
rect 7956 33756 8252 33776
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8034 33702 8036 33754
rect 8098 33702 8110 33754
rect 8172 33702 8174 33754
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 7956 33680 8252 33700
rect 5622 33212 5918 33232
rect 5678 33210 5702 33212
rect 5758 33210 5782 33212
rect 5838 33210 5862 33212
rect 5700 33158 5702 33210
rect 5764 33158 5776 33210
rect 5838 33158 5840 33210
rect 5678 33156 5702 33158
rect 5758 33156 5782 33158
rect 5838 33156 5862 33158
rect 5622 33136 5918 33156
rect 3289 32668 3585 32688
rect 3345 32666 3369 32668
rect 3425 32666 3449 32668
rect 3505 32666 3529 32668
rect 3367 32614 3369 32666
rect 3431 32614 3443 32666
rect 3505 32614 3507 32666
rect 3345 32612 3369 32614
rect 3425 32612 3449 32614
rect 3505 32612 3529 32614
rect 3289 32592 3585 32612
rect 7956 32668 8252 32688
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8034 32614 8036 32666
rect 8098 32614 8110 32666
rect 8172 32614 8174 32666
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 7956 32592 8252 32612
rect 5622 32124 5918 32144
rect 5678 32122 5702 32124
rect 5758 32122 5782 32124
rect 5838 32122 5862 32124
rect 5700 32070 5702 32122
rect 5764 32070 5776 32122
rect 5838 32070 5840 32122
rect 5678 32068 5702 32070
rect 5758 32068 5782 32070
rect 5838 32068 5862 32070
rect 5622 32048 5918 32068
rect 3289 31580 3585 31600
rect 3345 31578 3369 31580
rect 3425 31578 3449 31580
rect 3505 31578 3529 31580
rect 3367 31526 3369 31578
rect 3431 31526 3443 31578
rect 3505 31526 3507 31578
rect 3345 31524 3369 31526
rect 3425 31524 3449 31526
rect 3505 31524 3529 31526
rect 3289 31504 3585 31524
rect 7956 31580 8252 31600
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8034 31526 8036 31578
rect 8098 31526 8110 31578
rect 8172 31526 8174 31578
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 7956 31504 8252 31524
rect 110 31240 166 31249
rect 110 31175 166 31184
rect 5622 31036 5918 31056
rect 5678 31034 5702 31036
rect 5758 31034 5782 31036
rect 5838 31034 5862 31036
rect 5700 30982 5702 31034
rect 5764 30982 5776 31034
rect 5838 30982 5840 31034
rect 5678 30980 5702 30982
rect 5758 30980 5782 30982
rect 5838 30980 5862 30982
rect 5622 30960 5918 30980
rect 3289 30492 3585 30512
rect 3345 30490 3369 30492
rect 3425 30490 3449 30492
rect 3505 30490 3529 30492
rect 3367 30438 3369 30490
rect 3431 30438 3443 30490
rect 3505 30438 3507 30490
rect 3345 30436 3369 30438
rect 3425 30436 3449 30438
rect 3505 30436 3529 30438
rect 3289 30416 3585 30436
rect 7956 30492 8252 30512
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8034 30438 8036 30490
rect 8098 30438 8110 30490
rect 8172 30438 8174 30490
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 7956 30416 8252 30436
rect 5622 29948 5918 29968
rect 5678 29946 5702 29948
rect 5758 29946 5782 29948
rect 5838 29946 5862 29948
rect 5700 29894 5702 29946
rect 5764 29894 5776 29946
rect 5838 29894 5840 29946
rect 5678 29892 5702 29894
rect 5758 29892 5782 29894
rect 5838 29892 5862 29894
rect 5622 29872 5918 29892
rect 3289 29404 3585 29424
rect 3345 29402 3369 29404
rect 3425 29402 3449 29404
rect 3505 29402 3529 29404
rect 3367 29350 3369 29402
rect 3431 29350 3443 29402
rect 3505 29350 3507 29402
rect 3345 29348 3369 29350
rect 3425 29348 3449 29350
rect 3505 29348 3529 29350
rect 3289 29328 3585 29348
rect 7956 29404 8252 29424
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8034 29350 8036 29402
rect 8098 29350 8110 29402
rect 8172 29350 8174 29402
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 7956 29328 8252 29348
rect 5622 28860 5918 28880
rect 5678 28858 5702 28860
rect 5758 28858 5782 28860
rect 5838 28858 5862 28860
rect 5700 28806 5702 28858
rect 5764 28806 5776 28858
rect 5838 28806 5840 28858
rect 5678 28804 5702 28806
rect 5758 28804 5782 28806
rect 5838 28804 5862 28806
rect 5622 28784 5918 28804
rect 3289 28316 3585 28336
rect 3345 28314 3369 28316
rect 3425 28314 3449 28316
rect 3505 28314 3529 28316
rect 3367 28262 3369 28314
rect 3431 28262 3443 28314
rect 3505 28262 3507 28314
rect 3345 28260 3369 28262
rect 3425 28260 3449 28262
rect 3505 28260 3529 28262
rect 3289 28240 3585 28260
rect 7956 28316 8252 28336
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8034 28262 8036 28314
rect 8098 28262 8110 28314
rect 8172 28262 8174 28314
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 7956 28240 8252 28260
rect 5622 27772 5918 27792
rect 5678 27770 5702 27772
rect 5758 27770 5782 27772
rect 5838 27770 5862 27772
rect 5700 27718 5702 27770
rect 5764 27718 5776 27770
rect 5838 27718 5840 27770
rect 5678 27716 5702 27718
rect 5758 27716 5782 27718
rect 5838 27716 5862 27718
rect 5622 27696 5918 27716
rect 3289 27228 3585 27248
rect 3345 27226 3369 27228
rect 3425 27226 3449 27228
rect 3505 27226 3529 27228
rect 3367 27174 3369 27226
rect 3431 27174 3443 27226
rect 3505 27174 3507 27226
rect 3345 27172 3369 27174
rect 3425 27172 3449 27174
rect 3505 27172 3529 27174
rect 3289 27152 3585 27172
rect 7956 27228 8252 27248
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8034 27174 8036 27226
rect 8098 27174 8110 27226
rect 8172 27174 8174 27226
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 7956 27152 8252 27172
rect 5622 26684 5918 26704
rect 5678 26682 5702 26684
rect 5758 26682 5782 26684
rect 5838 26682 5862 26684
rect 5700 26630 5702 26682
rect 5764 26630 5776 26682
rect 5838 26630 5840 26682
rect 5678 26628 5702 26630
rect 5758 26628 5782 26630
rect 5838 26628 5862 26630
rect 5622 26608 5918 26628
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 3289 26140 3585 26160
rect 3345 26138 3369 26140
rect 3425 26138 3449 26140
rect 3505 26138 3529 26140
rect 3367 26086 3369 26138
rect 3431 26086 3443 26138
rect 3505 26086 3507 26138
rect 3345 26084 3369 26086
rect 3425 26084 3449 26086
rect 3505 26084 3529 26086
rect 3289 26064 3585 26084
rect 7956 26140 8252 26160
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8034 26086 8036 26138
rect 8098 26086 8110 26138
rect 8172 26086 8174 26138
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 7956 26064 8252 26084
rect 5622 25596 5918 25616
rect 5678 25594 5702 25596
rect 5758 25594 5782 25596
rect 5838 25594 5862 25596
rect 5700 25542 5702 25594
rect 5764 25542 5776 25594
rect 5838 25542 5840 25594
rect 5678 25540 5702 25542
rect 5758 25540 5782 25542
rect 5838 25540 5862 25542
rect 5622 25520 5918 25540
rect 3289 25052 3585 25072
rect 3345 25050 3369 25052
rect 3425 25050 3449 25052
rect 3505 25050 3529 25052
rect 3367 24998 3369 25050
rect 3431 24998 3443 25050
rect 3505 24998 3507 25050
rect 3345 24996 3369 24998
rect 3425 24996 3449 24998
rect 3505 24996 3529 24998
rect 3289 24976 3585 24996
rect 7956 25052 8252 25072
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8034 24998 8036 25050
rect 8098 24998 8110 25050
rect 8172 24998 8174 25050
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 7956 24976 8252 24996
rect 5622 24508 5918 24528
rect 5678 24506 5702 24508
rect 5758 24506 5782 24508
rect 5838 24506 5862 24508
rect 5700 24454 5702 24506
rect 5764 24454 5776 24506
rect 5838 24454 5840 24506
rect 5678 24452 5702 24454
rect 5758 24452 5782 24454
rect 5838 24452 5862 24454
rect 5622 24432 5918 24452
rect 3289 23964 3585 23984
rect 3345 23962 3369 23964
rect 3425 23962 3449 23964
rect 3505 23962 3529 23964
rect 3367 23910 3369 23962
rect 3431 23910 3443 23962
rect 3505 23910 3507 23962
rect 3345 23908 3369 23910
rect 3425 23908 3449 23910
rect 3505 23908 3529 23910
rect 3289 23888 3585 23908
rect 7956 23964 8252 23984
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8034 23910 8036 23962
rect 8098 23910 8110 23962
rect 8172 23910 8174 23962
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 7956 23888 8252 23908
rect 5622 23420 5918 23440
rect 5678 23418 5702 23420
rect 5758 23418 5782 23420
rect 5838 23418 5862 23420
rect 5700 23366 5702 23418
rect 5764 23366 5776 23418
rect 5838 23366 5840 23418
rect 5678 23364 5702 23366
rect 5758 23364 5782 23366
rect 5838 23364 5862 23366
rect 5622 23344 5918 23364
rect 3289 22876 3585 22896
rect 3345 22874 3369 22876
rect 3425 22874 3449 22876
rect 3505 22874 3529 22876
rect 3367 22822 3369 22874
rect 3431 22822 3443 22874
rect 3505 22822 3507 22874
rect 3345 22820 3369 22822
rect 3425 22820 3449 22822
rect 3505 22820 3529 22822
rect 3289 22800 3585 22820
rect 7956 22876 8252 22896
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8034 22822 8036 22874
rect 8098 22822 8110 22874
rect 8172 22822 8174 22874
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 7956 22800 8252 22820
rect 5622 22332 5918 22352
rect 5678 22330 5702 22332
rect 5758 22330 5782 22332
rect 5838 22330 5862 22332
rect 5700 22278 5702 22330
rect 5764 22278 5776 22330
rect 5838 22278 5840 22330
rect 5678 22276 5702 22278
rect 5758 22276 5782 22278
rect 5838 22276 5862 22278
rect 5622 22256 5918 22276
rect 3289 21788 3585 21808
rect 3345 21786 3369 21788
rect 3425 21786 3449 21788
rect 3505 21786 3529 21788
rect 3367 21734 3369 21786
rect 3431 21734 3443 21786
rect 3505 21734 3507 21786
rect 3345 21732 3369 21734
rect 3425 21732 3449 21734
rect 3505 21732 3529 21734
rect 3289 21712 3585 21732
rect 7956 21788 8252 21808
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8034 21734 8036 21786
rect 8098 21734 8110 21786
rect 8172 21734 8174 21786
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 7956 21712 8252 21732
rect 5622 21244 5918 21264
rect 5678 21242 5702 21244
rect 5758 21242 5782 21244
rect 5838 21242 5862 21244
rect 5700 21190 5702 21242
rect 5764 21190 5776 21242
rect 5838 21190 5840 21242
rect 5678 21188 5702 21190
rect 5758 21188 5782 21190
rect 5838 21188 5862 21190
rect 5622 21168 5918 21188
rect 3289 20700 3585 20720
rect 3345 20698 3369 20700
rect 3425 20698 3449 20700
rect 3505 20698 3529 20700
rect 3367 20646 3369 20698
rect 3431 20646 3443 20698
rect 3505 20646 3507 20698
rect 3345 20644 3369 20646
rect 3425 20644 3449 20646
rect 3505 20644 3529 20646
rect 3289 20624 3585 20644
rect 7956 20700 8252 20720
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8034 20646 8036 20698
rect 8098 20646 8110 20698
rect 8172 20646 8174 20698
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 7956 20624 8252 20644
rect 110 20496 166 20505
rect 110 20431 166 20440
rect 124 17241 152 20431
rect 5622 20156 5918 20176
rect 5678 20154 5702 20156
rect 5758 20154 5782 20156
rect 5838 20154 5862 20156
rect 5700 20102 5702 20154
rect 5764 20102 5776 20154
rect 5838 20102 5840 20154
rect 5678 20100 5702 20102
rect 5758 20100 5782 20102
rect 5838 20100 5862 20102
rect 5622 20080 5918 20100
rect 3289 19612 3585 19632
rect 3345 19610 3369 19612
rect 3425 19610 3449 19612
rect 3505 19610 3529 19612
rect 3367 19558 3369 19610
rect 3431 19558 3443 19610
rect 3505 19558 3507 19610
rect 3345 19556 3369 19558
rect 3425 19556 3449 19558
rect 3505 19556 3529 19558
rect 3289 19536 3585 19556
rect 7956 19612 8252 19632
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8034 19558 8036 19610
rect 8098 19558 8110 19610
rect 8172 19558 8174 19610
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 7956 19536 8252 19556
rect 5622 19068 5918 19088
rect 5678 19066 5702 19068
rect 5758 19066 5782 19068
rect 5838 19066 5862 19068
rect 5700 19014 5702 19066
rect 5764 19014 5776 19066
rect 5838 19014 5840 19066
rect 5678 19012 5702 19014
rect 5758 19012 5782 19014
rect 5838 19012 5862 19014
rect 5622 18992 5918 19012
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 3289 18524 3585 18544
rect 3345 18522 3369 18524
rect 3425 18522 3449 18524
rect 3505 18522 3529 18524
rect 3367 18470 3369 18522
rect 3431 18470 3443 18522
rect 3505 18470 3507 18522
rect 3345 18468 3369 18470
rect 3425 18468 3449 18470
rect 3505 18468 3529 18470
rect 3289 18448 3585 18468
rect 7956 18524 8252 18544
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8034 18470 8036 18522
rect 8098 18470 8110 18522
rect 8172 18470 8174 18522
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 7956 18448 8252 18468
rect 8588 18222 8616 18566
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 5622 17980 5918 18000
rect 5678 17978 5702 17980
rect 5758 17978 5782 17980
rect 5838 17978 5862 17980
rect 5700 17926 5702 17978
rect 5764 17926 5776 17978
rect 5838 17926 5840 17978
rect 5678 17924 5702 17926
rect 5758 17924 5782 17926
rect 5838 17924 5862 17926
rect 5622 17904 5918 17924
rect 3289 17436 3585 17456
rect 3345 17434 3369 17436
rect 3425 17434 3449 17436
rect 3505 17434 3529 17436
rect 3367 17382 3369 17434
rect 3431 17382 3443 17434
rect 3505 17382 3507 17434
rect 3345 17380 3369 17382
rect 3425 17380 3449 17382
rect 3505 17380 3529 17382
rect 3289 17360 3585 17380
rect 7956 17436 8252 17456
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8034 17382 8036 17434
rect 8098 17382 8110 17434
rect 8172 17382 8174 17434
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 7956 17360 8252 17380
rect 110 17232 166 17241
rect 110 17167 166 17176
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16998 8524 17070
rect 8588 16998 8616 18158
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 5622 16892 5918 16912
rect 5678 16890 5702 16892
rect 5758 16890 5782 16892
rect 5838 16890 5862 16892
rect 5700 16838 5702 16890
rect 5764 16838 5776 16890
rect 5838 16838 5840 16890
rect 5678 16836 5702 16838
rect 5758 16836 5782 16838
rect 5838 16836 5862 16838
rect 5622 16816 5918 16836
rect 3289 16348 3585 16368
rect 3345 16346 3369 16348
rect 3425 16346 3449 16348
rect 3505 16346 3529 16348
rect 3367 16294 3369 16346
rect 3431 16294 3443 16346
rect 3505 16294 3507 16346
rect 3345 16292 3369 16294
rect 3425 16292 3449 16294
rect 3505 16292 3529 16294
rect 3289 16272 3585 16292
rect 7956 16348 8252 16368
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8034 16294 8036 16346
rect 8098 16294 8110 16346
rect 8172 16294 8174 16346
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 7956 16272 8252 16292
rect 8312 16114 8340 16934
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 5622 15804 5918 15824
rect 5678 15802 5702 15804
rect 5758 15802 5782 15804
rect 5838 15802 5862 15804
rect 5700 15750 5702 15802
rect 5764 15750 5776 15802
rect 5838 15750 5840 15802
rect 5678 15748 5702 15750
rect 5758 15748 5782 15750
rect 5838 15748 5862 15750
rect 5622 15728 5918 15748
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 3289 15260 3585 15280
rect 3345 15258 3369 15260
rect 3425 15258 3449 15260
rect 3505 15258 3529 15260
rect 3367 15206 3369 15258
rect 3431 15206 3443 15258
rect 3505 15206 3507 15258
rect 3345 15204 3369 15206
rect 3425 15204 3449 15206
rect 3505 15204 3529 15206
rect 3289 15184 3585 15204
rect 7392 15162 7420 15574
rect 7852 15502 7880 15914
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7852 14890 7880 15438
rect 7956 15260 8252 15280
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8034 15206 8036 15258
rect 8098 15206 8110 15258
rect 8172 15206 8174 15258
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 7956 15184 8252 15204
rect 8312 15162 8340 15506
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 5622 14716 5918 14736
rect 5678 14714 5702 14716
rect 5758 14714 5782 14716
rect 5838 14714 5862 14716
rect 5700 14662 5702 14714
rect 5764 14662 5776 14714
rect 5838 14662 5840 14714
rect 5678 14660 5702 14662
rect 5758 14660 5782 14662
rect 5838 14660 5862 14662
rect 5622 14640 5918 14660
rect 8496 14482 8524 16934
rect 8576 16516 8628 16522
rect 8680 16504 8708 17478
rect 8628 16476 8708 16504
rect 8576 16458 8628 16464
rect 8588 15638 8616 16458
rect 8772 15638 8800 18702
rect 9416 18426 9444 26182
rect 10152 23474 10180 65962
rect 10289 65852 10585 65872
rect 10345 65850 10369 65852
rect 10425 65850 10449 65852
rect 10505 65850 10529 65852
rect 10367 65798 10369 65850
rect 10431 65798 10443 65850
rect 10505 65798 10507 65850
rect 10345 65796 10369 65798
rect 10425 65796 10449 65798
rect 10505 65796 10529 65798
rect 10289 65776 10585 65796
rect 10289 64764 10585 64784
rect 10345 64762 10369 64764
rect 10425 64762 10449 64764
rect 10505 64762 10529 64764
rect 10367 64710 10369 64762
rect 10431 64710 10443 64762
rect 10505 64710 10507 64762
rect 10345 64708 10369 64710
rect 10425 64708 10449 64710
rect 10505 64708 10529 64710
rect 10289 64688 10585 64708
rect 10289 63676 10585 63696
rect 10345 63674 10369 63676
rect 10425 63674 10449 63676
rect 10505 63674 10529 63676
rect 10367 63622 10369 63674
rect 10431 63622 10443 63674
rect 10505 63622 10507 63674
rect 10345 63620 10369 63622
rect 10425 63620 10449 63622
rect 10505 63620 10529 63622
rect 10289 63600 10585 63620
rect 10289 62588 10585 62608
rect 10345 62586 10369 62588
rect 10425 62586 10449 62588
rect 10505 62586 10529 62588
rect 10367 62534 10369 62586
rect 10431 62534 10443 62586
rect 10505 62534 10507 62586
rect 10345 62532 10369 62534
rect 10425 62532 10449 62534
rect 10505 62532 10529 62534
rect 10289 62512 10585 62532
rect 10289 61500 10585 61520
rect 10345 61498 10369 61500
rect 10425 61498 10449 61500
rect 10505 61498 10529 61500
rect 10367 61446 10369 61498
rect 10431 61446 10443 61498
rect 10505 61446 10507 61498
rect 10345 61444 10369 61446
rect 10425 61444 10449 61446
rect 10505 61444 10529 61446
rect 10289 61424 10585 61444
rect 10289 60412 10585 60432
rect 10345 60410 10369 60412
rect 10425 60410 10449 60412
rect 10505 60410 10529 60412
rect 10367 60358 10369 60410
rect 10431 60358 10443 60410
rect 10505 60358 10507 60410
rect 10345 60356 10369 60358
rect 10425 60356 10449 60358
rect 10505 60356 10529 60358
rect 10289 60336 10585 60356
rect 10289 59324 10585 59344
rect 10345 59322 10369 59324
rect 10425 59322 10449 59324
rect 10505 59322 10529 59324
rect 10367 59270 10369 59322
rect 10431 59270 10443 59322
rect 10505 59270 10507 59322
rect 10345 59268 10369 59270
rect 10425 59268 10449 59270
rect 10505 59268 10529 59270
rect 10289 59248 10585 59268
rect 10289 58236 10585 58256
rect 10345 58234 10369 58236
rect 10425 58234 10449 58236
rect 10505 58234 10529 58236
rect 10367 58182 10369 58234
rect 10431 58182 10443 58234
rect 10505 58182 10507 58234
rect 10345 58180 10369 58182
rect 10425 58180 10449 58182
rect 10505 58180 10529 58182
rect 10289 58160 10585 58180
rect 10289 57148 10585 57168
rect 10345 57146 10369 57148
rect 10425 57146 10449 57148
rect 10505 57146 10529 57148
rect 10367 57094 10369 57146
rect 10431 57094 10443 57146
rect 10505 57094 10507 57146
rect 10345 57092 10369 57094
rect 10425 57092 10449 57094
rect 10505 57092 10529 57094
rect 10289 57072 10585 57092
rect 10289 56060 10585 56080
rect 10345 56058 10369 56060
rect 10425 56058 10449 56060
rect 10505 56058 10529 56060
rect 10367 56006 10369 56058
rect 10431 56006 10443 56058
rect 10505 56006 10507 56058
rect 10345 56004 10369 56006
rect 10425 56004 10449 56006
rect 10505 56004 10529 56006
rect 10289 55984 10585 56004
rect 10289 54972 10585 54992
rect 10345 54970 10369 54972
rect 10425 54970 10449 54972
rect 10505 54970 10529 54972
rect 10367 54918 10369 54970
rect 10431 54918 10443 54970
rect 10505 54918 10507 54970
rect 10345 54916 10369 54918
rect 10425 54916 10449 54918
rect 10505 54916 10529 54918
rect 10289 54896 10585 54916
rect 10289 53884 10585 53904
rect 10345 53882 10369 53884
rect 10425 53882 10449 53884
rect 10505 53882 10529 53884
rect 10367 53830 10369 53882
rect 10431 53830 10443 53882
rect 10505 53830 10507 53882
rect 10345 53828 10369 53830
rect 10425 53828 10449 53830
rect 10505 53828 10529 53830
rect 10289 53808 10585 53828
rect 10289 52796 10585 52816
rect 10345 52794 10369 52796
rect 10425 52794 10449 52796
rect 10505 52794 10529 52796
rect 10367 52742 10369 52794
rect 10431 52742 10443 52794
rect 10505 52742 10507 52794
rect 10345 52740 10369 52742
rect 10425 52740 10449 52742
rect 10505 52740 10529 52742
rect 10289 52720 10585 52740
rect 10289 51708 10585 51728
rect 10345 51706 10369 51708
rect 10425 51706 10449 51708
rect 10505 51706 10529 51708
rect 10367 51654 10369 51706
rect 10431 51654 10443 51706
rect 10505 51654 10507 51706
rect 10345 51652 10369 51654
rect 10425 51652 10449 51654
rect 10505 51652 10529 51654
rect 10289 51632 10585 51652
rect 10289 50620 10585 50640
rect 10345 50618 10369 50620
rect 10425 50618 10449 50620
rect 10505 50618 10529 50620
rect 10367 50566 10369 50618
rect 10431 50566 10443 50618
rect 10505 50566 10507 50618
rect 10345 50564 10369 50566
rect 10425 50564 10449 50566
rect 10505 50564 10529 50566
rect 10289 50544 10585 50564
rect 10289 49532 10585 49552
rect 10345 49530 10369 49532
rect 10425 49530 10449 49532
rect 10505 49530 10529 49532
rect 10367 49478 10369 49530
rect 10431 49478 10443 49530
rect 10505 49478 10507 49530
rect 10345 49476 10369 49478
rect 10425 49476 10449 49478
rect 10505 49476 10529 49478
rect 10289 49456 10585 49476
rect 10289 48444 10585 48464
rect 10345 48442 10369 48444
rect 10425 48442 10449 48444
rect 10505 48442 10529 48444
rect 10367 48390 10369 48442
rect 10431 48390 10443 48442
rect 10505 48390 10507 48442
rect 10345 48388 10369 48390
rect 10425 48388 10449 48390
rect 10505 48388 10529 48390
rect 10289 48368 10585 48388
rect 10289 47356 10585 47376
rect 10345 47354 10369 47356
rect 10425 47354 10449 47356
rect 10505 47354 10529 47356
rect 10367 47302 10369 47354
rect 10431 47302 10443 47354
rect 10505 47302 10507 47354
rect 10345 47300 10369 47302
rect 10425 47300 10449 47302
rect 10505 47300 10529 47302
rect 10289 47280 10585 47300
rect 10289 46268 10585 46288
rect 10345 46266 10369 46268
rect 10425 46266 10449 46268
rect 10505 46266 10529 46268
rect 10367 46214 10369 46266
rect 10431 46214 10443 46266
rect 10505 46214 10507 46266
rect 10345 46212 10369 46214
rect 10425 46212 10449 46214
rect 10505 46212 10529 46214
rect 10289 46192 10585 46212
rect 10289 45180 10585 45200
rect 10345 45178 10369 45180
rect 10425 45178 10449 45180
rect 10505 45178 10529 45180
rect 10367 45126 10369 45178
rect 10431 45126 10443 45178
rect 10505 45126 10507 45178
rect 10345 45124 10369 45126
rect 10425 45124 10449 45126
rect 10505 45124 10529 45126
rect 10289 45104 10585 45124
rect 10782 44296 10838 44305
rect 10782 44231 10838 44240
rect 10289 44092 10585 44112
rect 10345 44090 10369 44092
rect 10425 44090 10449 44092
rect 10505 44090 10529 44092
rect 10367 44038 10369 44090
rect 10431 44038 10443 44090
rect 10505 44038 10507 44090
rect 10345 44036 10369 44038
rect 10425 44036 10449 44038
rect 10505 44036 10529 44038
rect 10289 44016 10585 44036
rect 10289 43004 10585 43024
rect 10345 43002 10369 43004
rect 10425 43002 10449 43004
rect 10505 43002 10529 43004
rect 10367 42950 10369 43002
rect 10431 42950 10443 43002
rect 10505 42950 10507 43002
rect 10345 42948 10369 42950
rect 10425 42948 10449 42950
rect 10505 42948 10529 42950
rect 10289 42928 10585 42948
rect 10289 41916 10585 41936
rect 10345 41914 10369 41916
rect 10425 41914 10449 41916
rect 10505 41914 10529 41916
rect 10367 41862 10369 41914
rect 10431 41862 10443 41914
rect 10505 41862 10507 41914
rect 10345 41860 10369 41862
rect 10425 41860 10449 41862
rect 10505 41860 10529 41862
rect 10289 41840 10585 41860
rect 10289 40828 10585 40848
rect 10345 40826 10369 40828
rect 10425 40826 10449 40828
rect 10505 40826 10529 40828
rect 10367 40774 10369 40826
rect 10431 40774 10443 40826
rect 10505 40774 10507 40826
rect 10345 40772 10369 40774
rect 10425 40772 10449 40774
rect 10505 40772 10529 40774
rect 10289 40752 10585 40772
rect 10796 40186 10824 44231
rect 10784 40180 10836 40186
rect 10784 40122 10836 40128
rect 10289 39740 10585 39760
rect 10345 39738 10369 39740
rect 10425 39738 10449 39740
rect 10505 39738 10529 39740
rect 10367 39686 10369 39738
rect 10431 39686 10443 39738
rect 10505 39686 10507 39738
rect 10345 39684 10369 39686
rect 10425 39684 10449 39686
rect 10505 39684 10529 39686
rect 10289 39664 10585 39684
rect 10289 38652 10585 38672
rect 10345 38650 10369 38652
rect 10425 38650 10449 38652
rect 10505 38650 10529 38652
rect 10367 38598 10369 38650
rect 10431 38598 10443 38650
rect 10505 38598 10507 38650
rect 10345 38596 10369 38598
rect 10425 38596 10449 38598
rect 10505 38596 10529 38598
rect 10289 38576 10585 38596
rect 10289 37564 10585 37584
rect 10345 37562 10369 37564
rect 10425 37562 10449 37564
rect 10505 37562 10529 37564
rect 10367 37510 10369 37562
rect 10431 37510 10443 37562
rect 10505 37510 10507 37562
rect 10345 37508 10369 37510
rect 10425 37508 10449 37510
rect 10505 37508 10529 37510
rect 10289 37488 10585 37508
rect 10289 36476 10585 36496
rect 10345 36474 10369 36476
rect 10425 36474 10449 36476
rect 10505 36474 10529 36476
rect 10367 36422 10369 36474
rect 10431 36422 10443 36474
rect 10505 36422 10507 36474
rect 10345 36420 10369 36422
rect 10425 36420 10449 36422
rect 10505 36420 10529 36422
rect 10289 36400 10585 36420
rect 10289 35388 10585 35408
rect 10345 35386 10369 35388
rect 10425 35386 10449 35388
rect 10505 35386 10529 35388
rect 10367 35334 10369 35386
rect 10431 35334 10443 35386
rect 10505 35334 10507 35386
rect 10345 35332 10369 35334
rect 10425 35332 10449 35334
rect 10505 35332 10529 35334
rect 10289 35312 10585 35332
rect 10289 34300 10585 34320
rect 10345 34298 10369 34300
rect 10425 34298 10449 34300
rect 10505 34298 10529 34300
rect 10367 34246 10369 34298
rect 10431 34246 10443 34298
rect 10505 34246 10507 34298
rect 10345 34244 10369 34246
rect 10425 34244 10449 34246
rect 10505 34244 10529 34246
rect 10289 34224 10585 34244
rect 10289 33212 10585 33232
rect 10345 33210 10369 33212
rect 10425 33210 10449 33212
rect 10505 33210 10529 33212
rect 10367 33158 10369 33210
rect 10431 33158 10443 33210
rect 10505 33158 10507 33210
rect 10345 33156 10369 33158
rect 10425 33156 10449 33158
rect 10505 33156 10529 33158
rect 10289 33136 10585 33156
rect 10289 32124 10585 32144
rect 10345 32122 10369 32124
rect 10425 32122 10449 32124
rect 10505 32122 10529 32124
rect 10367 32070 10369 32122
rect 10431 32070 10443 32122
rect 10505 32070 10507 32122
rect 10345 32068 10369 32070
rect 10425 32068 10449 32070
rect 10505 32068 10529 32070
rect 10289 32048 10585 32068
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10980 31249 11008 31282
rect 10966 31240 11022 31249
rect 10966 31175 11022 31184
rect 10289 31036 10585 31056
rect 10345 31034 10369 31036
rect 10425 31034 10449 31036
rect 10505 31034 10529 31036
rect 10367 30982 10369 31034
rect 10431 30982 10443 31034
rect 10505 30982 10507 31034
rect 10345 30980 10369 30982
rect 10425 30980 10449 30982
rect 10505 30980 10529 30982
rect 10289 30960 10585 30980
rect 10782 30696 10838 30705
rect 10782 30631 10838 30640
rect 10289 29948 10585 29968
rect 10345 29946 10369 29948
rect 10425 29946 10449 29948
rect 10505 29946 10529 29948
rect 10367 29894 10369 29946
rect 10431 29894 10443 29946
rect 10505 29894 10507 29946
rect 10345 29892 10369 29894
rect 10425 29892 10449 29894
rect 10505 29892 10529 29894
rect 10289 29872 10585 29892
rect 10289 28860 10585 28880
rect 10345 28858 10369 28860
rect 10425 28858 10449 28860
rect 10505 28858 10529 28860
rect 10367 28806 10369 28858
rect 10431 28806 10443 28858
rect 10505 28806 10507 28858
rect 10345 28804 10369 28806
rect 10425 28804 10449 28806
rect 10505 28804 10529 28806
rect 10289 28784 10585 28804
rect 10289 27772 10585 27792
rect 10345 27770 10369 27772
rect 10425 27770 10449 27772
rect 10505 27770 10529 27772
rect 10367 27718 10369 27770
rect 10431 27718 10443 27770
rect 10505 27718 10507 27770
rect 10345 27716 10369 27718
rect 10425 27716 10449 27718
rect 10505 27716 10529 27718
rect 10289 27696 10585 27716
rect 10796 27130 10824 30631
rect 10980 27130 11008 31175
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 10968 27124 11020 27130
rect 10968 27066 11020 27072
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10289 26684 10585 26704
rect 10345 26682 10369 26684
rect 10425 26682 10449 26684
rect 10505 26682 10529 26684
rect 10367 26630 10369 26682
rect 10431 26630 10443 26682
rect 10505 26630 10507 26682
rect 10345 26628 10369 26630
rect 10425 26628 10449 26630
rect 10505 26628 10529 26630
rect 10289 26608 10585 26628
rect 10980 26246 11008 26862
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10690 23896 10746 23905
rect 10690 23831 10746 23840
rect 9968 23446 10180 23474
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 15910 8984 16390
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 3289 14172 3585 14192
rect 3345 14170 3369 14172
rect 3425 14170 3449 14172
rect 3505 14170 3529 14172
rect 3367 14118 3369 14170
rect 3431 14118 3443 14170
rect 3505 14118 3507 14170
rect 3345 14116 3369 14118
rect 3425 14116 3449 14118
rect 3505 14116 3529 14118
rect 3289 14096 3585 14116
rect 7852 13734 7880 14418
rect 8588 14346 8616 15574
rect 8956 15366 8984 15846
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 14890 8984 15302
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8772 14414 8800 14758
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 7956 14172 8252 14192
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8034 14118 8036 14170
rect 8098 14118 8110 14170
rect 8172 14118 8174 14170
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 7956 14096 8252 14116
rect 8772 13734 8800 14350
rect 8956 13870 8984 14826
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 5622 13628 5918 13648
rect 5678 13626 5702 13628
rect 5758 13626 5782 13628
rect 5838 13626 5862 13628
rect 5700 13574 5702 13626
rect 5764 13574 5776 13626
rect 5838 13574 5840 13626
rect 5678 13572 5702 13574
rect 5758 13572 5782 13574
rect 5838 13572 5862 13574
rect 5622 13552 5918 13572
rect 3289 13084 3585 13104
rect 3345 13082 3369 13084
rect 3425 13082 3449 13084
rect 3505 13082 3529 13084
rect 3367 13030 3369 13082
rect 3431 13030 3443 13082
rect 3505 13030 3507 13082
rect 3345 13028 3369 13030
rect 3425 13028 3449 13030
rect 3505 13028 3529 13030
rect 3289 13008 3585 13028
rect 1308 12640 1360 12646
rect 1308 12582 1360 12588
rect 110 6896 166 6905
rect 110 6831 166 6840
rect 124 5681 152 6831
rect 110 5672 166 5681
rect 110 5607 166 5616
rect 1122 82 1178 480
rect 1320 82 1348 12582
rect 5622 12540 5918 12560
rect 5678 12538 5702 12540
rect 5758 12538 5782 12540
rect 5838 12538 5862 12540
rect 5700 12486 5702 12538
rect 5764 12486 5776 12538
rect 5838 12486 5840 12538
rect 5678 12484 5702 12486
rect 5758 12484 5782 12486
rect 5838 12484 5862 12486
rect 5622 12464 5918 12484
rect 3289 11996 3585 12016
rect 3345 11994 3369 11996
rect 3425 11994 3449 11996
rect 3505 11994 3529 11996
rect 3367 11942 3369 11994
rect 3431 11942 3443 11994
rect 3505 11942 3507 11994
rect 3345 11940 3369 11942
rect 3425 11940 3449 11942
rect 3505 11940 3529 11942
rect 3289 11920 3585 11940
rect 5622 11452 5918 11472
rect 5678 11450 5702 11452
rect 5758 11450 5782 11452
rect 5838 11450 5862 11452
rect 5700 11398 5702 11450
rect 5764 11398 5776 11450
rect 5838 11398 5840 11450
rect 5678 11396 5702 11398
rect 5758 11396 5782 11398
rect 5838 11396 5862 11398
rect 5622 11376 5918 11396
rect 3289 10908 3585 10928
rect 3345 10906 3369 10908
rect 3425 10906 3449 10908
rect 3505 10906 3529 10908
rect 3367 10854 3369 10906
rect 3431 10854 3443 10906
rect 3505 10854 3507 10906
rect 3345 10852 3369 10854
rect 3425 10852 3449 10854
rect 3505 10852 3529 10854
rect 3289 10832 3585 10852
rect 5622 10364 5918 10384
rect 5678 10362 5702 10364
rect 5758 10362 5782 10364
rect 5838 10362 5862 10364
rect 5700 10310 5702 10362
rect 5764 10310 5776 10362
rect 5838 10310 5840 10362
rect 5678 10308 5702 10310
rect 5758 10308 5782 10310
rect 5838 10308 5862 10310
rect 5622 10288 5918 10308
rect 3289 9820 3585 9840
rect 3345 9818 3369 9820
rect 3425 9818 3449 9820
rect 3505 9818 3529 9820
rect 3367 9766 3369 9818
rect 3431 9766 3443 9818
rect 3505 9766 3507 9818
rect 3345 9764 3369 9766
rect 3425 9764 3449 9766
rect 3505 9764 3529 9766
rect 3289 9744 3585 9764
rect 5622 9276 5918 9296
rect 5678 9274 5702 9276
rect 5758 9274 5782 9276
rect 5838 9274 5862 9276
rect 5700 9222 5702 9274
rect 5764 9222 5776 9274
rect 5838 9222 5840 9274
rect 5678 9220 5702 9222
rect 5758 9220 5782 9222
rect 5838 9220 5862 9222
rect 5622 9200 5918 9220
rect 3289 8732 3585 8752
rect 3345 8730 3369 8732
rect 3425 8730 3449 8732
rect 3505 8730 3529 8732
rect 3367 8678 3369 8730
rect 3431 8678 3443 8730
rect 3505 8678 3507 8730
rect 3345 8676 3369 8678
rect 3425 8676 3449 8678
rect 3505 8676 3529 8678
rect 3289 8656 3585 8676
rect 5622 8188 5918 8208
rect 5678 8186 5702 8188
rect 5758 8186 5782 8188
rect 5838 8186 5862 8188
rect 5700 8134 5702 8186
rect 5764 8134 5776 8186
rect 5838 8134 5840 8186
rect 5678 8132 5702 8134
rect 5758 8132 5782 8134
rect 5838 8132 5862 8134
rect 5622 8112 5918 8132
rect 3289 7644 3585 7664
rect 3345 7642 3369 7644
rect 3425 7642 3449 7644
rect 3505 7642 3529 7644
rect 3367 7590 3369 7642
rect 3431 7590 3443 7642
rect 3505 7590 3507 7642
rect 3345 7588 3369 7590
rect 3425 7588 3449 7590
rect 3505 7588 3529 7590
rect 3289 7568 3585 7588
rect 5622 7100 5918 7120
rect 5678 7098 5702 7100
rect 5758 7098 5782 7100
rect 5838 7098 5862 7100
rect 5700 7046 5702 7098
rect 5764 7046 5776 7098
rect 5838 7046 5840 7098
rect 5678 7044 5702 7046
rect 5758 7044 5782 7046
rect 5838 7044 5862 7046
rect 5622 7024 5918 7044
rect 3289 6556 3585 6576
rect 3345 6554 3369 6556
rect 3425 6554 3449 6556
rect 3505 6554 3529 6556
rect 3367 6502 3369 6554
rect 3431 6502 3443 6554
rect 3505 6502 3507 6554
rect 3345 6500 3369 6502
rect 3425 6500 3449 6502
rect 3505 6500 3529 6502
rect 3289 6480 3585 6500
rect 5622 6012 5918 6032
rect 5678 6010 5702 6012
rect 5758 6010 5782 6012
rect 5838 6010 5862 6012
rect 5700 5958 5702 6010
rect 5764 5958 5776 6010
rect 5838 5958 5840 6010
rect 5678 5956 5702 5958
rect 5758 5956 5782 5958
rect 5838 5956 5862 5958
rect 5622 5936 5918 5956
rect 3289 5468 3585 5488
rect 3345 5466 3369 5468
rect 3425 5466 3449 5468
rect 3505 5466 3529 5468
rect 3367 5414 3369 5466
rect 3431 5414 3443 5466
rect 3505 5414 3507 5466
rect 3345 5412 3369 5414
rect 3425 5412 3449 5414
rect 3505 5412 3529 5414
rect 3289 5392 3585 5412
rect 5622 4924 5918 4944
rect 5678 4922 5702 4924
rect 5758 4922 5782 4924
rect 5838 4922 5862 4924
rect 5700 4870 5702 4922
rect 5764 4870 5776 4922
rect 5838 4870 5840 4922
rect 5678 4868 5702 4870
rect 5758 4868 5782 4870
rect 5838 4868 5862 4870
rect 5622 4848 5918 4868
rect 3289 4380 3585 4400
rect 3345 4378 3369 4380
rect 3425 4378 3449 4380
rect 3505 4378 3529 4380
rect 3367 4326 3369 4378
rect 3431 4326 3443 4378
rect 3505 4326 3507 4378
rect 3345 4324 3369 4326
rect 3425 4324 3449 4326
rect 3505 4324 3529 4326
rect 3289 4304 3585 4324
rect 5622 3836 5918 3856
rect 5678 3834 5702 3836
rect 5758 3834 5782 3836
rect 5838 3834 5862 3836
rect 5700 3782 5702 3834
rect 5764 3782 5776 3834
rect 5838 3782 5840 3834
rect 5678 3780 5702 3782
rect 5758 3780 5782 3782
rect 5838 3780 5862 3782
rect 5622 3760 5918 3780
rect 3289 3292 3585 3312
rect 3345 3290 3369 3292
rect 3425 3290 3449 3292
rect 3505 3290 3529 3292
rect 3367 3238 3369 3290
rect 3431 3238 3443 3290
rect 3505 3238 3507 3290
rect 3345 3236 3369 3238
rect 3425 3236 3449 3238
rect 3505 3236 3529 3238
rect 3289 3216 3585 3236
rect 7852 2854 7880 13670
rect 7956 13084 8252 13104
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8034 13030 8036 13082
rect 8098 13030 8110 13082
rect 8172 13030 8174 13082
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 7956 13008 8252 13028
rect 8772 12102 8800 13670
rect 9048 12714 9076 15982
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9232 14550 9260 15098
rect 9692 15026 9720 18022
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9784 16046 9812 17070
rect 9876 16504 9904 17070
rect 9968 16794 9996 23446
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10060 18630 10088 19246
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9956 16516 10008 16522
rect 9876 16476 9956 16504
rect 9956 16458 10008 16464
rect 9968 16046 9996 16458
rect 10060 16182 10088 18566
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 17338 10180 17614
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9784 15502 9812 15982
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9324 14890 9352 14962
rect 9772 14952 9824 14958
rect 9876 14940 9904 15574
rect 9968 15162 9996 15642
rect 10152 15638 10180 17274
rect 10704 17270 10732 23831
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18902 10824 19110
rect 10784 18896 10836 18902
rect 10784 18838 10836 18844
rect 10796 18086 10824 18838
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17814 10824 18022
rect 11072 17882 11100 94250
rect 11518 85232 11574 85241
rect 11518 85167 11520 85176
rect 11572 85167 11574 85176
rect 11520 85138 11572 85144
rect 11150 85096 11206 85105
rect 11150 85031 11206 85040
rect 11164 80850 11192 85031
rect 11532 84794 11560 85138
rect 11520 84788 11572 84794
rect 11520 84730 11572 84736
rect 11796 84788 11848 84794
rect 11796 84730 11848 84736
rect 11808 80986 11836 84730
rect 11796 80980 11848 80986
rect 11796 80922 11848 80928
rect 11152 80844 11204 80850
rect 11152 80786 11204 80792
rect 11164 80442 11192 80786
rect 11336 80776 11388 80782
rect 11336 80718 11388 80724
rect 11152 80436 11204 80442
rect 11152 80378 11204 80384
rect 11348 80102 11376 80718
rect 11152 80096 11204 80102
rect 11152 80038 11204 80044
rect 11336 80096 11388 80102
rect 11336 80038 11388 80044
rect 11164 18426 11192 80038
rect 11242 71632 11298 71641
rect 11242 71567 11298 71576
rect 11256 71534 11284 71567
rect 11244 71528 11296 71534
rect 11796 71528 11848 71534
rect 11244 71470 11296 71476
rect 11426 71496 11482 71505
rect 11796 71470 11848 71476
rect 11426 71431 11482 71440
rect 11440 66706 11468 71431
rect 11808 66842 11836 71470
rect 11796 66836 11848 66842
rect 11796 66778 11848 66784
rect 11428 66700 11480 66706
rect 11428 66642 11480 66648
rect 11336 66632 11388 66638
rect 11336 66574 11388 66580
rect 11348 66026 11376 66574
rect 11440 66298 11468 66642
rect 11428 66292 11480 66298
rect 11428 66234 11480 66240
rect 11336 66020 11388 66026
rect 11336 65962 11388 65968
rect 11426 64696 11482 64705
rect 11426 64631 11482 64640
rect 11440 58682 11468 64631
rect 11428 58676 11480 58682
rect 11428 58618 11480 58624
rect 11242 58576 11298 58585
rect 11242 58511 11298 58520
rect 11256 58478 11284 58511
rect 11244 58472 11296 58478
rect 11244 58414 11296 58420
rect 11796 58472 11848 58478
rect 11796 58414 11848 58420
rect 11426 57896 11482 57905
rect 11426 57831 11482 57840
rect 11440 53650 11468 57831
rect 11808 53786 11836 58414
rect 11796 53780 11848 53786
rect 11796 53722 11848 53728
rect 11428 53644 11480 53650
rect 11428 53586 11480 53592
rect 11440 53242 11468 53586
rect 11612 53576 11664 53582
rect 11612 53518 11664 53524
rect 11428 53236 11480 53242
rect 11428 53178 11480 53184
rect 11624 52902 11652 53518
rect 11612 52896 11664 52902
rect 11612 52838 11664 52844
rect 11520 44940 11572 44946
rect 11520 44882 11572 44888
rect 11532 44849 11560 44882
rect 11518 44840 11574 44849
rect 11518 44775 11574 44784
rect 11532 44538 11560 44775
rect 11520 44532 11572 44538
rect 11520 44474 11572 44480
rect 11532 40186 11560 44474
rect 11520 40180 11572 40186
rect 11520 40122 11572 40128
rect 11244 39976 11296 39982
rect 11244 39918 11296 39924
rect 11256 39302 11284 39918
rect 11244 39296 11296 39302
rect 11244 39238 11296 39244
rect 11256 19514 11284 39238
rect 11426 37496 11482 37505
rect 11426 37431 11482 37440
rect 11440 31482 11468 37431
rect 11428 31476 11480 31482
rect 11428 31418 11480 31424
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11624 18970 11652 52838
rect 11702 51096 11758 51105
rect 11702 51031 11758 51040
rect 11716 45082 11744 51031
rect 11704 45076 11756 45082
rect 11704 45018 11756 45024
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11808 18426 11836 18702
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10796 16998 10824 17750
rect 11242 17232 11298 17241
rect 11242 17167 11298 17176
rect 11256 17134 11284 17167
rect 11244 17128 11296 17134
rect 11150 17096 11206 17105
rect 11244 17070 11296 17076
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11150 17031 11206 17040
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10796 16726 10824 16934
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10704 16250 10732 16526
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10692 15904 10744 15910
rect 10796 15892 10824 16662
rect 10744 15864 10824 15892
rect 10692 15846 10744 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15688 10732 15846
rect 10612 15660 10732 15688
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9824 14912 9904 14940
rect 9772 14894 9824 14900
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9324 14618 9352 14826
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 7956 11996 8252 12016
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8034 11942 8036 11994
rect 8098 11942 8110 11994
rect 8172 11942 8174 11994
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 7956 11920 8252 11940
rect 8772 11694 8800 12038
rect 9048 11694 9076 12650
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 7956 10908 8252 10928
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8034 10854 8036 10906
rect 8098 10854 8110 10906
rect 8172 10854 8174 10906
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 7956 10832 8252 10852
rect 7956 9820 8252 9840
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8034 9766 8036 9818
rect 8098 9766 8110 9818
rect 8172 9766 8174 9818
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 7956 9744 8252 9764
rect 7956 8732 8252 8752
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8034 8678 8036 8730
rect 8098 8678 8110 8730
rect 8172 8678 8174 8730
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 7956 8656 8252 8676
rect 7956 7644 8252 7664
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8034 7590 8036 7642
rect 8098 7590 8110 7642
rect 8172 7590 8174 7642
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 7956 7568 8252 7588
rect 7956 6556 8252 6576
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8034 6502 8036 6554
rect 8098 6502 8110 6554
rect 8172 6502 8174 6554
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 7956 6480 8252 6500
rect 7956 5468 8252 5488
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8034 5414 8036 5466
rect 8098 5414 8110 5466
rect 8172 5414 8174 5466
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 7956 5392 8252 5412
rect 7956 4380 8252 4400
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8034 4326 8036 4378
rect 8098 4326 8110 4378
rect 8172 4326 8174 4378
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 7956 4304 8252 4324
rect 7956 3292 8252 3312
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8034 3238 8036 3290
rect 8098 3238 8110 3290
rect 8172 3238 8174 3290
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 7956 3216 8252 3236
rect 9048 2990 9076 11630
rect 9232 4078 9260 14486
rect 9312 14476 9364 14482
rect 9416 14464 9444 14758
rect 9364 14436 9444 14464
rect 9312 14418 9364 14424
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9416 11694 9444 13806
rect 9600 12782 9628 14826
rect 9784 14482 9812 14894
rect 9968 14822 9996 15098
rect 9956 14816 10008 14822
rect 10612 14804 10640 15660
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10704 15366 10732 15506
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 14958 10732 15302
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10784 14816 10836 14822
rect 10612 14776 10732 14804
rect 9956 14758 10008 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 13734 9812 14418
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10060 13734 10088 13806
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9784 11762 9812 13670
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11014 9444 11630
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 4214 9444 10950
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9416 3738 9444 4150
rect 9508 3738 9536 10406
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9416 2990 9444 3674
rect 9784 2990 9812 11698
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 11218 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11354 10732 14776
rect 10784 14758 10836 14764
rect 10796 14550 10824 14758
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10888 14414 10916 14826
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 11164 13394 11192 17031
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11256 15026 11284 16186
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11808 13530 11836 17070
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11164 12986 11192 13330
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12646 11284 13262
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 11354 11284 12582
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10810 10180 11154
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10704 10470 10732 11290
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 11426 10296 11482 10305
rect 11426 10231 11482 10240
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 11256 4078 11284 5607
rect 11440 4282 11468 10231
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 5622 2748 5918 2768
rect 5678 2746 5702 2748
rect 5758 2746 5782 2748
rect 5838 2746 5862 2748
rect 5700 2694 5702 2746
rect 5764 2694 5776 2746
rect 5838 2694 5840 2746
rect 5678 2692 5702 2694
rect 5758 2692 5782 2694
rect 5838 2692 5862 2694
rect 5622 2672 5918 2692
rect 3289 2204 3585 2224
rect 3345 2202 3369 2204
rect 3425 2202 3449 2204
rect 3505 2202 3529 2204
rect 3367 2150 3369 2202
rect 3431 2150 3443 2202
rect 3505 2150 3507 2202
rect 3345 2148 3369 2150
rect 3425 2148 3449 2150
rect 3505 2148 3529 2150
rect 3289 2128 3585 2148
rect 1122 54 1348 82
rect 1122 0 1178 54
rect 3422 0 3478 480
rect 5722 82 5778 480
rect 6012 82 6040 2790
rect 9784 2310 9812 2926
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 7956 2204 8252 2224
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8034 2150 8036 2202
rect 8098 2150 8110 2202
rect 8172 2150 8174 2202
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 7956 2128 8252 2148
rect 5722 54 6040 82
rect 8114 82 8170 480
rect 8404 82 8432 2246
rect 8114 54 8432 82
rect 10060 82 10088 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10152 3058 10180 3470
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10704 2854 10732 3674
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10980 2650 11008 3431
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10980 2446 11008 2586
rect 11256 2514 11284 3334
rect 11716 2650 11744 3878
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10414 82 10470 480
rect 10060 54 10470 82
rect 12360 82 12388 2790
rect 12714 82 12770 480
rect 12360 54 12770 82
rect 5722 0 5778 54
rect 8114 0 8170 54
rect 10414 0 10470 54
rect 12714 0 12770 54
<< via2 >>
rect 3289 106650 3345 106652
rect 3369 106650 3425 106652
rect 3449 106650 3505 106652
rect 3529 106650 3585 106652
rect 3289 106598 3315 106650
rect 3315 106598 3345 106650
rect 3369 106598 3379 106650
rect 3379 106598 3425 106650
rect 3449 106598 3495 106650
rect 3495 106598 3505 106650
rect 3529 106598 3559 106650
rect 3559 106598 3585 106650
rect 3289 106596 3345 106598
rect 3369 106596 3425 106598
rect 3449 106596 3505 106598
rect 3529 106596 3585 106598
rect 7956 106650 8012 106652
rect 8036 106650 8092 106652
rect 8116 106650 8172 106652
rect 8196 106650 8252 106652
rect 7956 106598 7982 106650
rect 7982 106598 8012 106650
rect 8036 106598 8046 106650
rect 8046 106598 8092 106650
rect 8116 106598 8162 106650
rect 8162 106598 8172 106650
rect 8196 106598 8226 106650
rect 8226 106598 8252 106650
rect 7956 106596 8012 106598
rect 8036 106596 8092 106598
rect 8116 106596 8172 106598
rect 8196 106596 8252 106598
rect 5622 106106 5678 106108
rect 5702 106106 5758 106108
rect 5782 106106 5838 106108
rect 5862 106106 5918 106108
rect 5622 106054 5648 106106
rect 5648 106054 5678 106106
rect 5702 106054 5712 106106
rect 5712 106054 5758 106106
rect 5782 106054 5828 106106
rect 5828 106054 5838 106106
rect 5862 106054 5892 106106
rect 5892 106054 5918 106106
rect 5622 106052 5678 106054
rect 5702 106052 5758 106054
rect 5782 106052 5838 106054
rect 5862 106052 5918 106054
rect 10289 106106 10345 106108
rect 10369 106106 10425 106108
rect 10449 106106 10505 106108
rect 10529 106106 10585 106108
rect 10289 106054 10315 106106
rect 10315 106054 10345 106106
rect 10369 106054 10379 106106
rect 10379 106054 10425 106106
rect 10449 106054 10495 106106
rect 10495 106054 10505 106106
rect 10529 106054 10559 106106
rect 10559 106054 10585 106106
rect 10289 106052 10345 106054
rect 10369 106052 10425 106054
rect 10449 106052 10505 106054
rect 10529 106052 10585 106054
rect 3289 105562 3345 105564
rect 3369 105562 3425 105564
rect 3449 105562 3505 105564
rect 3529 105562 3585 105564
rect 3289 105510 3315 105562
rect 3315 105510 3345 105562
rect 3369 105510 3379 105562
rect 3379 105510 3425 105562
rect 3449 105510 3495 105562
rect 3495 105510 3505 105562
rect 3529 105510 3559 105562
rect 3559 105510 3585 105562
rect 3289 105508 3345 105510
rect 3369 105508 3425 105510
rect 3449 105508 3505 105510
rect 3529 105508 3585 105510
rect 7956 105562 8012 105564
rect 8036 105562 8092 105564
rect 8116 105562 8172 105564
rect 8196 105562 8252 105564
rect 7956 105510 7982 105562
rect 7982 105510 8012 105562
rect 8036 105510 8046 105562
rect 8046 105510 8092 105562
rect 8116 105510 8162 105562
rect 8162 105510 8172 105562
rect 8196 105510 8226 105562
rect 8226 105510 8252 105562
rect 7956 105508 8012 105510
rect 8036 105508 8092 105510
rect 8116 105508 8172 105510
rect 8196 105508 8252 105510
rect 11426 105440 11482 105496
rect 5622 105018 5678 105020
rect 5702 105018 5758 105020
rect 5782 105018 5838 105020
rect 5862 105018 5918 105020
rect 5622 104966 5648 105018
rect 5648 104966 5678 105018
rect 5702 104966 5712 105018
rect 5712 104966 5758 105018
rect 5782 104966 5828 105018
rect 5828 104966 5838 105018
rect 5862 104966 5892 105018
rect 5892 104966 5918 105018
rect 5622 104964 5678 104966
rect 5702 104964 5758 104966
rect 5782 104964 5838 104966
rect 5862 104964 5918 104966
rect 10289 105018 10345 105020
rect 10369 105018 10425 105020
rect 10449 105018 10505 105020
rect 10529 105018 10585 105020
rect 10289 104966 10315 105018
rect 10315 104966 10345 105018
rect 10369 104966 10379 105018
rect 10379 104966 10425 105018
rect 10449 104966 10495 105018
rect 10495 104966 10505 105018
rect 10529 104966 10559 105018
rect 10559 104966 10585 105018
rect 10289 104964 10345 104966
rect 10369 104964 10425 104966
rect 10449 104964 10505 104966
rect 10529 104964 10585 104966
rect 3289 104474 3345 104476
rect 3369 104474 3425 104476
rect 3449 104474 3505 104476
rect 3529 104474 3585 104476
rect 3289 104422 3315 104474
rect 3315 104422 3345 104474
rect 3369 104422 3379 104474
rect 3379 104422 3425 104474
rect 3449 104422 3495 104474
rect 3495 104422 3505 104474
rect 3529 104422 3559 104474
rect 3559 104422 3585 104474
rect 3289 104420 3345 104422
rect 3369 104420 3425 104422
rect 3449 104420 3505 104422
rect 3529 104420 3585 104422
rect 7956 104474 8012 104476
rect 8036 104474 8092 104476
rect 8116 104474 8172 104476
rect 8196 104474 8252 104476
rect 7956 104422 7982 104474
rect 7982 104422 8012 104474
rect 8036 104422 8046 104474
rect 8046 104422 8092 104474
rect 8116 104422 8162 104474
rect 8162 104422 8172 104474
rect 8196 104422 8226 104474
rect 8226 104422 8252 104474
rect 7956 104420 8012 104422
rect 8036 104420 8092 104422
rect 8116 104420 8172 104422
rect 8196 104420 8252 104422
rect 5622 103930 5678 103932
rect 5702 103930 5758 103932
rect 5782 103930 5838 103932
rect 5862 103930 5918 103932
rect 5622 103878 5648 103930
rect 5648 103878 5678 103930
rect 5702 103878 5712 103930
rect 5712 103878 5758 103930
rect 5782 103878 5828 103930
rect 5828 103878 5838 103930
rect 5862 103878 5892 103930
rect 5892 103878 5918 103930
rect 5622 103876 5678 103878
rect 5702 103876 5758 103878
rect 5782 103876 5838 103878
rect 5862 103876 5918 103878
rect 10289 103930 10345 103932
rect 10369 103930 10425 103932
rect 10449 103930 10505 103932
rect 10529 103930 10585 103932
rect 10289 103878 10315 103930
rect 10315 103878 10345 103930
rect 10369 103878 10379 103930
rect 10379 103878 10425 103930
rect 10449 103878 10495 103930
rect 10495 103878 10505 103930
rect 10529 103878 10559 103930
rect 10559 103878 10585 103930
rect 10289 103876 10345 103878
rect 10369 103876 10425 103878
rect 10449 103876 10505 103878
rect 10529 103876 10585 103878
rect 3289 103386 3345 103388
rect 3369 103386 3425 103388
rect 3449 103386 3505 103388
rect 3529 103386 3585 103388
rect 3289 103334 3315 103386
rect 3315 103334 3345 103386
rect 3369 103334 3379 103386
rect 3379 103334 3425 103386
rect 3449 103334 3495 103386
rect 3495 103334 3505 103386
rect 3529 103334 3559 103386
rect 3559 103334 3585 103386
rect 3289 103332 3345 103334
rect 3369 103332 3425 103334
rect 3449 103332 3505 103334
rect 3529 103332 3585 103334
rect 7956 103386 8012 103388
rect 8036 103386 8092 103388
rect 8116 103386 8172 103388
rect 8196 103386 8252 103388
rect 7956 103334 7982 103386
rect 7982 103334 8012 103386
rect 8036 103334 8046 103386
rect 8046 103334 8092 103386
rect 8116 103334 8162 103386
rect 8162 103334 8172 103386
rect 8196 103334 8226 103386
rect 8226 103334 8252 103386
rect 7956 103332 8012 103334
rect 8036 103332 8092 103334
rect 8116 103332 8172 103334
rect 8196 103332 8252 103334
rect 5622 102842 5678 102844
rect 5702 102842 5758 102844
rect 5782 102842 5838 102844
rect 5862 102842 5918 102844
rect 5622 102790 5648 102842
rect 5648 102790 5678 102842
rect 5702 102790 5712 102842
rect 5712 102790 5758 102842
rect 5782 102790 5828 102842
rect 5828 102790 5838 102842
rect 5862 102790 5892 102842
rect 5892 102790 5918 102842
rect 5622 102788 5678 102790
rect 5702 102788 5758 102790
rect 5782 102788 5838 102790
rect 5862 102788 5918 102790
rect 10289 102842 10345 102844
rect 10369 102842 10425 102844
rect 10449 102842 10505 102844
rect 10529 102842 10585 102844
rect 10289 102790 10315 102842
rect 10315 102790 10345 102842
rect 10369 102790 10379 102842
rect 10379 102790 10425 102842
rect 10449 102790 10495 102842
rect 10495 102790 10505 102842
rect 10529 102790 10559 102842
rect 10559 102790 10585 102842
rect 10289 102788 10345 102790
rect 10369 102788 10425 102790
rect 10449 102788 10505 102790
rect 10529 102788 10585 102790
rect 3289 102298 3345 102300
rect 3369 102298 3425 102300
rect 3449 102298 3505 102300
rect 3529 102298 3585 102300
rect 3289 102246 3315 102298
rect 3315 102246 3345 102298
rect 3369 102246 3379 102298
rect 3379 102246 3425 102298
rect 3449 102246 3495 102298
rect 3495 102246 3505 102298
rect 3529 102246 3559 102298
rect 3559 102246 3585 102298
rect 3289 102244 3345 102246
rect 3369 102244 3425 102246
rect 3449 102244 3505 102246
rect 3529 102244 3585 102246
rect 7956 102298 8012 102300
rect 8036 102298 8092 102300
rect 8116 102298 8172 102300
rect 8196 102298 8252 102300
rect 7956 102246 7982 102298
rect 7982 102246 8012 102298
rect 8036 102246 8046 102298
rect 8046 102246 8092 102298
rect 8116 102246 8162 102298
rect 8162 102246 8172 102298
rect 8196 102246 8226 102298
rect 8226 102246 8252 102298
rect 7956 102244 8012 102246
rect 8036 102244 8092 102246
rect 8116 102244 8172 102246
rect 8196 102244 8252 102246
rect 110 102040 166 102096
rect 5622 101754 5678 101756
rect 5702 101754 5758 101756
rect 5782 101754 5838 101756
rect 5862 101754 5918 101756
rect 5622 101702 5648 101754
rect 5648 101702 5678 101754
rect 5702 101702 5712 101754
rect 5712 101702 5758 101754
rect 5782 101702 5828 101754
rect 5828 101702 5838 101754
rect 5862 101702 5892 101754
rect 5892 101702 5918 101754
rect 5622 101700 5678 101702
rect 5702 101700 5758 101702
rect 5782 101700 5838 101702
rect 5862 101700 5918 101702
rect 10289 101754 10345 101756
rect 10369 101754 10425 101756
rect 10449 101754 10505 101756
rect 10529 101754 10585 101756
rect 10289 101702 10315 101754
rect 10315 101702 10345 101754
rect 10369 101702 10379 101754
rect 10379 101702 10425 101754
rect 10449 101702 10495 101754
rect 10495 101702 10505 101754
rect 10529 101702 10559 101754
rect 10559 101702 10585 101754
rect 10289 101700 10345 101702
rect 10369 101700 10425 101702
rect 10449 101700 10505 101702
rect 10529 101700 10585 101702
rect 3289 101210 3345 101212
rect 3369 101210 3425 101212
rect 3449 101210 3505 101212
rect 3529 101210 3585 101212
rect 3289 101158 3315 101210
rect 3315 101158 3345 101210
rect 3369 101158 3379 101210
rect 3379 101158 3425 101210
rect 3449 101158 3495 101210
rect 3495 101158 3505 101210
rect 3529 101158 3559 101210
rect 3559 101158 3585 101210
rect 3289 101156 3345 101158
rect 3369 101156 3425 101158
rect 3449 101156 3505 101158
rect 3529 101156 3585 101158
rect 7956 101210 8012 101212
rect 8036 101210 8092 101212
rect 8116 101210 8172 101212
rect 8196 101210 8252 101212
rect 7956 101158 7982 101210
rect 7982 101158 8012 101210
rect 8036 101158 8046 101210
rect 8046 101158 8092 101210
rect 8116 101158 8162 101210
rect 8162 101158 8172 101210
rect 8196 101158 8226 101210
rect 8226 101158 8252 101210
rect 7956 101156 8012 101158
rect 8036 101156 8092 101158
rect 8116 101156 8172 101158
rect 8196 101156 8252 101158
rect 5622 100666 5678 100668
rect 5702 100666 5758 100668
rect 5782 100666 5838 100668
rect 5862 100666 5918 100668
rect 5622 100614 5648 100666
rect 5648 100614 5678 100666
rect 5702 100614 5712 100666
rect 5712 100614 5758 100666
rect 5782 100614 5828 100666
rect 5828 100614 5838 100666
rect 5862 100614 5892 100666
rect 5892 100614 5918 100666
rect 5622 100612 5678 100614
rect 5702 100612 5758 100614
rect 5782 100612 5838 100614
rect 5862 100612 5918 100614
rect 10289 100666 10345 100668
rect 10369 100666 10425 100668
rect 10449 100666 10505 100668
rect 10529 100666 10585 100668
rect 10289 100614 10315 100666
rect 10315 100614 10345 100666
rect 10369 100614 10379 100666
rect 10379 100614 10425 100666
rect 10449 100614 10495 100666
rect 10495 100614 10505 100666
rect 10529 100614 10559 100666
rect 10559 100614 10585 100666
rect 10289 100612 10345 100614
rect 10369 100612 10425 100614
rect 10449 100612 10505 100614
rect 10529 100612 10585 100614
rect 3289 100122 3345 100124
rect 3369 100122 3425 100124
rect 3449 100122 3505 100124
rect 3529 100122 3585 100124
rect 3289 100070 3315 100122
rect 3315 100070 3345 100122
rect 3369 100070 3379 100122
rect 3379 100070 3425 100122
rect 3449 100070 3495 100122
rect 3495 100070 3505 100122
rect 3529 100070 3559 100122
rect 3559 100070 3585 100122
rect 3289 100068 3345 100070
rect 3369 100068 3425 100070
rect 3449 100068 3505 100070
rect 3529 100068 3585 100070
rect 7956 100122 8012 100124
rect 8036 100122 8092 100124
rect 8116 100122 8172 100124
rect 8196 100122 8252 100124
rect 7956 100070 7982 100122
rect 7982 100070 8012 100122
rect 8036 100070 8046 100122
rect 8046 100070 8092 100122
rect 8116 100070 8162 100122
rect 8162 100070 8172 100122
rect 8196 100070 8226 100122
rect 8226 100070 8252 100122
rect 7956 100068 8012 100070
rect 8036 100068 8092 100070
rect 8116 100068 8172 100070
rect 8196 100068 8252 100070
rect 5622 99578 5678 99580
rect 5702 99578 5758 99580
rect 5782 99578 5838 99580
rect 5862 99578 5918 99580
rect 5622 99526 5648 99578
rect 5648 99526 5678 99578
rect 5702 99526 5712 99578
rect 5712 99526 5758 99578
rect 5782 99526 5828 99578
rect 5828 99526 5838 99578
rect 5862 99526 5892 99578
rect 5892 99526 5918 99578
rect 5622 99524 5678 99526
rect 5702 99524 5758 99526
rect 5782 99524 5838 99526
rect 5862 99524 5918 99526
rect 10289 99578 10345 99580
rect 10369 99578 10425 99580
rect 10449 99578 10505 99580
rect 10529 99578 10585 99580
rect 10289 99526 10315 99578
rect 10315 99526 10345 99578
rect 10369 99526 10379 99578
rect 10379 99526 10425 99578
rect 10449 99526 10495 99578
rect 10495 99526 10505 99578
rect 10529 99526 10559 99578
rect 10559 99526 10585 99578
rect 10289 99524 10345 99526
rect 10369 99524 10425 99526
rect 10449 99524 10505 99526
rect 10529 99524 10585 99526
rect 3289 99034 3345 99036
rect 3369 99034 3425 99036
rect 3449 99034 3505 99036
rect 3529 99034 3585 99036
rect 3289 98982 3315 99034
rect 3315 98982 3345 99034
rect 3369 98982 3379 99034
rect 3379 98982 3425 99034
rect 3449 98982 3495 99034
rect 3495 98982 3505 99034
rect 3529 98982 3559 99034
rect 3559 98982 3585 99034
rect 3289 98980 3345 98982
rect 3369 98980 3425 98982
rect 3449 98980 3505 98982
rect 3529 98980 3585 98982
rect 7956 99034 8012 99036
rect 8036 99034 8092 99036
rect 8116 99034 8172 99036
rect 8196 99034 8252 99036
rect 7956 98982 7982 99034
rect 7982 98982 8012 99034
rect 8036 98982 8046 99034
rect 8046 98982 8092 99034
rect 8116 98982 8162 99034
rect 8162 98982 8172 99034
rect 8196 98982 8226 99034
rect 8226 98982 8252 99034
rect 7956 98980 8012 98982
rect 8036 98980 8092 98982
rect 8116 98980 8172 98982
rect 8196 98980 8252 98982
rect 11150 98640 11206 98696
rect 5622 98490 5678 98492
rect 5702 98490 5758 98492
rect 5782 98490 5838 98492
rect 5862 98490 5918 98492
rect 5622 98438 5648 98490
rect 5648 98438 5678 98490
rect 5702 98438 5712 98490
rect 5712 98438 5758 98490
rect 5782 98438 5828 98490
rect 5828 98438 5838 98490
rect 5862 98438 5892 98490
rect 5892 98438 5918 98490
rect 5622 98436 5678 98438
rect 5702 98436 5758 98438
rect 5782 98436 5838 98438
rect 5862 98436 5918 98438
rect 10289 98490 10345 98492
rect 10369 98490 10425 98492
rect 10449 98490 10505 98492
rect 10529 98490 10585 98492
rect 10289 98438 10315 98490
rect 10315 98438 10345 98490
rect 10369 98438 10379 98490
rect 10379 98438 10425 98490
rect 10449 98438 10495 98490
rect 10495 98438 10505 98490
rect 10529 98438 10559 98490
rect 10559 98438 10585 98490
rect 10289 98436 10345 98438
rect 10369 98436 10425 98438
rect 10449 98436 10505 98438
rect 10529 98436 10585 98438
rect 3289 97946 3345 97948
rect 3369 97946 3425 97948
rect 3449 97946 3505 97948
rect 3529 97946 3585 97948
rect 3289 97894 3315 97946
rect 3315 97894 3345 97946
rect 3369 97894 3379 97946
rect 3379 97894 3425 97946
rect 3449 97894 3495 97946
rect 3495 97894 3505 97946
rect 3529 97894 3559 97946
rect 3559 97894 3585 97946
rect 3289 97892 3345 97894
rect 3369 97892 3425 97894
rect 3449 97892 3505 97894
rect 3529 97892 3585 97894
rect 7956 97946 8012 97948
rect 8036 97946 8092 97948
rect 8116 97946 8172 97948
rect 8196 97946 8252 97948
rect 7956 97894 7982 97946
rect 7982 97894 8012 97946
rect 8036 97894 8046 97946
rect 8046 97894 8092 97946
rect 8116 97894 8162 97946
rect 8162 97894 8172 97946
rect 8196 97894 8226 97946
rect 8226 97894 8252 97946
rect 7956 97892 8012 97894
rect 8036 97892 8092 97894
rect 8116 97892 8172 97894
rect 8196 97892 8252 97894
rect 5622 97402 5678 97404
rect 5702 97402 5758 97404
rect 5782 97402 5838 97404
rect 5862 97402 5918 97404
rect 5622 97350 5648 97402
rect 5648 97350 5678 97402
rect 5702 97350 5712 97402
rect 5712 97350 5758 97402
rect 5782 97350 5828 97402
rect 5828 97350 5838 97402
rect 5862 97350 5892 97402
rect 5892 97350 5918 97402
rect 5622 97348 5678 97350
rect 5702 97348 5758 97350
rect 5782 97348 5838 97350
rect 5862 97348 5918 97350
rect 10289 97402 10345 97404
rect 10369 97402 10425 97404
rect 10449 97402 10505 97404
rect 10529 97402 10585 97404
rect 10289 97350 10315 97402
rect 10315 97350 10345 97402
rect 10369 97350 10379 97402
rect 10379 97350 10425 97402
rect 10449 97350 10495 97402
rect 10495 97350 10505 97402
rect 10529 97350 10559 97402
rect 10559 97350 10585 97402
rect 10289 97348 10345 97350
rect 10369 97348 10425 97350
rect 10449 97348 10505 97350
rect 10529 97348 10585 97350
rect 110 97144 166 97200
rect 3289 96858 3345 96860
rect 3369 96858 3425 96860
rect 3449 96858 3505 96860
rect 3529 96858 3585 96860
rect 3289 96806 3315 96858
rect 3315 96806 3345 96858
rect 3369 96806 3379 96858
rect 3379 96806 3425 96858
rect 3449 96806 3495 96858
rect 3495 96806 3505 96858
rect 3529 96806 3559 96858
rect 3559 96806 3585 96858
rect 3289 96804 3345 96806
rect 3369 96804 3425 96806
rect 3449 96804 3505 96806
rect 3529 96804 3585 96806
rect 7956 96858 8012 96860
rect 8036 96858 8092 96860
rect 8116 96858 8172 96860
rect 8196 96858 8252 96860
rect 7956 96806 7982 96858
rect 7982 96806 8012 96858
rect 8036 96806 8046 96858
rect 8046 96806 8092 96858
rect 8116 96806 8162 96858
rect 8162 96806 8172 96858
rect 8196 96806 8226 96858
rect 8226 96806 8252 96858
rect 7956 96804 8012 96806
rect 8036 96804 8092 96806
rect 8116 96804 8172 96806
rect 8196 96804 8252 96806
rect 5622 96314 5678 96316
rect 5702 96314 5758 96316
rect 5782 96314 5838 96316
rect 5862 96314 5918 96316
rect 5622 96262 5648 96314
rect 5648 96262 5678 96314
rect 5702 96262 5712 96314
rect 5712 96262 5758 96314
rect 5782 96262 5828 96314
rect 5828 96262 5838 96314
rect 5862 96262 5892 96314
rect 5892 96262 5918 96314
rect 5622 96260 5678 96262
rect 5702 96260 5758 96262
rect 5782 96260 5838 96262
rect 5862 96260 5918 96262
rect 10289 96314 10345 96316
rect 10369 96314 10425 96316
rect 10449 96314 10505 96316
rect 10529 96314 10585 96316
rect 10289 96262 10315 96314
rect 10315 96262 10345 96314
rect 10369 96262 10379 96314
rect 10379 96262 10425 96314
rect 10449 96262 10495 96314
rect 10495 96262 10505 96314
rect 10529 96262 10559 96314
rect 10559 96262 10585 96314
rect 10289 96260 10345 96262
rect 10369 96260 10425 96262
rect 10449 96260 10505 96262
rect 10529 96260 10585 96262
rect 3289 95770 3345 95772
rect 3369 95770 3425 95772
rect 3449 95770 3505 95772
rect 3529 95770 3585 95772
rect 3289 95718 3315 95770
rect 3315 95718 3345 95770
rect 3369 95718 3379 95770
rect 3379 95718 3425 95770
rect 3449 95718 3495 95770
rect 3495 95718 3505 95770
rect 3529 95718 3559 95770
rect 3559 95718 3585 95770
rect 3289 95716 3345 95718
rect 3369 95716 3425 95718
rect 3449 95716 3505 95718
rect 3529 95716 3585 95718
rect 7956 95770 8012 95772
rect 8036 95770 8092 95772
rect 8116 95770 8172 95772
rect 8196 95770 8252 95772
rect 7956 95718 7982 95770
rect 7982 95718 8012 95770
rect 8036 95718 8046 95770
rect 8046 95718 8092 95770
rect 8116 95718 8162 95770
rect 8162 95718 8172 95770
rect 8196 95718 8226 95770
rect 8226 95718 8252 95770
rect 7956 95716 8012 95718
rect 8036 95716 8092 95718
rect 8116 95716 8172 95718
rect 8196 95716 8252 95718
rect 5622 95226 5678 95228
rect 5702 95226 5758 95228
rect 5782 95226 5838 95228
rect 5862 95226 5918 95228
rect 5622 95174 5648 95226
rect 5648 95174 5678 95226
rect 5702 95174 5712 95226
rect 5712 95174 5758 95226
rect 5782 95174 5828 95226
rect 5828 95174 5838 95226
rect 5862 95174 5892 95226
rect 5892 95174 5918 95226
rect 5622 95172 5678 95174
rect 5702 95172 5758 95174
rect 5782 95172 5838 95174
rect 5862 95172 5918 95174
rect 10289 95226 10345 95228
rect 10369 95226 10425 95228
rect 10449 95226 10505 95228
rect 10529 95226 10585 95228
rect 10289 95174 10315 95226
rect 10315 95174 10345 95226
rect 10369 95174 10379 95226
rect 10379 95174 10425 95226
rect 10449 95174 10495 95226
rect 10495 95174 10505 95226
rect 10529 95174 10559 95226
rect 10559 95174 10585 95226
rect 10289 95172 10345 95174
rect 10369 95172 10425 95174
rect 10449 95172 10505 95174
rect 10529 95172 10585 95174
rect 3289 94682 3345 94684
rect 3369 94682 3425 94684
rect 3449 94682 3505 94684
rect 3529 94682 3585 94684
rect 3289 94630 3315 94682
rect 3315 94630 3345 94682
rect 3369 94630 3379 94682
rect 3379 94630 3425 94682
rect 3449 94630 3495 94682
rect 3495 94630 3505 94682
rect 3529 94630 3559 94682
rect 3559 94630 3585 94682
rect 3289 94628 3345 94630
rect 3369 94628 3425 94630
rect 3449 94628 3505 94630
rect 3529 94628 3585 94630
rect 7956 94682 8012 94684
rect 8036 94682 8092 94684
rect 8116 94682 8172 94684
rect 8196 94682 8252 94684
rect 7956 94630 7982 94682
rect 7982 94630 8012 94682
rect 8036 94630 8046 94682
rect 8046 94630 8092 94682
rect 8116 94630 8162 94682
rect 8162 94630 8172 94682
rect 8196 94630 8226 94682
rect 8226 94630 8252 94682
rect 7956 94628 8012 94630
rect 8036 94628 8092 94630
rect 8116 94628 8172 94630
rect 8196 94628 8252 94630
rect 11242 97144 11298 97200
rect 5622 94138 5678 94140
rect 5702 94138 5758 94140
rect 5782 94138 5838 94140
rect 5862 94138 5918 94140
rect 5622 94086 5648 94138
rect 5648 94086 5678 94138
rect 5702 94086 5712 94138
rect 5712 94086 5758 94138
rect 5782 94086 5828 94138
rect 5828 94086 5838 94138
rect 5862 94086 5892 94138
rect 5892 94086 5918 94138
rect 5622 94084 5678 94086
rect 5702 94084 5758 94086
rect 5782 94084 5838 94086
rect 5862 94084 5918 94086
rect 10289 94138 10345 94140
rect 10369 94138 10425 94140
rect 10449 94138 10505 94140
rect 10529 94138 10585 94140
rect 10289 94086 10315 94138
rect 10315 94086 10345 94138
rect 10369 94086 10379 94138
rect 10379 94086 10425 94138
rect 10449 94086 10495 94138
rect 10495 94086 10505 94138
rect 10529 94086 10559 94138
rect 10559 94086 10585 94138
rect 10289 94084 10345 94086
rect 10369 94084 10425 94086
rect 10449 94084 10505 94086
rect 10529 94084 10585 94086
rect 3289 93594 3345 93596
rect 3369 93594 3425 93596
rect 3449 93594 3505 93596
rect 3529 93594 3585 93596
rect 3289 93542 3315 93594
rect 3315 93542 3345 93594
rect 3369 93542 3379 93594
rect 3379 93542 3425 93594
rect 3449 93542 3495 93594
rect 3495 93542 3505 93594
rect 3529 93542 3559 93594
rect 3559 93542 3585 93594
rect 3289 93540 3345 93542
rect 3369 93540 3425 93542
rect 3449 93540 3505 93542
rect 3529 93540 3585 93542
rect 7956 93594 8012 93596
rect 8036 93594 8092 93596
rect 8116 93594 8172 93596
rect 8196 93594 8252 93596
rect 7956 93542 7982 93594
rect 7982 93542 8012 93594
rect 8036 93542 8046 93594
rect 8046 93542 8092 93594
rect 8116 93542 8162 93594
rect 8162 93542 8172 93594
rect 8196 93542 8226 93594
rect 8226 93542 8252 93594
rect 7956 93540 8012 93542
rect 8036 93540 8092 93542
rect 8116 93540 8172 93542
rect 8196 93540 8252 93542
rect 5622 93050 5678 93052
rect 5702 93050 5758 93052
rect 5782 93050 5838 93052
rect 5862 93050 5918 93052
rect 5622 92998 5648 93050
rect 5648 92998 5678 93050
rect 5702 92998 5712 93050
rect 5712 92998 5758 93050
rect 5782 92998 5828 93050
rect 5828 92998 5838 93050
rect 5862 92998 5892 93050
rect 5892 92998 5918 93050
rect 5622 92996 5678 92998
rect 5702 92996 5758 92998
rect 5782 92996 5838 92998
rect 5862 92996 5918 92998
rect 10289 93050 10345 93052
rect 10369 93050 10425 93052
rect 10449 93050 10505 93052
rect 10529 93050 10585 93052
rect 10289 92998 10315 93050
rect 10315 92998 10345 93050
rect 10369 92998 10379 93050
rect 10379 92998 10425 93050
rect 10449 92998 10495 93050
rect 10495 92998 10505 93050
rect 10529 92998 10559 93050
rect 10559 92998 10585 93050
rect 10289 92996 10345 92998
rect 10369 92996 10425 92998
rect 10449 92996 10505 92998
rect 10529 92996 10585 92998
rect 3289 92506 3345 92508
rect 3369 92506 3425 92508
rect 3449 92506 3505 92508
rect 3529 92506 3585 92508
rect 3289 92454 3315 92506
rect 3315 92454 3345 92506
rect 3369 92454 3379 92506
rect 3379 92454 3425 92506
rect 3449 92454 3495 92506
rect 3495 92454 3505 92506
rect 3529 92454 3559 92506
rect 3559 92454 3585 92506
rect 3289 92452 3345 92454
rect 3369 92452 3425 92454
rect 3449 92452 3505 92454
rect 3529 92452 3585 92454
rect 7956 92506 8012 92508
rect 8036 92506 8092 92508
rect 8116 92506 8172 92508
rect 8196 92506 8252 92508
rect 7956 92454 7982 92506
rect 7982 92454 8012 92506
rect 8036 92454 8046 92506
rect 8046 92454 8092 92506
rect 8116 92454 8162 92506
rect 8162 92454 8172 92506
rect 8196 92454 8226 92506
rect 8226 92454 8252 92506
rect 7956 92452 8012 92454
rect 8036 92452 8092 92454
rect 8116 92452 8172 92454
rect 8196 92452 8252 92454
rect 5622 91962 5678 91964
rect 5702 91962 5758 91964
rect 5782 91962 5838 91964
rect 5862 91962 5918 91964
rect 5622 91910 5648 91962
rect 5648 91910 5678 91962
rect 5702 91910 5712 91962
rect 5712 91910 5758 91962
rect 5782 91910 5828 91962
rect 5828 91910 5838 91962
rect 5862 91910 5892 91962
rect 5892 91910 5918 91962
rect 5622 91908 5678 91910
rect 5702 91908 5758 91910
rect 5782 91908 5838 91910
rect 5862 91908 5918 91910
rect 10289 91962 10345 91964
rect 10369 91962 10425 91964
rect 10449 91962 10505 91964
rect 10529 91962 10585 91964
rect 10289 91910 10315 91962
rect 10315 91910 10345 91962
rect 10369 91910 10379 91962
rect 10379 91910 10425 91962
rect 10449 91910 10495 91962
rect 10495 91910 10505 91962
rect 10529 91910 10559 91962
rect 10559 91910 10585 91962
rect 10289 91908 10345 91910
rect 10369 91908 10425 91910
rect 10449 91908 10505 91910
rect 10529 91908 10585 91910
rect 10690 91840 10746 91896
rect 3289 91418 3345 91420
rect 3369 91418 3425 91420
rect 3449 91418 3505 91420
rect 3529 91418 3585 91420
rect 3289 91366 3315 91418
rect 3315 91366 3345 91418
rect 3369 91366 3379 91418
rect 3379 91366 3425 91418
rect 3449 91366 3495 91418
rect 3495 91366 3505 91418
rect 3529 91366 3559 91418
rect 3559 91366 3585 91418
rect 3289 91364 3345 91366
rect 3369 91364 3425 91366
rect 3449 91364 3505 91366
rect 3529 91364 3585 91366
rect 7956 91418 8012 91420
rect 8036 91418 8092 91420
rect 8116 91418 8172 91420
rect 8196 91418 8252 91420
rect 7956 91366 7982 91418
rect 7982 91366 8012 91418
rect 8036 91366 8046 91418
rect 8046 91366 8092 91418
rect 8116 91366 8162 91418
rect 8162 91366 8172 91418
rect 8196 91366 8226 91418
rect 8226 91366 8252 91418
rect 7956 91364 8012 91366
rect 8036 91364 8092 91366
rect 8116 91364 8172 91366
rect 8196 91364 8252 91366
rect 5622 90874 5678 90876
rect 5702 90874 5758 90876
rect 5782 90874 5838 90876
rect 5862 90874 5918 90876
rect 5622 90822 5648 90874
rect 5648 90822 5678 90874
rect 5702 90822 5712 90874
rect 5712 90822 5758 90874
rect 5782 90822 5828 90874
rect 5828 90822 5838 90874
rect 5862 90822 5892 90874
rect 5892 90822 5918 90874
rect 5622 90820 5678 90822
rect 5702 90820 5758 90822
rect 5782 90820 5838 90822
rect 5862 90820 5918 90822
rect 10289 90874 10345 90876
rect 10369 90874 10425 90876
rect 10449 90874 10505 90876
rect 10529 90874 10585 90876
rect 10289 90822 10315 90874
rect 10315 90822 10345 90874
rect 10369 90822 10379 90874
rect 10379 90822 10425 90874
rect 10449 90822 10495 90874
rect 10495 90822 10505 90874
rect 10529 90822 10559 90874
rect 10559 90822 10585 90874
rect 10289 90820 10345 90822
rect 10369 90820 10425 90822
rect 10449 90820 10505 90822
rect 10529 90820 10585 90822
rect 3289 90330 3345 90332
rect 3369 90330 3425 90332
rect 3449 90330 3505 90332
rect 3529 90330 3585 90332
rect 3289 90278 3315 90330
rect 3315 90278 3345 90330
rect 3369 90278 3379 90330
rect 3379 90278 3425 90330
rect 3449 90278 3495 90330
rect 3495 90278 3505 90330
rect 3529 90278 3559 90330
rect 3559 90278 3585 90330
rect 3289 90276 3345 90278
rect 3369 90276 3425 90278
rect 3449 90276 3505 90278
rect 3529 90276 3585 90278
rect 7956 90330 8012 90332
rect 8036 90330 8092 90332
rect 8116 90330 8172 90332
rect 8196 90330 8252 90332
rect 7956 90278 7982 90330
rect 7982 90278 8012 90330
rect 8036 90278 8046 90330
rect 8046 90278 8092 90330
rect 8116 90278 8162 90330
rect 8162 90278 8172 90330
rect 8196 90278 8226 90330
rect 8226 90278 8252 90330
rect 7956 90276 8012 90278
rect 8036 90276 8092 90278
rect 8116 90276 8172 90278
rect 8196 90276 8252 90278
rect 5622 89786 5678 89788
rect 5702 89786 5758 89788
rect 5782 89786 5838 89788
rect 5862 89786 5918 89788
rect 5622 89734 5648 89786
rect 5648 89734 5678 89786
rect 5702 89734 5712 89786
rect 5712 89734 5758 89786
rect 5782 89734 5828 89786
rect 5828 89734 5838 89786
rect 5862 89734 5892 89786
rect 5892 89734 5918 89786
rect 5622 89732 5678 89734
rect 5702 89732 5758 89734
rect 5782 89732 5838 89734
rect 5862 89732 5918 89734
rect 10289 89786 10345 89788
rect 10369 89786 10425 89788
rect 10449 89786 10505 89788
rect 10529 89786 10585 89788
rect 10289 89734 10315 89786
rect 10315 89734 10345 89786
rect 10369 89734 10379 89786
rect 10379 89734 10425 89786
rect 10449 89734 10495 89786
rect 10495 89734 10505 89786
rect 10529 89734 10559 89786
rect 10559 89734 10585 89786
rect 10289 89732 10345 89734
rect 10369 89732 10425 89734
rect 10449 89732 10505 89734
rect 10529 89732 10585 89734
rect 3289 89242 3345 89244
rect 3369 89242 3425 89244
rect 3449 89242 3505 89244
rect 3529 89242 3585 89244
rect 3289 89190 3315 89242
rect 3315 89190 3345 89242
rect 3369 89190 3379 89242
rect 3379 89190 3425 89242
rect 3449 89190 3495 89242
rect 3495 89190 3505 89242
rect 3529 89190 3559 89242
rect 3559 89190 3585 89242
rect 3289 89188 3345 89190
rect 3369 89188 3425 89190
rect 3449 89188 3505 89190
rect 3529 89188 3585 89190
rect 7956 89242 8012 89244
rect 8036 89242 8092 89244
rect 8116 89242 8172 89244
rect 8196 89242 8252 89244
rect 7956 89190 7982 89242
rect 7982 89190 8012 89242
rect 8036 89190 8046 89242
rect 8046 89190 8092 89242
rect 8116 89190 8162 89242
rect 8162 89190 8172 89242
rect 8196 89190 8226 89242
rect 8226 89190 8252 89242
rect 7956 89188 8012 89190
rect 8036 89188 8092 89190
rect 8116 89188 8172 89190
rect 8196 89188 8252 89190
rect 5622 88698 5678 88700
rect 5702 88698 5758 88700
rect 5782 88698 5838 88700
rect 5862 88698 5918 88700
rect 5622 88646 5648 88698
rect 5648 88646 5678 88698
rect 5702 88646 5712 88698
rect 5712 88646 5758 88698
rect 5782 88646 5828 88698
rect 5828 88646 5838 88698
rect 5862 88646 5892 88698
rect 5892 88646 5918 88698
rect 5622 88644 5678 88646
rect 5702 88644 5758 88646
rect 5782 88644 5838 88646
rect 5862 88644 5918 88646
rect 10289 88698 10345 88700
rect 10369 88698 10425 88700
rect 10449 88698 10505 88700
rect 10529 88698 10585 88700
rect 10289 88646 10315 88698
rect 10315 88646 10345 88698
rect 10369 88646 10379 88698
rect 10379 88646 10425 88698
rect 10449 88646 10495 88698
rect 10495 88646 10505 88698
rect 10529 88646 10559 88698
rect 10559 88646 10585 88698
rect 10289 88644 10345 88646
rect 10369 88644 10425 88646
rect 10449 88644 10505 88646
rect 10529 88644 10585 88646
rect 110 88440 166 88496
rect 3289 88154 3345 88156
rect 3369 88154 3425 88156
rect 3449 88154 3505 88156
rect 3529 88154 3585 88156
rect 3289 88102 3315 88154
rect 3315 88102 3345 88154
rect 3369 88102 3379 88154
rect 3379 88102 3425 88154
rect 3449 88102 3495 88154
rect 3495 88102 3505 88154
rect 3529 88102 3559 88154
rect 3559 88102 3585 88154
rect 3289 88100 3345 88102
rect 3369 88100 3425 88102
rect 3449 88100 3505 88102
rect 3529 88100 3585 88102
rect 7956 88154 8012 88156
rect 8036 88154 8092 88156
rect 8116 88154 8172 88156
rect 8196 88154 8252 88156
rect 7956 88102 7982 88154
rect 7982 88102 8012 88154
rect 8036 88102 8046 88154
rect 8046 88102 8092 88154
rect 8116 88102 8162 88154
rect 8162 88102 8172 88154
rect 8196 88102 8226 88154
rect 8226 88102 8252 88154
rect 7956 88100 8012 88102
rect 8036 88100 8092 88102
rect 8116 88100 8172 88102
rect 8196 88100 8252 88102
rect 5622 87610 5678 87612
rect 5702 87610 5758 87612
rect 5782 87610 5838 87612
rect 5862 87610 5918 87612
rect 5622 87558 5648 87610
rect 5648 87558 5678 87610
rect 5702 87558 5712 87610
rect 5712 87558 5758 87610
rect 5782 87558 5828 87610
rect 5828 87558 5838 87610
rect 5862 87558 5892 87610
rect 5892 87558 5918 87610
rect 5622 87556 5678 87558
rect 5702 87556 5758 87558
rect 5782 87556 5838 87558
rect 5862 87556 5918 87558
rect 10289 87610 10345 87612
rect 10369 87610 10425 87612
rect 10449 87610 10505 87612
rect 10529 87610 10585 87612
rect 10289 87558 10315 87610
rect 10315 87558 10345 87610
rect 10369 87558 10379 87610
rect 10379 87558 10425 87610
rect 10449 87558 10495 87610
rect 10495 87558 10505 87610
rect 10529 87558 10559 87610
rect 10559 87558 10585 87610
rect 10289 87556 10345 87558
rect 10369 87556 10425 87558
rect 10449 87556 10505 87558
rect 10529 87556 10585 87558
rect 3289 87066 3345 87068
rect 3369 87066 3425 87068
rect 3449 87066 3505 87068
rect 3529 87066 3585 87068
rect 3289 87014 3315 87066
rect 3315 87014 3345 87066
rect 3369 87014 3379 87066
rect 3379 87014 3425 87066
rect 3449 87014 3495 87066
rect 3495 87014 3505 87066
rect 3529 87014 3559 87066
rect 3559 87014 3585 87066
rect 3289 87012 3345 87014
rect 3369 87012 3425 87014
rect 3449 87012 3505 87014
rect 3529 87012 3585 87014
rect 7956 87066 8012 87068
rect 8036 87066 8092 87068
rect 8116 87066 8172 87068
rect 8196 87066 8252 87068
rect 7956 87014 7982 87066
rect 7982 87014 8012 87066
rect 8036 87014 8046 87066
rect 8046 87014 8092 87066
rect 8116 87014 8162 87066
rect 8162 87014 8172 87066
rect 8196 87014 8226 87066
rect 8226 87014 8252 87066
rect 7956 87012 8012 87014
rect 8036 87012 8092 87014
rect 8116 87012 8172 87014
rect 8196 87012 8252 87014
rect 5622 86522 5678 86524
rect 5702 86522 5758 86524
rect 5782 86522 5838 86524
rect 5862 86522 5918 86524
rect 5622 86470 5648 86522
rect 5648 86470 5678 86522
rect 5702 86470 5712 86522
rect 5712 86470 5758 86522
rect 5782 86470 5828 86522
rect 5828 86470 5838 86522
rect 5862 86470 5892 86522
rect 5892 86470 5918 86522
rect 5622 86468 5678 86470
rect 5702 86468 5758 86470
rect 5782 86468 5838 86470
rect 5862 86468 5918 86470
rect 10289 86522 10345 86524
rect 10369 86522 10425 86524
rect 10449 86522 10505 86524
rect 10529 86522 10585 86524
rect 10289 86470 10315 86522
rect 10315 86470 10345 86522
rect 10369 86470 10379 86522
rect 10379 86470 10425 86522
rect 10449 86470 10495 86522
rect 10495 86470 10505 86522
rect 10529 86470 10559 86522
rect 10559 86470 10585 86522
rect 10289 86468 10345 86470
rect 10369 86468 10425 86470
rect 10449 86468 10505 86470
rect 10529 86468 10585 86470
rect 3289 85978 3345 85980
rect 3369 85978 3425 85980
rect 3449 85978 3505 85980
rect 3529 85978 3585 85980
rect 3289 85926 3315 85978
rect 3315 85926 3345 85978
rect 3369 85926 3379 85978
rect 3379 85926 3425 85978
rect 3449 85926 3495 85978
rect 3495 85926 3505 85978
rect 3529 85926 3559 85978
rect 3559 85926 3585 85978
rect 3289 85924 3345 85926
rect 3369 85924 3425 85926
rect 3449 85924 3505 85926
rect 3529 85924 3585 85926
rect 7956 85978 8012 85980
rect 8036 85978 8092 85980
rect 8116 85978 8172 85980
rect 8196 85978 8252 85980
rect 7956 85926 7982 85978
rect 7982 85926 8012 85978
rect 8036 85926 8046 85978
rect 8046 85926 8092 85978
rect 8116 85926 8162 85978
rect 8162 85926 8172 85978
rect 8196 85926 8226 85978
rect 8226 85926 8252 85978
rect 7956 85924 8012 85926
rect 8036 85924 8092 85926
rect 8116 85924 8172 85926
rect 8196 85924 8252 85926
rect 5622 85434 5678 85436
rect 5702 85434 5758 85436
rect 5782 85434 5838 85436
rect 5862 85434 5918 85436
rect 5622 85382 5648 85434
rect 5648 85382 5678 85434
rect 5702 85382 5712 85434
rect 5712 85382 5758 85434
rect 5782 85382 5828 85434
rect 5828 85382 5838 85434
rect 5862 85382 5892 85434
rect 5892 85382 5918 85434
rect 5622 85380 5678 85382
rect 5702 85380 5758 85382
rect 5782 85380 5838 85382
rect 5862 85380 5918 85382
rect 10289 85434 10345 85436
rect 10369 85434 10425 85436
rect 10449 85434 10505 85436
rect 10529 85434 10585 85436
rect 10289 85382 10315 85434
rect 10315 85382 10345 85434
rect 10369 85382 10379 85434
rect 10379 85382 10425 85434
rect 10449 85382 10495 85434
rect 10495 85382 10505 85434
rect 10529 85382 10559 85434
rect 10559 85382 10585 85434
rect 10289 85380 10345 85382
rect 10369 85380 10425 85382
rect 10449 85380 10505 85382
rect 10529 85380 10585 85382
rect 110 85176 166 85232
rect 3289 84890 3345 84892
rect 3369 84890 3425 84892
rect 3449 84890 3505 84892
rect 3529 84890 3585 84892
rect 3289 84838 3315 84890
rect 3315 84838 3345 84890
rect 3369 84838 3379 84890
rect 3379 84838 3425 84890
rect 3449 84838 3495 84890
rect 3495 84838 3505 84890
rect 3529 84838 3559 84890
rect 3559 84838 3585 84890
rect 3289 84836 3345 84838
rect 3369 84836 3425 84838
rect 3449 84836 3505 84838
rect 3529 84836 3585 84838
rect 7956 84890 8012 84892
rect 8036 84890 8092 84892
rect 8116 84890 8172 84892
rect 8196 84890 8252 84892
rect 7956 84838 7982 84890
rect 7982 84838 8012 84890
rect 8036 84838 8046 84890
rect 8046 84838 8092 84890
rect 8116 84838 8162 84890
rect 8162 84838 8172 84890
rect 8196 84838 8226 84890
rect 8226 84838 8252 84890
rect 7956 84836 8012 84838
rect 8036 84836 8092 84838
rect 8116 84836 8172 84838
rect 8196 84836 8252 84838
rect 5622 84346 5678 84348
rect 5702 84346 5758 84348
rect 5782 84346 5838 84348
rect 5862 84346 5918 84348
rect 5622 84294 5648 84346
rect 5648 84294 5678 84346
rect 5702 84294 5712 84346
rect 5712 84294 5758 84346
rect 5782 84294 5828 84346
rect 5828 84294 5838 84346
rect 5862 84294 5892 84346
rect 5892 84294 5918 84346
rect 5622 84292 5678 84294
rect 5702 84292 5758 84294
rect 5782 84292 5838 84294
rect 5862 84292 5918 84294
rect 10289 84346 10345 84348
rect 10369 84346 10425 84348
rect 10449 84346 10505 84348
rect 10529 84346 10585 84348
rect 10289 84294 10315 84346
rect 10315 84294 10345 84346
rect 10369 84294 10379 84346
rect 10379 84294 10425 84346
rect 10449 84294 10495 84346
rect 10495 84294 10505 84346
rect 10529 84294 10559 84346
rect 10559 84294 10585 84346
rect 10289 84292 10345 84294
rect 10369 84292 10425 84294
rect 10449 84292 10505 84294
rect 10529 84292 10585 84294
rect 3289 83802 3345 83804
rect 3369 83802 3425 83804
rect 3449 83802 3505 83804
rect 3529 83802 3585 83804
rect 3289 83750 3315 83802
rect 3315 83750 3345 83802
rect 3369 83750 3379 83802
rect 3379 83750 3425 83802
rect 3449 83750 3495 83802
rect 3495 83750 3505 83802
rect 3529 83750 3559 83802
rect 3559 83750 3585 83802
rect 3289 83748 3345 83750
rect 3369 83748 3425 83750
rect 3449 83748 3505 83750
rect 3529 83748 3585 83750
rect 7956 83802 8012 83804
rect 8036 83802 8092 83804
rect 8116 83802 8172 83804
rect 8196 83802 8252 83804
rect 7956 83750 7982 83802
rect 7982 83750 8012 83802
rect 8036 83750 8046 83802
rect 8046 83750 8092 83802
rect 8116 83750 8162 83802
rect 8162 83750 8172 83802
rect 8196 83750 8226 83802
rect 8226 83750 8252 83802
rect 7956 83748 8012 83750
rect 8036 83748 8092 83750
rect 8116 83748 8172 83750
rect 8196 83748 8252 83750
rect 5622 83258 5678 83260
rect 5702 83258 5758 83260
rect 5782 83258 5838 83260
rect 5862 83258 5918 83260
rect 5622 83206 5648 83258
rect 5648 83206 5678 83258
rect 5702 83206 5712 83258
rect 5712 83206 5758 83258
rect 5782 83206 5828 83258
rect 5828 83206 5838 83258
rect 5862 83206 5892 83258
rect 5892 83206 5918 83258
rect 5622 83204 5678 83206
rect 5702 83204 5758 83206
rect 5782 83204 5838 83206
rect 5862 83204 5918 83206
rect 10289 83258 10345 83260
rect 10369 83258 10425 83260
rect 10449 83258 10505 83260
rect 10529 83258 10585 83260
rect 10289 83206 10315 83258
rect 10315 83206 10345 83258
rect 10369 83206 10379 83258
rect 10379 83206 10425 83258
rect 10449 83206 10495 83258
rect 10495 83206 10505 83258
rect 10529 83206 10559 83258
rect 10559 83206 10585 83258
rect 10289 83204 10345 83206
rect 10369 83204 10425 83206
rect 10449 83204 10505 83206
rect 10529 83204 10585 83206
rect 3289 82714 3345 82716
rect 3369 82714 3425 82716
rect 3449 82714 3505 82716
rect 3529 82714 3585 82716
rect 3289 82662 3315 82714
rect 3315 82662 3345 82714
rect 3369 82662 3379 82714
rect 3379 82662 3425 82714
rect 3449 82662 3495 82714
rect 3495 82662 3505 82714
rect 3529 82662 3559 82714
rect 3559 82662 3585 82714
rect 3289 82660 3345 82662
rect 3369 82660 3425 82662
rect 3449 82660 3505 82662
rect 3529 82660 3585 82662
rect 7956 82714 8012 82716
rect 8036 82714 8092 82716
rect 8116 82714 8172 82716
rect 8196 82714 8252 82716
rect 7956 82662 7982 82714
rect 7982 82662 8012 82714
rect 8036 82662 8046 82714
rect 8046 82662 8092 82714
rect 8116 82662 8162 82714
rect 8162 82662 8172 82714
rect 8196 82662 8226 82714
rect 8226 82662 8252 82714
rect 7956 82660 8012 82662
rect 8036 82660 8092 82662
rect 8116 82660 8172 82662
rect 8196 82660 8252 82662
rect 5622 82170 5678 82172
rect 5702 82170 5758 82172
rect 5782 82170 5838 82172
rect 5862 82170 5918 82172
rect 5622 82118 5648 82170
rect 5648 82118 5678 82170
rect 5702 82118 5712 82170
rect 5712 82118 5758 82170
rect 5782 82118 5828 82170
rect 5828 82118 5838 82170
rect 5862 82118 5892 82170
rect 5892 82118 5918 82170
rect 5622 82116 5678 82118
rect 5702 82116 5758 82118
rect 5782 82116 5838 82118
rect 5862 82116 5918 82118
rect 10289 82170 10345 82172
rect 10369 82170 10425 82172
rect 10449 82170 10505 82172
rect 10529 82170 10585 82172
rect 10289 82118 10315 82170
rect 10315 82118 10345 82170
rect 10369 82118 10379 82170
rect 10379 82118 10425 82170
rect 10449 82118 10495 82170
rect 10495 82118 10505 82170
rect 10529 82118 10559 82170
rect 10559 82118 10585 82170
rect 10289 82116 10345 82118
rect 10369 82116 10425 82118
rect 10449 82116 10505 82118
rect 10529 82116 10585 82118
rect 3289 81626 3345 81628
rect 3369 81626 3425 81628
rect 3449 81626 3505 81628
rect 3529 81626 3585 81628
rect 3289 81574 3315 81626
rect 3315 81574 3345 81626
rect 3369 81574 3379 81626
rect 3379 81574 3425 81626
rect 3449 81574 3495 81626
rect 3495 81574 3505 81626
rect 3529 81574 3559 81626
rect 3559 81574 3585 81626
rect 3289 81572 3345 81574
rect 3369 81572 3425 81574
rect 3449 81572 3505 81574
rect 3529 81572 3585 81574
rect 7956 81626 8012 81628
rect 8036 81626 8092 81628
rect 8116 81626 8172 81628
rect 8196 81626 8252 81628
rect 7956 81574 7982 81626
rect 7982 81574 8012 81626
rect 8036 81574 8046 81626
rect 8046 81574 8092 81626
rect 8116 81574 8162 81626
rect 8162 81574 8172 81626
rect 8196 81574 8226 81626
rect 8226 81574 8252 81626
rect 7956 81572 8012 81574
rect 8036 81572 8092 81574
rect 8116 81572 8172 81574
rect 8196 81572 8252 81574
rect 5622 81082 5678 81084
rect 5702 81082 5758 81084
rect 5782 81082 5838 81084
rect 5862 81082 5918 81084
rect 5622 81030 5648 81082
rect 5648 81030 5678 81082
rect 5702 81030 5712 81082
rect 5712 81030 5758 81082
rect 5782 81030 5828 81082
rect 5828 81030 5838 81082
rect 5862 81030 5892 81082
rect 5892 81030 5918 81082
rect 5622 81028 5678 81030
rect 5702 81028 5758 81030
rect 5782 81028 5838 81030
rect 5862 81028 5918 81030
rect 10289 81082 10345 81084
rect 10369 81082 10425 81084
rect 10449 81082 10505 81084
rect 10529 81082 10585 81084
rect 10289 81030 10315 81082
rect 10315 81030 10345 81082
rect 10369 81030 10379 81082
rect 10379 81030 10425 81082
rect 10449 81030 10495 81082
rect 10495 81030 10505 81082
rect 10529 81030 10559 81082
rect 10559 81030 10585 81082
rect 10289 81028 10345 81030
rect 10369 81028 10425 81030
rect 10449 81028 10505 81030
rect 10529 81028 10585 81030
rect 3289 80538 3345 80540
rect 3369 80538 3425 80540
rect 3449 80538 3505 80540
rect 3529 80538 3585 80540
rect 3289 80486 3315 80538
rect 3315 80486 3345 80538
rect 3369 80486 3379 80538
rect 3379 80486 3425 80538
rect 3449 80486 3495 80538
rect 3495 80486 3505 80538
rect 3529 80486 3559 80538
rect 3559 80486 3585 80538
rect 3289 80484 3345 80486
rect 3369 80484 3425 80486
rect 3449 80484 3505 80486
rect 3529 80484 3585 80486
rect 7956 80538 8012 80540
rect 8036 80538 8092 80540
rect 8116 80538 8172 80540
rect 8196 80538 8252 80540
rect 7956 80486 7982 80538
rect 7982 80486 8012 80538
rect 8036 80486 8046 80538
rect 8046 80486 8092 80538
rect 8116 80486 8162 80538
rect 8162 80486 8172 80538
rect 8196 80486 8226 80538
rect 8226 80486 8252 80538
rect 7956 80484 8012 80486
rect 8036 80484 8092 80486
rect 8116 80484 8172 80486
rect 8196 80484 8252 80486
rect 5622 79994 5678 79996
rect 5702 79994 5758 79996
rect 5782 79994 5838 79996
rect 5862 79994 5918 79996
rect 5622 79942 5648 79994
rect 5648 79942 5678 79994
rect 5702 79942 5712 79994
rect 5712 79942 5758 79994
rect 5782 79942 5828 79994
rect 5828 79942 5838 79994
rect 5862 79942 5892 79994
rect 5892 79942 5918 79994
rect 5622 79940 5678 79942
rect 5702 79940 5758 79942
rect 5782 79940 5838 79942
rect 5862 79940 5918 79942
rect 10289 79994 10345 79996
rect 10369 79994 10425 79996
rect 10449 79994 10505 79996
rect 10529 79994 10585 79996
rect 10289 79942 10315 79994
rect 10315 79942 10345 79994
rect 10369 79942 10379 79994
rect 10379 79942 10425 79994
rect 10449 79942 10495 79994
rect 10495 79942 10505 79994
rect 10529 79942 10559 79994
rect 10559 79942 10585 79994
rect 10289 79940 10345 79942
rect 10369 79940 10425 79942
rect 10449 79940 10505 79942
rect 10529 79940 10585 79942
rect 3289 79450 3345 79452
rect 3369 79450 3425 79452
rect 3449 79450 3505 79452
rect 3529 79450 3585 79452
rect 3289 79398 3315 79450
rect 3315 79398 3345 79450
rect 3369 79398 3379 79450
rect 3379 79398 3425 79450
rect 3449 79398 3495 79450
rect 3495 79398 3505 79450
rect 3529 79398 3559 79450
rect 3559 79398 3585 79450
rect 3289 79396 3345 79398
rect 3369 79396 3425 79398
rect 3449 79396 3505 79398
rect 3529 79396 3585 79398
rect 7956 79450 8012 79452
rect 8036 79450 8092 79452
rect 8116 79450 8172 79452
rect 8196 79450 8252 79452
rect 7956 79398 7982 79450
rect 7982 79398 8012 79450
rect 8036 79398 8046 79450
rect 8046 79398 8092 79450
rect 8116 79398 8162 79450
rect 8162 79398 8172 79450
rect 8196 79398 8226 79450
rect 8226 79398 8252 79450
rect 7956 79396 8012 79398
rect 8036 79396 8092 79398
rect 8116 79396 8172 79398
rect 8196 79396 8252 79398
rect 5622 78906 5678 78908
rect 5702 78906 5758 78908
rect 5782 78906 5838 78908
rect 5862 78906 5918 78908
rect 5622 78854 5648 78906
rect 5648 78854 5678 78906
rect 5702 78854 5712 78906
rect 5712 78854 5758 78906
rect 5782 78854 5828 78906
rect 5828 78854 5838 78906
rect 5862 78854 5892 78906
rect 5892 78854 5918 78906
rect 5622 78852 5678 78854
rect 5702 78852 5758 78854
rect 5782 78852 5838 78854
rect 5862 78852 5918 78854
rect 10289 78906 10345 78908
rect 10369 78906 10425 78908
rect 10449 78906 10505 78908
rect 10529 78906 10585 78908
rect 10289 78854 10315 78906
rect 10315 78854 10345 78906
rect 10369 78854 10379 78906
rect 10379 78854 10425 78906
rect 10449 78854 10495 78906
rect 10495 78854 10505 78906
rect 10529 78854 10559 78906
rect 10559 78854 10585 78906
rect 10289 78852 10345 78854
rect 10369 78852 10425 78854
rect 10449 78852 10505 78854
rect 10529 78852 10585 78854
rect 3289 78362 3345 78364
rect 3369 78362 3425 78364
rect 3449 78362 3505 78364
rect 3529 78362 3585 78364
rect 3289 78310 3315 78362
rect 3315 78310 3345 78362
rect 3369 78310 3379 78362
rect 3379 78310 3425 78362
rect 3449 78310 3495 78362
rect 3495 78310 3505 78362
rect 3529 78310 3559 78362
rect 3559 78310 3585 78362
rect 3289 78308 3345 78310
rect 3369 78308 3425 78310
rect 3449 78308 3505 78310
rect 3529 78308 3585 78310
rect 7956 78362 8012 78364
rect 8036 78362 8092 78364
rect 8116 78362 8172 78364
rect 8196 78362 8252 78364
rect 7956 78310 7982 78362
rect 7982 78310 8012 78362
rect 8036 78310 8046 78362
rect 8046 78310 8092 78362
rect 8116 78310 8162 78362
rect 8162 78310 8172 78362
rect 8196 78310 8226 78362
rect 8226 78310 8252 78362
rect 7956 78308 8012 78310
rect 8036 78308 8092 78310
rect 8116 78308 8172 78310
rect 8196 78308 8252 78310
rect 10966 78240 11022 78296
rect 5622 77818 5678 77820
rect 5702 77818 5758 77820
rect 5782 77818 5838 77820
rect 5862 77818 5918 77820
rect 5622 77766 5648 77818
rect 5648 77766 5678 77818
rect 5702 77766 5712 77818
rect 5712 77766 5758 77818
rect 5782 77766 5828 77818
rect 5828 77766 5838 77818
rect 5862 77766 5892 77818
rect 5892 77766 5918 77818
rect 5622 77764 5678 77766
rect 5702 77764 5758 77766
rect 5782 77764 5838 77766
rect 5862 77764 5918 77766
rect 10289 77818 10345 77820
rect 10369 77818 10425 77820
rect 10449 77818 10505 77820
rect 10529 77818 10585 77820
rect 10289 77766 10315 77818
rect 10315 77766 10345 77818
rect 10369 77766 10379 77818
rect 10379 77766 10425 77818
rect 10449 77766 10495 77818
rect 10495 77766 10505 77818
rect 10529 77766 10559 77818
rect 10559 77766 10585 77818
rect 10289 77764 10345 77766
rect 10369 77764 10425 77766
rect 10449 77764 10505 77766
rect 10529 77764 10585 77766
rect 3289 77274 3345 77276
rect 3369 77274 3425 77276
rect 3449 77274 3505 77276
rect 3529 77274 3585 77276
rect 3289 77222 3315 77274
rect 3315 77222 3345 77274
rect 3369 77222 3379 77274
rect 3379 77222 3425 77274
rect 3449 77222 3495 77274
rect 3495 77222 3505 77274
rect 3529 77222 3559 77274
rect 3559 77222 3585 77274
rect 3289 77220 3345 77222
rect 3369 77220 3425 77222
rect 3449 77220 3505 77222
rect 3529 77220 3585 77222
rect 7956 77274 8012 77276
rect 8036 77274 8092 77276
rect 8116 77274 8172 77276
rect 8196 77274 8252 77276
rect 7956 77222 7982 77274
rect 7982 77222 8012 77274
rect 8036 77222 8046 77274
rect 8046 77222 8092 77274
rect 8116 77222 8162 77274
rect 8162 77222 8172 77274
rect 8196 77222 8226 77274
rect 8226 77222 8252 77274
rect 7956 77220 8012 77222
rect 8036 77220 8092 77222
rect 8116 77220 8172 77222
rect 8196 77220 8252 77222
rect 5622 76730 5678 76732
rect 5702 76730 5758 76732
rect 5782 76730 5838 76732
rect 5862 76730 5918 76732
rect 5622 76678 5648 76730
rect 5648 76678 5678 76730
rect 5702 76678 5712 76730
rect 5712 76678 5758 76730
rect 5782 76678 5828 76730
rect 5828 76678 5838 76730
rect 5862 76678 5892 76730
rect 5892 76678 5918 76730
rect 5622 76676 5678 76678
rect 5702 76676 5758 76678
rect 5782 76676 5838 76678
rect 5862 76676 5918 76678
rect 10289 76730 10345 76732
rect 10369 76730 10425 76732
rect 10449 76730 10505 76732
rect 10529 76730 10585 76732
rect 10289 76678 10315 76730
rect 10315 76678 10345 76730
rect 10369 76678 10379 76730
rect 10379 76678 10425 76730
rect 10449 76678 10495 76730
rect 10495 76678 10505 76730
rect 10529 76678 10559 76730
rect 10559 76678 10585 76730
rect 10289 76676 10345 76678
rect 10369 76676 10425 76678
rect 10449 76676 10505 76678
rect 10529 76676 10585 76678
rect 3289 76186 3345 76188
rect 3369 76186 3425 76188
rect 3449 76186 3505 76188
rect 3529 76186 3585 76188
rect 3289 76134 3315 76186
rect 3315 76134 3345 76186
rect 3369 76134 3379 76186
rect 3379 76134 3425 76186
rect 3449 76134 3495 76186
rect 3495 76134 3505 76186
rect 3529 76134 3559 76186
rect 3559 76134 3585 76186
rect 3289 76132 3345 76134
rect 3369 76132 3425 76134
rect 3449 76132 3505 76134
rect 3529 76132 3585 76134
rect 7956 76186 8012 76188
rect 8036 76186 8092 76188
rect 8116 76186 8172 76188
rect 8196 76186 8252 76188
rect 7956 76134 7982 76186
rect 7982 76134 8012 76186
rect 8036 76134 8046 76186
rect 8046 76134 8092 76186
rect 8116 76134 8162 76186
rect 8162 76134 8172 76186
rect 8196 76134 8226 76186
rect 8226 76134 8252 76186
rect 7956 76132 8012 76134
rect 8036 76132 8092 76134
rect 8116 76132 8172 76134
rect 8196 76132 8252 76134
rect 5622 75642 5678 75644
rect 5702 75642 5758 75644
rect 5782 75642 5838 75644
rect 5862 75642 5918 75644
rect 5622 75590 5648 75642
rect 5648 75590 5678 75642
rect 5702 75590 5712 75642
rect 5712 75590 5758 75642
rect 5782 75590 5828 75642
rect 5828 75590 5838 75642
rect 5862 75590 5892 75642
rect 5892 75590 5918 75642
rect 5622 75588 5678 75590
rect 5702 75588 5758 75590
rect 5782 75588 5838 75590
rect 5862 75588 5918 75590
rect 10289 75642 10345 75644
rect 10369 75642 10425 75644
rect 10449 75642 10505 75644
rect 10529 75642 10585 75644
rect 10289 75590 10315 75642
rect 10315 75590 10345 75642
rect 10369 75590 10379 75642
rect 10379 75590 10425 75642
rect 10449 75590 10495 75642
rect 10495 75590 10505 75642
rect 10529 75590 10559 75642
rect 10559 75590 10585 75642
rect 10289 75588 10345 75590
rect 10369 75588 10425 75590
rect 10449 75588 10505 75590
rect 10529 75588 10585 75590
rect 3289 75098 3345 75100
rect 3369 75098 3425 75100
rect 3449 75098 3505 75100
rect 3529 75098 3585 75100
rect 3289 75046 3315 75098
rect 3315 75046 3345 75098
rect 3369 75046 3379 75098
rect 3379 75046 3425 75098
rect 3449 75046 3495 75098
rect 3495 75046 3505 75098
rect 3529 75046 3559 75098
rect 3559 75046 3585 75098
rect 3289 75044 3345 75046
rect 3369 75044 3425 75046
rect 3449 75044 3505 75046
rect 3529 75044 3585 75046
rect 7956 75098 8012 75100
rect 8036 75098 8092 75100
rect 8116 75098 8172 75100
rect 8196 75098 8252 75100
rect 7956 75046 7982 75098
rect 7982 75046 8012 75098
rect 8036 75046 8046 75098
rect 8046 75046 8092 75098
rect 8116 75046 8162 75098
rect 8162 75046 8172 75098
rect 8196 75046 8226 75098
rect 8226 75046 8252 75098
rect 7956 75044 8012 75046
rect 8036 75044 8092 75046
rect 8116 75044 8172 75046
rect 8196 75044 8252 75046
rect 110 74840 166 74896
rect 5622 74554 5678 74556
rect 5702 74554 5758 74556
rect 5782 74554 5838 74556
rect 5862 74554 5918 74556
rect 5622 74502 5648 74554
rect 5648 74502 5678 74554
rect 5702 74502 5712 74554
rect 5712 74502 5758 74554
rect 5782 74502 5828 74554
rect 5828 74502 5838 74554
rect 5862 74502 5892 74554
rect 5892 74502 5918 74554
rect 5622 74500 5678 74502
rect 5702 74500 5758 74502
rect 5782 74500 5838 74502
rect 5862 74500 5918 74502
rect 10289 74554 10345 74556
rect 10369 74554 10425 74556
rect 10449 74554 10505 74556
rect 10529 74554 10585 74556
rect 10289 74502 10315 74554
rect 10315 74502 10345 74554
rect 10369 74502 10379 74554
rect 10379 74502 10425 74554
rect 10449 74502 10495 74554
rect 10495 74502 10505 74554
rect 10529 74502 10559 74554
rect 10559 74502 10585 74554
rect 10289 74500 10345 74502
rect 10369 74500 10425 74502
rect 10449 74500 10505 74502
rect 10529 74500 10585 74502
rect 3289 74010 3345 74012
rect 3369 74010 3425 74012
rect 3449 74010 3505 74012
rect 3529 74010 3585 74012
rect 3289 73958 3315 74010
rect 3315 73958 3345 74010
rect 3369 73958 3379 74010
rect 3379 73958 3425 74010
rect 3449 73958 3495 74010
rect 3495 73958 3505 74010
rect 3529 73958 3559 74010
rect 3559 73958 3585 74010
rect 3289 73956 3345 73958
rect 3369 73956 3425 73958
rect 3449 73956 3505 73958
rect 3529 73956 3585 73958
rect 7956 74010 8012 74012
rect 8036 74010 8092 74012
rect 8116 74010 8172 74012
rect 8196 74010 8252 74012
rect 7956 73958 7982 74010
rect 7982 73958 8012 74010
rect 8036 73958 8046 74010
rect 8046 73958 8092 74010
rect 8116 73958 8162 74010
rect 8162 73958 8172 74010
rect 8196 73958 8226 74010
rect 8226 73958 8252 74010
rect 7956 73956 8012 73958
rect 8036 73956 8092 73958
rect 8116 73956 8172 73958
rect 8196 73956 8252 73958
rect 5622 73466 5678 73468
rect 5702 73466 5758 73468
rect 5782 73466 5838 73468
rect 5862 73466 5918 73468
rect 5622 73414 5648 73466
rect 5648 73414 5678 73466
rect 5702 73414 5712 73466
rect 5712 73414 5758 73466
rect 5782 73414 5828 73466
rect 5828 73414 5838 73466
rect 5862 73414 5892 73466
rect 5892 73414 5918 73466
rect 5622 73412 5678 73414
rect 5702 73412 5758 73414
rect 5782 73412 5838 73414
rect 5862 73412 5918 73414
rect 10289 73466 10345 73468
rect 10369 73466 10425 73468
rect 10449 73466 10505 73468
rect 10529 73466 10585 73468
rect 10289 73414 10315 73466
rect 10315 73414 10345 73466
rect 10369 73414 10379 73466
rect 10379 73414 10425 73466
rect 10449 73414 10495 73466
rect 10495 73414 10505 73466
rect 10529 73414 10559 73466
rect 10559 73414 10585 73466
rect 10289 73412 10345 73414
rect 10369 73412 10425 73414
rect 10449 73412 10505 73414
rect 10529 73412 10585 73414
rect 3289 72922 3345 72924
rect 3369 72922 3425 72924
rect 3449 72922 3505 72924
rect 3529 72922 3585 72924
rect 3289 72870 3315 72922
rect 3315 72870 3345 72922
rect 3369 72870 3379 72922
rect 3379 72870 3425 72922
rect 3449 72870 3495 72922
rect 3495 72870 3505 72922
rect 3529 72870 3559 72922
rect 3559 72870 3585 72922
rect 3289 72868 3345 72870
rect 3369 72868 3425 72870
rect 3449 72868 3505 72870
rect 3529 72868 3585 72870
rect 7956 72922 8012 72924
rect 8036 72922 8092 72924
rect 8116 72922 8172 72924
rect 8196 72922 8252 72924
rect 7956 72870 7982 72922
rect 7982 72870 8012 72922
rect 8036 72870 8046 72922
rect 8046 72870 8092 72922
rect 8116 72870 8162 72922
rect 8162 72870 8172 72922
rect 8196 72870 8226 72922
rect 8226 72870 8252 72922
rect 7956 72868 8012 72870
rect 8036 72868 8092 72870
rect 8116 72868 8172 72870
rect 8196 72868 8252 72870
rect 5622 72378 5678 72380
rect 5702 72378 5758 72380
rect 5782 72378 5838 72380
rect 5862 72378 5918 72380
rect 5622 72326 5648 72378
rect 5648 72326 5678 72378
rect 5702 72326 5712 72378
rect 5712 72326 5758 72378
rect 5782 72326 5828 72378
rect 5828 72326 5838 72378
rect 5862 72326 5892 72378
rect 5892 72326 5918 72378
rect 5622 72324 5678 72326
rect 5702 72324 5758 72326
rect 5782 72324 5838 72326
rect 5862 72324 5918 72326
rect 10289 72378 10345 72380
rect 10369 72378 10425 72380
rect 10449 72378 10505 72380
rect 10529 72378 10585 72380
rect 10289 72326 10315 72378
rect 10315 72326 10345 72378
rect 10369 72326 10379 72378
rect 10379 72326 10425 72378
rect 10449 72326 10495 72378
rect 10495 72326 10505 72378
rect 10529 72326 10559 72378
rect 10559 72326 10585 72378
rect 10289 72324 10345 72326
rect 10369 72324 10425 72326
rect 10449 72324 10505 72326
rect 10529 72324 10585 72326
rect 3289 71834 3345 71836
rect 3369 71834 3425 71836
rect 3449 71834 3505 71836
rect 3529 71834 3585 71836
rect 3289 71782 3315 71834
rect 3315 71782 3345 71834
rect 3369 71782 3379 71834
rect 3379 71782 3425 71834
rect 3449 71782 3495 71834
rect 3495 71782 3505 71834
rect 3529 71782 3559 71834
rect 3559 71782 3585 71834
rect 3289 71780 3345 71782
rect 3369 71780 3425 71782
rect 3449 71780 3505 71782
rect 3529 71780 3585 71782
rect 7956 71834 8012 71836
rect 8036 71834 8092 71836
rect 8116 71834 8172 71836
rect 8196 71834 8252 71836
rect 7956 71782 7982 71834
rect 7982 71782 8012 71834
rect 8036 71782 8046 71834
rect 8046 71782 8092 71834
rect 8116 71782 8162 71834
rect 8162 71782 8172 71834
rect 8196 71782 8226 71834
rect 8226 71782 8252 71834
rect 7956 71780 8012 71782
rect 8036 71780 8092 71782
rect 8116 71780 8172 71782
rect 8196 71780 8252 71782
rect 110 71576 166 71632
rect 5622 71290 5678 71292
rect 5702 71290 5758 71292
rect 5782 71290 5838 71292
rect 5862 71290 5918 71292
rect 5622 71238 5648 71290
rect 5648 71238 5678 71290
rect 5702 71238 5712 71290
rect 5712 71238 5758 71290
rect 5782 71238 5828 71290
rect 5828 71238 5838 71290
rect 5862 71238 5892 71290
rect 5892 71238 5918 71290
rect 5622 71236 5678 71238
rect 5702 71236 5758 71238
rect 5782 71236 5838 71238
rect 5862 71236 5918 71238
rect 10289 71290 10345 71292
rect 10369 71290 10425 71292
rect 10449 71290 10505 71292
rect 10529 71290 10585 71292
rect 10289 71238 10315 71290
rect 10315 71238 10345 71290
rect 10369 71238 10379 71290
rect 10379 71238 10425 71290
rect 10449 71238 10495 71290
rect 10495 71238 10505 71290
rect 10529 71238 10559 71290
rect 10559 71238 10585 71290
rect 10289 71236 10345 71238
rect 10369 71236 10425 71238
rect 10449 71236 10505 71238
rect 10529 71236 10585 71238
rect 3289 70746 3345 70748
rect 3369 70746 3425 70748
rect 3449 70746 3505 70748
rect 3529 70746 3585 70748
rect 3289 70694 3315 70746
rect 3315 70694 3345 70746
rect 3369 70694 3379 70746
rect 3379 70694 3425 70746
rect 3449 70694 3495 70746
rect 3495 70694 3505 70746
rect 3529 70694 3559 70746
rect 3559 70694 3585 70746
rect 3289 70692 3345 70694
rect 3369 70692 3425 70694
rect 3449 70692 3505 70694
rect 3529 70692 3585 70694
rect 7956 70746 8012 70748
rect 8036 70746 8092 70748
rect 8116 70746 8172 70748
rect 8196 70746 8252 70748
rect 7956 70694 7982 70746
rect 7982 70694 8012 70746
rect 8036 70694 8046 70746
rect 8046 70694 8092 70746
rect 8116 70694 8162 70746
rect 8162 70694 8172 70746
rect 8196 70694 8226 70746
rect 8226 70694 8252 70746
rect 7956 70692 8012 70694
rect 8036 70692 8092 70694
rect 8116 70692 8172 70694
rect 8196 70692 8252 70694
rect 5622 70202 5678 70204
rect 5702 70202 5758 70204
rect 5782 70202 5838 70204
rect 5862 70202 5918 70204
rect 5622 70150 5648 70202
rect 5648 70150 5678 70202
rect 5702 70150 5712 70202
rect 5712 70150 5758 70202
rect 5782 70150 5828 70202
rect 5828 70150 5838 70202
rect 5862 70150 5892 70202
rect 5892 70150 5918 70202
rect 5622 70148 5678 70150
rect 5702 70148 5758 70150
rect 5782 70148 5838 70150
rect 5862 70148 5918 70150
rect 10289 70202 10345 70204
rect 10369 70202 10425 70204
rect 10449 70202 10505 70204
rect 10529 70202 10585 70204
rect 10289 70150 10315 70202
rect 10315 70150 10345 70202
rect 10369 70150 10379 70202
rect 10379 70150 10425 70202
rect 10449 70150 10495 70202
rect 10495 70150 10505 70202
rect 10529 70150 10559 70202
rect 10559 70150 10585 70202
rect 10289 70148 10345 70150
rect 10369 70148 10425 70150
rect 10449 70148 10505 70150
rect 10529 70148 10585 70150
rect 3289 69658 3345 69660
rect 3369 69658 3425 69660
rect 3449 69658 3505 69660
rect 3529 69658 3585 69660
rect 3289 69606 3315 69658
rect 3315 69606 3345 69658
rect 3369 69606 3379 69658
rect 3379 69606 3425 69658
rect 3449 69606 3495 69658
rect 3495 69606 3505 69658
rect 3529 69606 3559 69658
rect 3559 69606 3585 69658
rect 3289 69604 3345 69606
rect 3369 69604 3425 69606
rect 3449 69604 3505 69606
rect 3529 69604 3585 69606
rect 7956 69658 8012 69660
rect 8036 69658 8092 69660
rect 8116 69658 8172 69660
rect 8196 69658 8252 69660
rect 7956 69606 7982 69658
rect 7982 69606 8012 69658
rect 8036 69606 8046 69658
rect 8046 69606 8092 69658
rect 8116 69606 8162 69658
rect 8162 69606 8172 69658
rect 8196 69606 8226 69658
rect 8226 69606 8252 69658
rect 7956 69604 8012 69606
rect 8036 69604 8092 69606
rect 8116 69604 8172 69606
rect 8196 69604 8252 69606
rect 5622 69114 5678 69116
rect 5702 69114 5758 69116
rect 5782 69114 5838 69116
rect 5862 69114 5918 69116
rect 5622 69062 5648 69114
rect 5648 69062 5678 69114
rect 5702 69062 5712 69114
rect 5712 69062 5758 69114
rect 5782 69062 5828 69114
rect 5828 69062 5838 69114
rect 5862 69062 5892 69114
rect 5892 69062 5918 69114
rect 5622 69060 5678 69062
rect 5702 69060 5758 69062
rect 5782 69060 5838 69062
rect 5862 69060 5918 69062
rect 10289 69114 10345 69116
rect 10369 69114 10425 69116
rect 10449 69114 10505 69116
rect 10529 69114 10585 69116
rect 10289 69062 10315 69114
rect 10315 69062 10345 69114
rect 10369 69062 10379 69114
rect 10379 69062 10425 69114
rect 10449 69062 10495 69114
rect 10495 69062 10505 69114
rect 10529 69062 10559 69114
rect 10559 69062 10585 69114
rect 10289 69060 10345 69062
rect 10369 69060 10425 69062
rect 10449 69060 10505 69062
rect 10529 69060 10585 69062
rect 3289 68570 3345 68572
rect 3369 68570 3425 68572
rect 3449 68570 3505 68572
rect 3529 68570 3585 68572
rect 3289 68518 3315 68570
rect 3315 68518 3345 68570
rect 3369 68518 3379 68570
rect 3379 68518 3425 68570
rect 3449 68518 3495 68570
rect 3495 68518 3505 68570
rect 3529 68518 3559 68570
rect 3559 68518 3585 68570
rect 3289 68516 3345 68518
rect 3369 68516 3425 68518
rect 3449 68516 3505 68518
rect 3529 68516 3585 68518
rect 7956 68570 8012 68572
rect 8036 68570 8092 68572
rect 8116 68570 8172 68572
rect 8196 68570 8252 68572
rect 7956 68518 7982 68570
rect 7982 68518 8012 68570
rect 8036 68518 8046 68570
rect 8046 68518 8092 68570
rect 8116 68518 8162 68570
rect 8162 68518 8172 68570
rect 8196 68518 8226 68570
rect 8226 68518 8252 68570
rect 7956 68516 8012 68518
rect 8036 68516 8092 68518
rect 8116 68516 8172 68518
rect 8196 68516 8252 68518
rect 5622 68026 5678 68028
rect 5702 68026 5758 68028
rect 5782 68026 5838 68028
rect 5862 68026 5918 68028
rect 5622 67974 5648 68026
rect 5648 67974 5678 68026
rect 5702 67974 5712 68026
rect 5712 67974 5758 68026
rect 5782 67974 5828 68026
rect 5828 67974 5838 68026
rect 5862 67974 5892 68026
rect 5892 67974 5918 68026
rect 5622 67972 5678 67974
rect 5702 67972 5758 67974
rect 5782 67972 5838 67974
rect 5862 67972 5918 67974
rect 10289 68026 10345 68028
rect 10369 68026 10425 68028
rect 10449 68026 10505 68028
rect 10529 68026 10585 68028
rect 10289 67974 10315 68026
rect 10315 67974 10345 68026
rect 10369 67974 10379 68026
rect 10379 67974 10425 68026
rect 10449 67974 10495 68026
rect 10495 67974 10505 68026
rect 10529 67974 10559 68026
rect 10559 67974 10585 68026
rect 10289 67972 10345 67974
rect 10369 67972 10425 67974
rect 10449 67972 10505 67974
rect 10529 67972 10585 67974
rect 3289 67482 3345 67484
rect 3369 67482 3425 67484
rect 3449 67482 3505 67484
rect 3529 67482 3585 67484
rect 3289 67430 3315 67482
rect 3315 67430 3345 67482
rect 3369 67430 3379 67482
rect 3379 67430 3425 67482
rect 3449 67430 3495 67482
rect 3495 67430 3505 67482
rect 3529 67430 3559 67482
rect 3559 67430 3585 67482
rect 3289 67428 3345 67430
rect 3369 67428 3425 67430
rect 3449 67428 3505 67430
rect 3529 67428 3585 67430
rect 7956 67482 8012 67484
rect 8036 67482 8092 67484
rect 8116 67482 8172 67484
rect 8196 67482 8252 67484
rect 7956 67430 7982 67482
rect 7982 67430 8012 67482
rect 8036 67430 8046 67482
rect 8046 67430 8092 67482
rect 8116 67430 8162 67482
rect 8162 67430 8172 67482
rect 8196 67430 8226 67482
rect 8226 67430 8252 67482
rect 7956 67428 8012 67430
rect 8036 67428 8092 67430
rect 8116 67428 8172 67430
rect 8196 67428 8252 67430
rect 5622 66938 5678 66940
rect 5702 66938 5758 66940
rect 5782 66938 5838 66940
rect 5862 66938 5918 66940
rect 5622 66886 5648 66938
rect 5648 66886 5678 66938
rect 5702 66886 5712 66938
rect 5712 66886 5758 66938
rect 5782 66886 5828 66938
rect 5828 66886 5838 66938
rect 5862 66886 5892 66938
rect 5892 66886 5918 66938
rect 5622 66884 5678 66886
rect 5702 66884 5758 66886
rect 5782 66884 5838 66886
rect 5862 66884 5918 66886
rect 10289 66938 10345 66940
rect 10369 66938 10425 66940
rect 10449 66938 10505 66940
rect 10529 66938 10585 66940
rect 10289 66886 10315 66938
rect 10315 66886 10345 66938
rect 10369 66886 10379 66938
rect 10379 66886 10425 66938
rect 10449 66886 10495 66938
rect 10495 66886 10505 66938
rect 10529 66886 10559 66938
rect 10559 66886 10585 66938
rect 10289 66884 10345 66886
rect 10369 66884 10425 66886
rect 10449 66884 10505 66886
rect 10529 66884 10585 66886
rect 3289 66394 3345 66396
rect 3369 66394 3425 66396
rect 3449 66394 3505 66396
rect 3529 66394 3585 66396
rect 3289 66342 3315 66394
rect 3315 66342 3345 66394
rect 3369 66342 3379 66394
rect 3379 66342 3425 66394
rect 3449 66342 3495 66394
rect 3495 66342 3505 66394
rect 3529 66342 3559 66394
rect 3559 66342 3585 66394
rect 3289 66340 3345 66342
rect 3369 66340 3425 66342
rect 3449 66340 3505 66342
rect 3529 66340 3585 66342
rect 7956 66394 8012 66396
rect 8036 66394 8092 66396
rect 8116 66394 8172 66396
rect 8196 66394 8252 66396
rect 7956 66342 7982 66394
rect 7982 66342 8012 66394
rect 8036 66342 8046 66394
rect 8046 66342 8092 66394
rect 8116 66342 8162 66394
rect 8162 66342 8172 66394
rect 8196 66342 8226 66394
rect 8226 66342 8252 66394
rect 7956 66340 8012 66342
rect 8036 66340 8092 66342
rect 8116 66340 8172 66342
rect 8196 66340 8252 66342
rect 5622 65850 5678 65852
rect 5702 65850 5758 65852
rect 5782 65850 5838 65852
rect 5862 65850 5918 65852
rect 5622 65798 5648 65850
rect 5648 65798 5678 65850
rect 5702 65798 5712 65850
rect 5712 65798 5758 65850
rect 5782 65798 5828 65850
rect 5828 65798 5838 65850
rect 5862 65798 5892 65850
rect 5892 65798 5918 65850
rect 5622 65796 5678 65798
rect 5702 65796 5758 65798
rect 5782 65796 5838 65798
rect 5862 65796 5918 65798
rect 3289 65306 3345 65308
rect 3369 65306 3425 65308
rect 3449 65306 3505 65308
rect 3529 65306 3585 65308
rect 3289 65254 3315 65306
rect 3315 65254 3345 65306
rect 3369 65254 3379 65306
rect 3379 65254 3425 65306
rect 3449 65254 3495 65306
rect 3495 65254 3505 65306
rect 3529 65254 3559 65306
rect 3559 65254 3585 65306
rect 3289 65252 3345 65254
rect 3369 65252 3425 65254
rect 3449 65252 3505 65254
rect 3529 65252 3585 65254
rect 7956 65306 8012 65308
rect 8036 65306 8092 65308
rect 8116 65306 8172 65308
rect 8196 65306 8252 65308
rect 7956 65254 7982 65306
rect 7982 65254 8012 65306
rect 8036 65254 8046 65306
rect 8046 65254 8092 65306
rect 8116 65254 8162 65306
rect 8162 65254 8172 65306
rect 8196 65254 8226 65306
rect 8226 65254 8252 65306
rect 7956 65252 8012 65254
rect 8036 65252 8092 65254
rect 8116 65252 8172 65254
rect 8196 65252 8252 65254
rect 5622 64762 5678 64764
rect 5702 64762 5758 64764
rect 5782 64762 5838 64764
rect 5862 64762 5918 64764
rect 5622 64710 5648 64762
rect 5648 64710 5678 64762
rect 5702 64710 5712 64762
rect 5712 64710 5758 64762
rect 5782 64710 5828 64762
rect 5828 64710 5838 64762
rect 5862 64710 5892 64762
rect 5892 64710 5918 64762
rect 5622 64708 5678 64710
rect 5702 64708 5758 64710
rect 5782 64708 5838 64710
rect 5862 64708 5918 64710
rect 3289 64218 3345 64220
rect 3369 64218 3425 64220
rect 3449 64218 3505 64220
rect 3529 64218 3585 64220
rect 3289 64166 3315 64218
rect 3315 64166 3345 64218
rect 3369 64166 3379 64218
rect 3379 64166 3425 64218
rect 3449 64166 3495 64218
rect 3495 64166 3505 64218
rect 3529 64166 3559 64218
rect 3559 64166 3585 64218
rect 3289 64164 3345 64166
rect 3369 64164 3425 64166
rect 3449 64164 3505 64166
rect 3529 64164 3585 64166
rect 7956 64218 8012 64220
rect 8036 64218 8092 64220
rect 8116 64218 8172 64220
rect 8196 64218 8252 64220
rect 7956 64166 7982 64218
rect 7982 64166 8012 64218
rect 8036 64166 8046 64218
rect 8046 64166 8092 64218
rect 8116 64166 8162 64218
rect 8162 64166 8172 64218
rect 8196 64166 8226 64218
rect 8226 64166 8252 64218
rect 7956 64164 8012 64166
rect 8036 64164 8092 64166
rect 8116 64164 8172 64166
rect 8196 64164 8252 64166
rect 5622 63674 5678 63676
rect 5702 63674 5758 63676
rect 5782 63674 5838 63676
rect 5862 63674 5918 63676
rect 5622 63622 5648 63674
rect 5648 63622 5678 63674
rect 5702 63622 5712 63674
rect 5712 63622 5758 63674
rect 5782 63622 5828 63674
rect 5828 63622 5838 63674
rect 5862 63622 5892 63674
rect 5892 63622 5918 63674
rect 5622 63620 5678 63622
rect 5702 63620 5758 63622
rect 5782 63620 5838 63622
rect 5862 63620 5918 63622
rect 3289 63130 3345 63132
rect 3369 63130 3425 63132
rect 3449 63130 3505 63132
rect 3529 63130 3585 63132
rect 3289 63078 3315 63130
rect 3315 63078 3345 63130
rect 3369 63078 3379 63130
rect 3379 63078 3425 63130
rect 3449 63078 3495 63130
rect 3495 63078 3505 63130
rect 3529 63078 3559 63130
rect 3559 63078 3585 63130
rect 3289 63076 3345 63078
rect 3369 63076 3425 63078
rect 3449 63076 3505 63078
rect 3529 63076 3585 63078
rect 7956 63130 8012 63132
rect 8036 63130 8092 63132
rect 8116 63130 8172 63132
rect 8196 63130 8252 63132
rect 7956 63078 7982 63130
rect 7982 63078 8012 63130
rect 8036 63078 8046 63130
rect 8046 63078 8092 63130
rect 8116 63078 8162 63130
rect 8162 63078 8172 63130
rect 8196 63078 8226 63130
rect 8226 63078 8252 63130
rect 7956 63076 8012 63078
rect 8036 63076 8092 63078
rect 8116 63076 8172 63078
rect 8196 63076 8252 63078
rect 5622 62586 5678 62588
rect 5702 62586 5758 62588
rect 5782 62586 5838 62588
rect 5862 62586 5918 62588
rect 5622 62534 5648 62586
rect 5648 62534 5678 62586
rect 5702 62534 5712 62586
rect 5712 62534 5758 62586
rect 5782 62534 5828 62586
rect 5828 62534 5838 62586
rect 5862 62534 5892 62586
rect 5892 62534 5918 62586
rect 5622 62532 5678 62534
rect 5702 62532 5758 62534
rect 5782 62532 5838 62534
rect 5862 62532 5918 62534
rect 3289 62042 3345 62044
rect 3369 62042 3425 62044
rect 3449 62042 3505 62044
rect 3529 62042 3585 62044
rect 3289 61990 3315 62042
rect 3315 61990 3345 62042
rect 3369 61990 3379 62042
rect 3379 61990 3425 62042
rect 3449 61990 3495 62042
rect 3495 61990 3505 62042
rect 3529 61990 3559 62042
rect 3559 61990 3585 62042
rect 3289 61988 3345 61990
rect 3369 61988 3425 61990
rect 3449 61988 3505 61990
rect 3529 61988 3585 61990
rect 7956 62042 8012 62044
rect 8036 62042 8092 62044
rect 8116 62042 8172 62044
rect 8196 62042 8252 62044
rect 7956 61990 7982 62042
rect 7982 61990 8012 62042
rect 8036 61990 8046 62042
rect 8046 61990 8092 62042
rect 8116 61990 8162 62042
rect 8162 61990 8172 62042
rect 8196 61990 8226 62042
rect 8226 61990 8252 62042
rect 7956 61988 8012 61990
rect 8036 61988 8092 61990
rect 8116 61988 8172 61990
rect 8196 61988 8252 61990
rect 5622 61498 5678 61500
rect 5702 61498 5758 61500
rect 5782 61498 5838 61500
rect 5862 61498 5918 61500
rect 5622 61446 5648 61498
rect 5648 61446 5678 61498
rect 5702 61446 5712 61498
rect 5712 61446 5758 61498
rect 5782 61446 5828 61498
rect 5828 61446 5838 61498
rect 5862 61446 5892 61498
rect 5892 61446 5918 61498
rect 5622 61444 5678 61446
rect 5702 61444 5758 61446
rect 5782 61444 5838 61446
rect 5862 61444 5918 61446
rect 110 61240 166 61296
rect 3289 60954 3345 60956
rect 3369 60954 3425 60956
rect 3449 60954 3505 60956
rect 3529 60954 3585 60956
rect 3289 60902 3315 60954
rect 3315 60902 3345 60954
rect 3369 60902 3379 60954
rect 3379 60902 3425 60954
rect 3449 60902 3495 60954
rect 3495 60902 3505 60954
rect 3529 60902 3559 60954
rect 3559 60902 3585 60954
rect 3289 60900 3345 60902
rect 3369 60900 3425 60902
rect 3449 60900 3505 60902
rect 3529 60900 3585 60902
rect 7956 60954 8012 60956
rect 8036 60954 8092 60956
rect 8116 60954 8172 60956
rect 8196 60954 8252 60956
rect 7956 60902 7982 60954
rect 7982 60902 8012 60954
rect 8036 60902 8046 60954
rect 8046 60902 8092 60954
rect 8116 60902 8162 60954
rect 8162 60902 8172 60954
rect 8196 60902 8226 60954
rect 8226 60902 8252 60954
rect 7956 60900 8012 60902
rect 8036 60900 8092 60902
rect 8116 60900 8172 60902
rect 8196 60900 8252 60902
rect 5622 60410 5678 60412
rect 5702 60410 5758 60412
rect 5782 60410 5838 60412
rect 5862 60410 5918 60412
rect 5622 60358 5648 60410
rect 5648 60358 5678 60410
rect 5702 60358 5712 60410
rect 5712 60358 5758 60410
rect 5782 60358 5828 60410
rect 5828 60358 5838 60410
rect 5862 60358 5892 60410
rect 5892 60358 5918 60410
rect 5622 60356 5678 60358
rect 5702 60356 5758 60358
rect 5782 60356 5838 60358
rect 5862 60356 5918 60358
rect 3289 59866 3345 59868
rect 3369 59866 3425 59868
rect 3449 59866 3505 59868
rect 3529 59866 3585 59868
rect 3289 59814 3315 59866
rect 3315 59814 3345 59866
rect 3369 59814 3379 59866
rect 3379 59814 3425 59866
rect 3449 59814 3495 59866
rect 3495 59814 3505 59866
rect 3529 59814 3559 59866
rect 3559 59814 3585 59866
rect 3289 59812 3345 59814
rect 3369 59812 3425 59814
rect 3449 59812 3505 59814
rect 3529 59812 3585 59814
rect 7956 59866 8012 59868
rect 8036 59866 8092 59868
rect 8116 59866 8172 59868
rect 8196 59866 8252 59868
rect 7956 59814 7982 59866
rect 7982 59814 8012 59866
rect 8036 59814 8046 59866
rect 8046 59814 8092 59866
rect 8116 59814 8162 59866
rect 8162 59814 8172 59866
rect 8196 59814 8226 59866
rect 8226 59814 8252 59866
rect 7956 59812 8012 59814
rect 8036 59812 8092 59814
rect 8116 59812 8172 59814
rect 8196 59812 8252 59814
rect 5622 59322 5678 59324
rect 5702 59322 5758 59324
rect 5782 59322 5838 59324
rect 5862 59322 5918 59324
rect 5622 59270 5648 59322
rect 5648 59270 5678 59322
rect 5702 59270 5712 59322
rect 5712 59270 5758 59322
rect 5782 59270 5828 59322
rect 5828 59270 5838 59322
rect 5862 59270 5892 59322
rect 5892 59270 5918 59322
rect 5622 59268 5678 59270
rect 5702 59268 5758 59270
rect 5782 59268 5838 59270
rect 5862 59268 5918 59270
rect 3289 58778 3345 58780
rect 3369 58778 3425 58780
rect 3449 58778 3505 58780
rect 3529 58778 3585 58780
rect 3289 58726 3315 58778
rect 3315 58726 3345 58778
rect 3369 58726 3379 58778
rect 3379 58726 3425 58778
rect 3449 58726 3495 58778
rect 3495 58726 3505 58778
rect 3529 58726 3559 58778
rect 3559 58726 3585 58778
rect 3289 58724 3345 58726
rect 3369 58724 3425 58726
rect 3449 58724 3505 58726
rect 3529 58724 3585 58726
rect 7956 58778 8012 58780
rect 8036 58778 8092 58780
rect 8116 58778 8172 58780
rect 8196 58778 8252 58780
rect 7956 58726 7982 58778
rect 7982 58726 8012 58778
rect 8036 58726 8046 58778
rect 8046 58726 8092 58778
rect 8116 58726 8162 58778
rect 8162 58726 8172 58778
rect 8196 58726 8226 58778
rect 8226 58726 8252 58778
rect 7956 58724 8012 58726
rect 8036 58724 8092 58726
rect 8116 58724 8172 58726
rect 8196 58724 8252 58726
rect 110 58520 166 58576
rect 5622 58234 5678 58236
rect 5702 58234 5758 58236
rect 5782 58234 5838 58236
rect 5862 58234 5918 58236
rect 5622 58182 5648 58234
rect 5648 58182 5678 58234
rect 5702 58182 5712 58234
rect 5712 58182 5758 58234
rect 5782 58182 5828 58234
rect 5828 58182 5838 58234
rect 5862 58182 5892 58234
rect 5892 58182 5918 58234
rect 5622 58180 5678 58182
rect 5702 58180 5758 58182
rect 5782 58180 5838 58182
rect 5862 58180 5918 58182
rect 3289 57690 3345 57692
rect 3369 57690 3425 57692
rect 3449 57690 3505 57692
rect 3529 57690 3585 57692
rect 3289 57638 3315 57690
rect 3315 57638 3345 57690
rect 3369 57638 3379 57690
rect 3379 57638 3425 57690
rect 3449 57638 3495 57690
rect 3495 57638 3505 57690
rect 3529 57638 3559 57690
rect 3559 57638 3585 57690
rect 3289 57636 3345 57638
rect 3369 57636 3425 57638
rect 3449 57636 3505 57638
rect 3529 57636 3585 57638
rect 7956 57690 8012 57692
rect 8036 57690 8092 57692
rect 8116 57690 8172 57692
rect 8196 57690 8252 57692
rect 7956 57638 7982 57690
rect 7982 57638 8012 57690
rect 8036 57638 8046 57690
rect 8046 57638 8092 57690
rect 8116 57638 8162 57690
rect 8162 57638 8172 57690
rect 8196 57638 8226 57690
rect 8226 57638 8252 57690
rect 7956 57636 8012 57638
rect 8036 57636 8092 57638
rect 8116 57636 8172 57638
rect 8196 57636 8252 57638
rect 5622 57146 5678 57148
rect 5702 57146 5758 57148
rect 5782 57146 5838 57148
rect 5862 57146 5918 57148
rect 5622 57094 5648 57146
rect 5648 57094 5678 57146
rect 5702 57094 5712 57146
rect 5712 57094 5758 57146
rect 5782 57094 5828 57146
rect 5828 57094 5838 57146
rect 5862 57094 5892 57146
rect 5892 57094 5918 57146
rect 5622 57092 5678 57094
rect 5702 57092 5758 57094
rect 5782 57092 5838 57094
rect 5862 57092 5918 57094
rect 3289 56602 3345 56604
rect 3369 56602 3425 56604
rect 3449 56602 3505 56604
rect 3529 56602 3585 56604
rect 3289 56550 3315 56602
rect 3315 56550 3345 56602
rect 3369 56550 3379 56602
rect 3379 56550 3425 56602
rect 3449 56550 3495 56602
rect 3495 56550 3505 56602
rect 3529 56550 3559 56602
rect 3559 56550 3585 56602
rect 3289 56548 3345 56550
rect 3369 56548 3425 56550
rect 3449 56548 3505 56550
rect 3529 56548 3585 56550
rect 7956 56602 8012 56604
rect 8036 56602 8092 56604
rect 8116 56602 8172 56604
rect 8196 56602 8252 56604
rect 7956 56550 7982 56602
rect 7982 56550 8012 56602
rect 8036 56550 8046 56602
rect 8046 56550 8092 56602
rect 8116 56550 8162 56602
rect 8162 56550 8172 56602
rect 8196 56550 8226 56602
rect 8226 56550 8252 56602
rect 7956 56548 8012 56550
rect 8036 56548 8092 56550
rect 8116 56548 8172 56550
rect 8196 56548 8252 56550
rect 5622 56058 5678 56060
rect 5702 56058 5758 56060
rect 5782 56058 5838 56060
rect 5862 56058 5918 56060
rect 5622 56006 5648 56058
rect 5648 56006 5678 56058
rect 5702 56006 5712 56058
rect 5712 56006 5758 56058
rect 5782 56006 5828 56058
rect 5828 56006 5838 56058
rect 5862 56006 5892 56058
rect 5892 56006 5918 56058
rect 5622 56004 5678 56006
rect 5702 56004 5758 56006
rect 5782 56004 5838 56006
rect 5862 56004 5918 56006
rect 3289 55514 3345 55516
rect 3369 55514 3425 55516
rect 3449 55514 3505 55516
rect 3529 55514 3585 55516
rect 3289 55462 3315 55514
rect 3315 55462 3345 55514
rect 3369 55462 3379 55514
rect 3379 55462 3425 55514
rect 3449 55462 3495 55514
rect 3495 55462 3505 55514
rect 3529 55462 3559 55514
rect 3559 55462 3585 55514
rect 3289 55460 3345 55462
rect 3369 55460 3425 55462
rect 3449 55460 3505 55462
rect 3529 55460 3585 55462
rect 7956 55514 8012 55516
rect 8036 55514 8092 55516
rect 8116 55514 8172 55516
rect 8196 55514 8252 55516
rect 7956 55462 7982 55514
rect 7982 55462 8012 55514
rect 8036 55462 8046 55514
rect 8046 55462 8092 55514
rect 8116 55462 8162 55514
rect 8162 55462 8172 55514
rect 8196 55462 8226 55514
rect 8226 55462 8252 55514
rect 7956 55460 8012 55462
rect 8036 55460 8092 55462
rect 8116 55460 8172 55462
rect 8196 55460 8252 55462
rect 5622 54970 5678 54972
rect 5702 54970 5758 54972
rect 5782 54970 5838 54972
rect 5862 54970 5918 54972
rect 5622 54918 5648 54970
rect 5648 54918 5678 54970
rect 5702 54918 5712 54970
rect 5712 54918 5758 54970
rect 5782 54918 5828 54970
rect 5828 54918 5838 54970
rect 5862 54918 5892 54970
rect 5892 54918 5918 54970
rect 5622 54916 5678 54918
rect 5702 54916 5758 54918
rect 5782 54916 5838 54918
rect 5862 54916 5918 54918
rect 3289 54426 3345 54428
rect 3369 54426 3425 54428
rect 3449 54426 3505 54428
rect 3529 54426 3585 54428
rect 3289 54374 3315 54426
rect 3315 54374 3345 54426
rect 3369 54374 3379 54426
rect 3379 54374 3425 54426
rect 3449 54374 3495 54426
rect 3495 54374 3505 54426
rect 3529 54374 3559 54426
rect 3559 54374 3585 54426
rect 3289 54372 3345 54374
rect 3369 54372 3425 54374
rect 3449 54372 3505 54374
rect 3529 54372 3585 54374
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 7982 54426
rect 7982 54374 8012 54426
rect 8036 54374 8046 54426
rect 8046 54374 8092 54426
rect 8116 54374 8162 54426
rect 8162 54374 8172 54426
rect 8196 54374 8226 54426
rect 8226 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 5622 53882 5678 53884
rect 5702 53882 5758 53884
rect 5782 53882 5838 53884
rect 5862 53882 5918 53884
rect 5622 53830 5648 53882
rect 5648 53830 5678 53882
rect 5702 53830 5712 53882
rect 5712 53830 5758 53882
rect 5782 53830 5828 53882
rect 5828 53830 5838 53882
rect 5862 53830 5892 53882
rect 5892 53830 5918 53882
rect 5622 53828 5678 53830
rect 5702 53828 5758 53830
rect 5782 53828 5838 53830
rect 5862 53828 5918 53830
rect 3289 53338 3345 53340
rect 3369 53338 3425 53340
rect 3449 53338 3505 53340
rect 3529 53338 3585 53340
rect 3289 53286 3315 53338
rect 3315 53286 3345 53338
rect 3369 53286 3379 53338
rect 3379 53286 3425 53338
rect 3449 53286 3495 53338
rect 3495 53286 3505 53338
rect 3529 53286 3559 53338
rect 3559 53286 3585 53338
rect 3289 53284 3345 53286
rect 3369 53284 3425 53286
rect 3449 53284 3505 53286
rect 3529 53284 3585 53286
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 7982 53338
rect 7982 53286 8012 53338
rect 8036 53286 8046 53338
rect 8046 53286 8092 53338
rect 8116 53286 8162 53338
rect 8162 53286 8172 53338
rect 8196 53286 8226 53338
rect 8226 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 5622 52794 5678 52796
rect 5702 52794 5758 52796
rect 5782 52794 5838 52796
rect 5862 52794 5918 52796
rect 5622 52742 5648 52794
rect 5648 52742 5678 52794
rect 5702 52742 5712 52794
rect 5712 52742 5758 52794
rect 5782 52742 5828 52794
rect 5828 52742 5838 52794
rect 5862 52742 5892 52794
rect 5892 52742 5918 52794
rect 5622 52740 5678 52742
rect 5702 52740 5758 52742
rect 5782 52740 5838 52742
rect 5862 52740 5918 52742
rect 3289 52250 3345 52252
rect 3369 52250 3425 52252
rect 3449 52250 3505 52252
rect 3529 52250 3585 52252
rect 3289 52198 3315 52250
rect 3315 52198 3345 52250
rect 3369 52198 3379 52250
rect 3379 52198 3425 52250
rect 3449 52198 3495 52250
rect 3495 52198 3505 52250
rect 3529 52198 3559 52250
rect 3559 52198 3585 52250
rect 3289 52196 3345 52198
rect 3369 52196 3425 52198
rect 3449 52196 3505 52198
rect 3529 52196 3585 52198
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 7982 52250
rect 7982 52198 8012 52250
rect 8036 52198 8046 52250
rect 8046 52198 8092 52250
rect 8116 52198 8162 52250
rect 8162 52198 8172 52250
rect 8196 52198 8226 52250
rect 8226 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 5622 51706 5678 51708
rect 5702 51706 5758 51708
rect 5782 51706 5838 51708
rect 5862 51706 5918 51708
rect 5622 51654 5648 51706
rect 5648 51654 5678 51706
rect 5702 51654 5712 51706
rect 5712 51654 5758 51706
rect 5782 51654 5828 51706
rect 5828 51654 5838 51706
rect 5862 51654 5892 51706
rect 5892 51654 5918 51706
rect 5622 51652 5678 51654
rect 5702 51652 5758 51654
rect 5782 51652 5838 51654
rect 5862 51652 5918 51654
rect 3289 51162 3345 51164
rect 3369 51162 3425 51164
rect 3449 51162 3505 51164
rect 3529 51162 3585 51164
rect 3289 51110 3315 51162
rect 3315 51110 3345 51162
rect 3369 51110 3379 51162
rect 3379 51110 3425 51162
rect 3449 51110 3495 51162
rect 3495 51110 3505 51162
rect 3529 51110 3559 51162
rect 3559 51110 3585 51162
rect 3289 51108 3345 51110
rect 3369 51108 3425 51110
rect 3449 51108 3505 51110
rect 3529 51108 3585 51110
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 7982 51162
rect 7982 51110 8012 51162
rect 8036 51110 8046 51162
rect 8046 51110 8092 51162
rect 8116 51110 8162 51162
rect 8162 51110 8172 51162
rect 8196 51110 8226 51162
rect 8226 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 5622 50618 5678 50620
rect 5702 50618 5758 50620
rect 5782 50618 5838 50620
rect 5862 50618 5918 50620
rect 5622 50566 5648 50618
rect 5648 50566 5678 50618
rect 5702 50566 5712 50618
rect 5712 50566 5758 50618
rect 5782 50566 5828 50618
rect 5828 50566 5838 50618
rect 5862 50566 5892 50618
rect 5892 50566 5918 50618
rect 5622 50564 5678 50566
rect 5702 50564 5758 50566
rect 5782 50564 5838 50566
rect 5862 50564 5918 50566
rect 3289 50074 3345 50076
rect 3369 50074 3425 50076
rect 3449 50074 3505 50076
rect 3529 50074 3585 50076
rect 3289 50022 3315 50074
rect 3315 50022 3345 50074
rect 3369 50022 3379 50074
rect 3379 50022 3425 50074
rect 3449 50022 3495 50074
rect 3495 50022 3505 50074
rect 3529 50022 3559 50074
rect 3559 50022 3585 50074
rect 3289 50020 3345 50022
rect 3369 50020 3425 50022
rect 3449 50020 3505 50022
rect 3529 50020 3585 50022
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 7982 50074
rect 7982 50022 8012 50074
rect 8036 50022 8046 50074
rect 8046 50022 8092 50074
rect 8116 50022 8162 50074
rect 8162 50022 8172 50074
rect 8196 50022 8226 50074
rect 8226 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 5622 49530 5678 49532
rect 5702 49530 5758 49532
rect 5782 49530 5838 49532
rect 5862 49530 5918 49532
rect 5622 49478 5648 49530
rect 5648 49478 5678 49530
rect 5702 49478 5712 49530
rect 5712 49478 5758 49530
rect 5782 49478 5828 49530
rect 5828 49478 5838 49530
rect 5862 49478 5892 49530
rect 5892 49478 5918 49530
rect 5622 49476 5678 49478
rect 5702 49476 5758 49478
rect 5782 49476 5838 49478
rect 5862 49476 5918 49478
rect 3289 48986 3345 48988
rect 3369 48986 3425 48988
rect 3449 48986 3505 48988
rect 3529 48986 3585 48988
rect 3289 48934 3315 48986
rect 3315 48934 3345 48986
rect 3369 48934 3379 48986
rect 3379 48934 3425 48986
rect 3449 48934 3495 48986
rect 3495 48934 3505 48986
rect 3529 48934 3559 48986
rect 3559 48934 3585 48986
rect 3289 48932 3345 48934
rect 3369 48932 3425 48934
rect 3449 48932 3505 48934
rect 3529 48932 3585 48934
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 7982 48986
rect 7982 48934 8012 48986
rect 8036 48934 8046 48986
rect 8046 48934 8092 48986
rect 8116 48934 8162 48986
rect 8162 48934 8172 48986
rect 8196 48934 8226 48986
rect 8226 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 5622 48442 5678 48444
rect 5702 48442 5758 48444
rect 5782 48442 5838 48444
rect 5862 48442 5918 48444
rect 5622 48390 5648 48442
rect 5648 48390 5678 48442
rect 5702 48390 5712 48442
rect 5712 48390 5758 48442
rect 5782 48390 5828 48442
rect 5828 48390 5838 48442
rect 5862 48390 5892 48442
rect 5892 48390 5918 48442
rect 5622 48388 5678 48390
rect 5702 48388 5758 48390
rect 5782 48388 5838 48390
rect 5862 48388 5918 48390
rect 3289 47898 3345 47900
rect 3369 47898 3425 47900
rect 3449 47898 3505 47900
rect 3529 47898 3585 47900
rect 3289 47846 3315 47898
rect 3315 47846 3345 47898
rect 3369 47846 3379 47898
rect 3379 47846 3425 47898
rect 3449 47846 3495 47898
rect 3495 47846 3505 47898
rect 3529 47846 3559 47898
rect 3559 47846 3585 47898
rect 3289 47844 3345 47846
rect 3369 47844 3425 47846
rect 3449 47844 3505 47846
rect 3529 47844 3585 47846
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 7982 47898
rect 7982 47846 8012 47898
rect 8036 47846 8046 47898
rect 8046 47846 8092 47898
rect 8116 47846 8162 47898
rect 8162 47846 8172 47898
rect 8196 47846 8226 47898
rect 8226 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 110 47640 166 47696
rect 5622 47354 5678 47356
rect 5702 47354 5758 47356
rect 5782 47354 5838 47356
rect 5862 47354 5918 47356
rect 5622 47302 5648 47354
rect 5648 47302 5678 47354
rect 5702 47302 5712 47354
rect 5712 47302 5758 47354
rect 5782 47302 5828 47354
rect 5828 47302 5838 47354
rect 5862 47302 5892 47354
rect 5892 47302 5918 47354
rect 5622 47300 5678 47302
rect 5702 47300 5758 47302
rect 5782 47300 5838 47302
rect 5862 47300 5918 47302
rect 3289 46810 3345 46812
rect 3369 46810 3425 46812
rect 3449 46810 3505 46812
rect 3529 46810 3585 46812
rect 3289 46758 3315 46810
rect 3315 46758 3345 46810
rect 3369 46758 3379 46810
rect 3379 46758 3425 46810
rect 3449 46758 3495 46810
rect 3495 46758 3505 46810
rect 3529 46758 3559 46810
rect 3559 46758 3585 46810
rect 3289 46756 3345 46758
rect 3369 46756 3425 46758
rect 3449 46756 3505 46758
rect 3529 46756 3585 46758
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 7982 46810
rect 7982 46758 8012 46810
rect 8036 46758 8046 46810
rect 8046 46758 8092 46810
rect 8116 46758 8162 46810
rect 8162 46758 8172 46810
rect 8196 46758 8226 46810
rect 8226 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 5622 46266 5678 46268
rect 5702 46266 5758 46268
rect 5782 46266 5838 46268
rect 5862 46266 5918 46268
rect 5622 46214 5648 46266
rect 5648 46214 5678 46266
rect 5702 46214 5712 46266
rect 5712 46214 5758 46266
rect 5782 46214 5828 46266
rect 5828 46214 5838 46266
rect 5862 46214 5892 46266
rect 5892 46214 5918 46266
rect 5622 46212 5678 46214
rect 5702 46212 5758 46214
rect 5782 46212 5838 46214
rect 5862 46212 5918 46214
rect 3289 45722 3345 45724
rect 3369 45722 3425 45724
rect 3449 45722 3505 45724
rect 3529 45722 3585 45724
rect 3289 45670 3315 45722
rect 3315 45670 3345 45722
rect 3369 45670 3379 45722
rect 3379 45670 3425 45722
rect 3449 45670 3495 45722
rect 3495 45670 3505 45722
rect 3529 45670 3559 45722
rect 3559 45670 3585 45722
rect 3289 45668 3345 45670
rect 3369 45668 3425 45670
rect 3449 45668 3505 45670
rect 3529 45668 3585 45670
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 7982 45722
rect 7982 45670 8012 45722
rect 8036 45670 8046 45722
rect 8046 45670 8092 45722
rect 8116 45670 8162 45722
rect 8162 45670 8172 45722
rect 8196 45670 8226 45722
rect 8226 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 5622 45178 5678 45180
rect 5702 45178 5758 45180
rect 5782 45178 5838 45180
rect 5862 45178 5918 45180
rect 5622 45126 5648 45178
rect 5648 45126 5678 45178
rect 5702 45126 5712 45178
rect 5712 45126 5758 45178
rect 5782 45126 5828 45178
rect 5828 45126 5838 45178
rect 5862 45126 5892 45178
rect 5892 45126 5918 45178
rect 5622 45124 5678 45126
rect 5702 45124 5758 45126
rect 5782 45124 5838 45126
rect 5862 45124 5918 45126
rect 110 44784 166 44840
rect 3289 44634 3345 44636
rect 3369 44634 3425 44636
rect 3449 44634 3505 44636
rect 3529 44634 3585 44636
rect 3289 44582 3315 44634
rect 3315 44582 3345 44634
rect 3369 44582 3379 44634
rect 3379 44582 3425 44634
rect 3449 44582 3495 44634
rect 3495 44582 3505 44634
rect 3529 44582 3559 44634
rect 3559 44582 3585 44634
rect 3289 44580 3345 44582
rect 3369 44580 3425 44582
rect 3449 44580 3505 44582
rect 3529 44580 3585 44582
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 7982 44634
rect 7982 44582 8012 44634
rect 8036 44582 8046 44634
rect 8046 44582 8092 44634
rect 8116 44582 8162 44634
rect 8162 44582 8172 44634
rect 8196 44582 8226 44634
rect 8226 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 5622 44090 5678 44092
rect 5702 44090 5758 44092
rect 5782 44090 5838 44092
rect 5862 44090 5918 44092
rect 5622 44038 5648 44090
rect 5648 44038 5678 44090
rect 5702 44038 5712 44090
rect 5712 44038 5758 44090
rect 5782 44038 5828 44090
rect 5828 44038 5838 44090
rect 5862 44038 5892 44090
rect 5892 44038 5918 44090
rect 5622 44036 5678 44038
rect 5702 44036 5758 44038
rect 5782 44036 5838 44038
rect 5862 44036 5918 44038
rect 3289 43546 3345 43548
rect 3369 43546 3425 43548
rect 3449 43546 3505 43548
rect 3529 43546 3585 43548
rect 3289 43494 3315 43546
rect 3315 43494 3345 43546
rect 3369 43494 3379 43546
rect 3379 43494 3425 43546
rect 3449 43494 3495 43546
rect 3495 43494 3505 43546
rect 3529 43494 3559 43546
rect 3559 43494 3585 43546
rect 3289 43492 3345 43494
rect 3369 43492 3425 43494
rect 3449 43492 3505 43494
rect 3529 43492 3585 43494
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 7982 43546
rect 7982 43494 8012 43546
rect 8036 43494 8046 43546
rect 8046 43494 8092 43546
rect 8116 43494 8162 43546
rect 8162 43494 8172 43546
rect 8196 43494 8226 43546
rect 8226 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 5622 43002 5678 43004
rect 5702 43002 5758 43004
rect 5782 43002 5838 43004
rect 5862 43002 5918 43004
rect 5622 42950 5648 43002
rect 5648 42950 5678 43002
rect 5702 42950 5712 43002
rect 5712 42950 5758 43002
rect 5782 42950 5828 43002
rect 5828 42950 5838 43002
rect 5862 42950 5892 43002
rect 5892 42950 5918 43002
rect 5622 42948 5678 42950
rect 5702 42948 5758 42950
rect 5782 42948 5838 42950
rect 5862 42948 5918 42950
rect 3289 42458 3345 42460
rect 3369 42458 3425 42460
rect 3449 42458 3505 42460
rect 3529 42458 3585 42460
rect 3289 42406 3315 42458
rect 3315 42406 3345 42458
rect 3369 42406 3379 42458
rect 3379 42406 3425 42458
rect 3449 42406 3495 42458
rect 3495 42406 3505 42458
rect 3529 42406 3559 42458
rect 3559 42406 3585 42458
rect 3289 42404 3345 42406
rect 3369 42404 3425 42406
rect 3449 42404 3505 42406
rect 3529 42404 3585 42406
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 7982 42458
rect 7982 42406 8012 42458
rect 8036 42406 8046 42458
rect 8046 42406 8092 42458
rect 8116 42406 8162 42458
rect 8162 42406 8172 42458
rect 8196 42406 8226 42458
rect 8226 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 5622 41914 5678 41916
rect 5702 41914 5758 41916
rect 5782 41914 5838 41916
rect 5862 41914 5918 41916
rect 5622 41862 5648 41914
rect 5648 41862 5678 41914
rect 5702 41862 5712 41914
rect 5712 41862 5758 41914
rect 5782 41862 5828 41914
rect 5828 41862 5838 41914
rect 5862 41862 5892 41914
rect 5892 41862 5918 41914
rect 5622 41860 5678 41862
rect 5702 41860 5758 41862
rect 5782 41860 5838 41862
rect 5862 41860 5918 41862
rect 3289 41370 3345 41372
rect 3369 41370 3425 41372
rect 3449 41370 3505 41372
rect 3529 41370 3585 41372
rect 3289 41318 3315 41370
rect 3315 41318 3345 41370
rect 3369 41318 3379 41370
rect 3379 41318 3425 41370
rect 3449 41318 3495 41370
rect 3495 41318 3505 41370
rect 3529 41318 3559 41370
rect 3559 41318 3585 41370
rect 3289 41316 3345 41318
rect 3369 41316 3425 41318
rect 3449 41316 3505 41318
rect 3529 41316 3585 41318
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 7982 41370
rect 7982 41318 8012 41370
rect 8036 41318 8046 41370
rect 8046 41318 8092 41370
rect 8116 41318 8162 41370
rect 8162 41318 8172 41370
rect 8196 41318 8226 41370
rect 8226 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 5622 40826 5678 40828
rect 5702 40826 5758 40828
rect 5782 40826 5838 40828
rect 5862 40826 5918 40828
rect 5622 40774 5648 40826
rect 5648 40774 5678 40826
rect 5702 40774 5712 40826
rect 5712 40774 5758 40826
rect 5782 40774 5828 40826
rect 5828 40774 5838 40826
rect 5862 40774 5892 40826
rect 5892 40774 5918 40826
rect 5622 40772 5678 40774
rect 5702 40772 5758 40774
rect 5782 40772 5838 40774
rect 5862 40772 5918 40774
rect 3289 40282 3345 40284
rect 3369 40282 3425 40284
rect 3449 40282 3505 40284
rect 3529 40282 3585 40284
rect 3289 40230 3315 40282
rect 3315 40230 3345 40282
rect 3369 40230 3379 40282
rect 3379 40230 3425 40282
rect 3449 40230 3495 40282
rect 3495 40230 3505 40282
rect 3529 40230 3559 40282
rect 3559 40230 3585 40282
rect 3289 40228 3345 40230
rect 3369 40228 3425 40230
rect 3449 40228 3505 40230
rect 3529 40228 3585 40230
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 7982 40282
rect 7982 40230 8012 40282
rect 8036 40230 8046 40282
rect 8046 40230 8092 40282
rect 8116 40230 8162 40282
rect 8162 40230 8172 40282
rect 8196 40230 8226 40282
rect 8226 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 5622 39738 5678 39740
rect 5702 39738 5758 39740
rect 5782 39738 5838 39740
rect 5862 39738 5918 39740
rect 5622 39686 5648 39738
rect 5648 39686 5678 39738
rect 5702 39686 5712 39738
rect 5712 39686 5758 39738
rect 5782 39686 5828 39738
rect 5828 39686 5838 39738
rect 5862 39686 5892 39738
rect 5892 39686 5918 39738
rect 5622 39684 5678 39686
rect 5702 39684 5758 39686
rect 5782 39684 5838 39686
rect 5862 39684 5918 39686
rect 3289 39194 3345 39196
rect 3369 39194 3425 39196
rect 3449 39194 3505 39196
rect 3529 39194 3585 39196
rect 3289 39142 3315 39194
rect 3315 39142 3345 39194
rect 3369 39142 3379 39194
rect 3379 39142 3425 39194
rect 3449 39142 3495 39194
rect 3495 39142 3505 39194
rect 3529 39142 3559 39194
rect 3559 39142 3585 39194
rect 3289 39140 3345 39142
rect 3369 39140 3425 39142
rect 3449 39140 3505 39142
rect 3529 39140 3585 39142
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 7982 39194
rect 7982 39142 8012 39194
rect 8036 39142 8046 39194
rect 8046 39142 8092 39194
rect 8116 39142 8162 39194
rect 8162 39142 8172 39194
rect 8196 39142 8226 39194
rect 8226 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 5622 38650 5678 38652
rect 5702 38650 5758 38652
rect 5782 38650 5838 38652
rect 5862 38650 5918 38652
rect 5622 38598 5648 38650
rect 5648 38598 5678 38650
rect 5702 38598 5712 38650
rect 5712 38598 5758 38650
rect 5782 38598 5828 38650
rect 5828 38598 5838 38650
rect 5862 38598 5892 38650
rect 5892 38598 5918 38650
rect 5622 38596 5678 38598
rect 5702 38596 5758 38598
rect 5782 38596 5838 38598
rect 5862 38596 5918 38598
rect 3289 38106 3345 38108
rect 3369 38106 3425 38108
rect 3449 38106 3505 38108
rect 3529 38106 3585 38108
rect 3289 38054 3315 38106
rect 3315 38054 3345 38106
rect 3369 38054 3379 38106
rect 3379 38054 3425 38106
rect 3449 38054 3495 38106
rect 3495 38054 3505 38106
rect 3529 38054 3559 38106
rect 3559 38054 3585 38106
rect 3289 38052 3345 38054
rect 3369 38052 3425 38054
rect 3449 38052 3505 38054
rect 3529 38052 3585 38054
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 7982 38106
rect 7982 38054 8012 38106
rect 8036 38054 8046 38106
rect 8046 38054 8092 38106
rect 8116 38054 8162 38106
rect 8162 38054 8172 38106
rect 8196 38054 8226 38106
rect 8226 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 5622 37562 5678 37564
rect 5702 37562 5758 37564
rect 5782 37562 5838 37564
rect 5862 37562 5918 37564
rect 5622 37510 5648 37562
rect 5648 37510 5678 37562
rect 5702 37510 5712 37562
rect 5712 37510 5758 37562
rect 5782 37510 5828 37562
rect 5828 37510 5838 37562
rect 5862 37510 5892 37562
rect 5892 37510 5918 37562
rect 5622 37508 5678 37510
rect 5702 37508 5758 37510
rect 5782 37508 5838 37510
rect 5862 37508 5918 37510
rect 3289 37018 3345 37020
rect 3369 37018 3425 37020
rect 3449 37018 3505 37020
rect 3529 37018 3585 37020
rect 3289 36966 3315 37018
rect 3315 36966 3345 37018
rect 3369 36966 3379 37018
rect 3379 36966 3425 37018
rect 3449 36966 3495 37018
rect 3495 36966 3505 37018
rect 3529 36966 3559 37018
rect 3559 36966 3585 37018
rect 3289 36964 3345 36966
rect 3369 36964 3425 36966
rect 3449 36964 3505 36966
rect 3529 36964 3585 36966
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 7982 37018
rect 7982 36966 8012 37018
rect 8036 36966 8046 37018
rect 8046 36966 8092 37018
rect 8116 36966 8162 37018
rect 8162 36966 8172 37018
rect 8196 36966 8226 37018
rect 8226 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 5622 36474 5678 36476
rect 5702 36474 5758 36476
rect 5782 36474 5838 36476
rect 5862 36474 5918 36476
rect 5622 36422 5648 36474
rect 5648 36422 5678 36474
rect 5702 36422 5712 36474
rect 5712 36422 5758 36474
rect 5782 36422 5828 36474
rect 5828 36422 5838 36474
rect 5862 36422 5892 36474
rect 5892 36422 5918 36474
rect 5622 36420 5678 36422
rect 5702 36420 5758 36422
rect 5782 36420 5838 36422
rect 5862 36420 5918 36422
rect 3289 35930 3345 35932
rect 3369 35930 3425 35932
rect 3449 35930 3505 35932
rect 3529 35930 3585 35932
rect 3289 35878 3315 35930
rect 3315 35878 3345 35930
rect 3369 35878 3379 35930
rect 3379 35878 3425 35930
rect 3449 35878 3495 35930
rect 3495 35878 3505 35930
rect 3529 35878 3559 35930
rect 3559 35878 3585 35930
rect 3289 35876 3345 35878
rect 3369 35876 3425 35878
rect 3449 35876 3505 35878
rect 3529 35876 3585 35878
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 7982 35930
rect 7982 35878 8012 35930
rect 8036 35878 8046 35930
rect 8046 35878 8092 35930
rect 8116 35878 8162 35930
rect 8162 35878 8172 35930
rect 8196 35878 8226 35930
rect 8226 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 5622 35386 5678 35388
rect 5702 35386 5758 35388
rect 5782 35386 5838 35388
rect 5862 35386 5918 35388
rect 5622 35334 5648 35386
rect 5648 35334 5678 35386
rect 5702 35334 5712 35386
rect 5712 35334 5758 35386
rect 5782 35334 5828 35386
rect 5828 35334 5838 35386
rect 5862 35334 5892 35386
rect 5892 35334 5918 35386
rect 5622 35332 5678 35334
rect 5702 35332 5758 35334
rect 5782 35332 5838 35334
rect 5862 35332 5918 35334
rect 3289 34842 3345 34844
rect 3369 34842 3425 34844
rect 3449 34842 3505 34844
rect 3529 34842 3585 34844
rect 3289 34790 3315 34842
rect 3315 34790 3345 34842
rect 3369 34790 3379 34842
rect 3379 34790 3425 34842
rect 3449 34790 3495 34842
rect 3495 34790 3505 34842
rect 3529 34790 3559 34842
rect 3559 34790 3585 34842
rect 3289 34788 3345 34790
rect 3369 34788 3425 34790
rect 3449 34788 3505 34790
rect 3529 34788 3585 34790
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 7982 34842
rect 7982 34790 8012 34842
rect 8036 34790 8046 34842
rect 8046 34790 8092 34842
rect 8116 34790 8162 34842
rect 8162 34790 8172 34842
rect 8196 34790 8226 34842
rect 8226 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 5622 34298 5678 34300
rect 5702 34298 5758 34300
rect 5782 34298 5838 34300
rect 5862 34298 5918 34300
rect 5622 34246 5648 34298
rect 5648 34246 5678 34298
rect 5702 34246 5712 34298
rect 5712 34246 5758 34298
rect 5782 34246 5828 34298
rect 5828 34246 5838 34298
rect 5862 34246 5892 34298
rect 5892 34246 5918 34298
rect 5622 34244 5678 34246
rect 5702 34244 5758 34246
rect 5782 34244 5838 34246
rect 5862 34244 5918 34246
rect 110 34040 166 34096
rect 3289 33754 3345 33756
rect 3369 33754 3425 33756
rect 3449 33754 3505 33756
rect 3529 33754 3585 33756
rect 3289 33702 3315 33754
rect 3315 33702 3345 33754
rect 3369 33702 3379 33754
rect 3379 33702 3425 33754
rect 3449 33702 3495 33754
rect 3495 33702 3505 33754
rect 3529 33702 3559 33754
rect 3559 33702 3585 33754
rect 3289 33700 3345 33702
rect 3369 33700 3425 33702
rect 3449 33700 3505 33702
rect 3529 33700 3585 33702
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 7982 33754
rect 7982 33702 8012 33754
rect 8036 33702 8046 33754
rect 8046 33702 8092 33754
rect 8116 33702 8162 33754
rect 8162 33702 8172 33754
rect 8196 33702 8226 33754
rect 8226 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 5622 33210 5678 33212
rect 5702 33210 5758 33212
rect 5782 33210 5838 33212
rect 5862 33210 5918 33212
rect 5622 33158 5648 33210
rect 5648 33158 5678 33210
rect 5702 33158 5712 33210
rect 5712 33158 5758 33210
rect 5782 33158 5828 33210
rect 5828 33158 5838 33210
rect 5862 33158 5892 33210
rect 5892 33158 5918 33210
rect 5622 33156 5678 33158
rect 5702 33156 5758 33158
rect 5782 33156 5838 33158
rect 5862 33156 5918 33158
rect 3289 32666 3345 32668
rect 3369 32666 3425 32668
rect 3449 32666 3505 32668
rect 3529 32666 3585 32668
rect 3289 32614 3315 32666
rect 3315 32614 3345 32666
rect 3369 32614 3379 32666
rect 3379 32614 3425 32666
rect 3449 32614 3495 32666
rect 3495 32614 3505 32666
rect 3529 32614 3559 32666
rect 3559 32614 3585 32666
rect 3289 32612 3345 32614
rect 3369 32612 3425 32614
rect 3449 32612 3505 32614
rect 3529 32612 3585 32614
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 7982 32666
rect 7982 32614 8012 32666
rect 8036 32614 8046 32666
rect 8046 32614 8092 32666
rect 8116 32614 8162 32666
rect 8162 32614 8172 32666
rect 8196 32614 8226 32666
rect 8226 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 5622 32122 5678 32124
rect 5702 32122 5758 32124
rect 5782 32122 5838 32124
rect 5862 32122 5918 32124
rect 5622 32070 5648 32122
rect 5648 32070 5678 32122
rect 5702 32070 5712 32122
rect 5712 32070 5758 32122
rect 5782 32070 5828 32122
rect 5828 32070 5838 32122
rect 5862 32070 5892 32122
rect 5892 32070 5918 32122
rect 5622 32068 5678 32070
rect 5702 32068 5758 32070
rect 5782 32068 5838 32070
rect 5862 32068 5918 32070
rect 3289 31578 3345 31580
rect 3369 31578 3425 31580
rect 3449 31578 3505 31580
rect 3529 31578 3585 31580
rect 3289 31526 3315 31578
rect 3315 31526 3345 31578
rect 3369 31526 3379 31578
rect 3379 31526 3425 31578
rect 3449 31526 3495 31578
rect 3495 31526 3505 31578
rect 3529 31526 3559 31578
rect 3559 31526 3585 31578
rect 3289 31524 3345 31526
rect 3369 31524 3425 31526
rect 3449 31524 3505 31526
rect 3529 31524 3585 31526
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 7982 31578
rect 7982 31526 8012 31578
rect 8036 31526 8046 31578
rect 8046 31526 8092 31578
rect 8116 31526 8162 31578
rect 8162 31526 8172 31578
rect 8196 31526 8226 31578
rect 8226 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 110 31184 166 31240
rect 5622 31034 5678 31036
rect 5702 31034 5758 31036
rect 5782 31034 5838 31036
rect 5862 31034 5918 31036
rect 5622 30982 5648 31034
rect 5648 30982 5678 31034
rect 5702 30982 5712 31034
rect 5712 30982 5758 31034
rect 5782 30982 5828 31034
rect 5828 30982 5838 31034
rect 5862 30982 5892 31034
rect 5892 30982 5918 31034
rect 5622 30980 5678 30982
rect 5702 30980 5758 30982
rect 5782 30980 5838 30982
rect 5862 30980 5918 30982
rect 3289 30490 3345 30492
rect 3369 30490 3425 30492
rect 3449 30490 3505 30492
rect 3529 30490 3585 30492
rect 3289 30438 3315 30490
rect 3315 30438 3345 30490
rect 3369 30438 3379 30490
rect 3379 30438 3425 30490
rect 3449 30438 3495 30490
rect 3495 30438 3505 30490
rect 3529 30438 3559 30490
rect 3559 30438 3585 30490
rect 3289 30436 3345 30438
rect 3369 30436 3425 30438
rect 3449 30436 3505 30438
rect 3529 30436 3585 30438
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 7982 30490
rect 7982 30438 8012 30490
rect 8036 30438 8046 30490
rect 8046 30438 8092 30490
rect 8116 30438 8162 30490
rect 8162 30438 8172 30490
rect 8196 30438 8226 30490
rect 8226 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 5622 29946 5678 29948
rect 5702 29946 5758 29948
rect 5782 29946 5838 29948
rect 5862 29946 5918 29948
rect 5622 29894 5648 29946
rect 5648 29894 5678 29946
rect 5702 29894 5712 29946
rect 5712 29894 5758 29946
rect 5782 29894 5828 29946
rect 5828 29894 5838 29946
rect 5862 29894 5892 29946
rect 5892 29894 5918 29946
rect 5622 29892 5678 29894
rect 5702 29892 5758 29894
rect 5782 29892 5838 29894
rect 5862 29892 5918 29894
rect 3289 29402 3345 29404
rect 3369 29402 3425 29404
rect 3449 29402 3505 29404
rect 3529 29402 3585 29404
rect 3289 29350 3315 29402
rect 3315 29350 3345 29402
rect 3369 29350 3379 29402
rect 3379 29350 3425 29402
rect 3449 29350 3495 29402
rect 3495 29350 3505 29402
rect 3529 29350 3559 29402
rect 3559 29350 3585 29402
rect 3289 29348 3345 29350
rect 3369 29348 3425 29350
rect 3449 29348 3505 29350
rect 3529 29348 3585 29350
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 7982 29402
rect 7982 29350 8012 29402
rect 8036 29350 8046 29402
rect 8046 29350 8092 29402
rect 8116 29350 8162 29402
rect 8162 29350 8172 29402
rect 8196 29350 8226 29402
rect 8226 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 5622 28858 5678 28860
rect 5702 28858 5758 28860
rect 5782 28858 5838 28860
rect 5862 28858 5918 28860
rect 5622 28806 5648 28858
rect 5648 28806 5678 28858
rect 5702 28806 5712 28858
rect 5712 28806 5758 28858
rect 5782 28806 5828 28858
rect 5828 28806 5838 28858
rect 5862 28806 5892 28858
rect 5892 28806 5918 28858
rect 5622 28804 5678 28806
rect 5702 28804 5758 28806
rect 5782 28804 5838 28806
rect 5862 28804 5918 28806
rect 3289 28314 3345 28316
rect 3369 28314 3425 28316
rect 3449 28314 3505 28316
rect 3529 28314 3585 28316
rect 3289 28262 3315 28314
rect 3315 28262 3345 28314
rect 3369 28262 3379 28314
rect 3379 28262 3425 28314
rect 3449 28262 3495 28314
rect 3495 28262 3505 28314
rect 3529 28262 3559 28314
rect 3559 28262 3585 28314
rect 3289 28260 3345 28262
rect 3369 28260 3425 28262
rect 3449 28260 3505 28262
rect 3529 28260 3585 28262
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 7982 28314
rect 7982 28262 8012 28314
rect 8036 28262 8046 28314
rect 8046 28262 8092 28314
rect 8116 28262 8162 28314
rect 8162 28262 8172 28314
rect 8196 28262 8226 28314
rect 8226 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 5622 27770 5678 27772
rect 5702 27770 5758 27772
rect 5782 27770 5838 27772
rect 5862 27770 5918 27772
rect 5622 27718 5648 27770
rect 5648 27718 5678 27770
rect 5702 27718 5712 27770
rect 5712 27718 5758 27770
rect 5782 27718 5828 27770
rect 5828 27718 5838 27770
rect 5862 27718 5892 27770
rect 5892 27718 5918 27770
rect 5622 27716 5678 27718
rect 5702 27716 5758 27718
rect 5782 27716 5838 27718
rect 5862 27716 5918 27718
rect 3289 27226 3345 27228
rect 3369 27226 3425 27228
rect 3449 27226 3505 27228
rect 3529 27226 3585 27228
rect 3289 27174 3315 27226
rect 3315 27174 3345 27226
rect 3369 27174 3379 27226
rect 3379 27174 3425 27226
rect 3449 27174 3495 27226
rect 3495 27174 3505 27226
rect 3529 27174 3559 27226
rect 3559 27174 3585 27226
rect 3289 27172 3345 27174
rect 3369 27172 3425 27174
rect 3449 27172 3505 27174
rect 3529 27172 3585 27174
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 7982 27226
rect 7982 27174 8012 27226
rect 8036 27174 8046 27226
rect 8046 27174 8092 27226
rect 8116 27174 8162 27226
rect 8162 27174 8172 27226
rect 8196 27174 8226 27226
rect 8226 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 5622 26682 5678 26684
rect 5702 26682 5758 26684
rect 5782 26682 5838 26684
rect 5862 26682 5918 26684
rect 5622 26630 5648 26682
rect 5648 26630 5678 26682
rect 5702 26630 5712 26682
rect 5712 26630 5758 26682
rect 5782 26630 5828 26682
rect 5828 26630 5838 26682
rect 5862 26630 5892 26682
rect 5892 26630 5918 26682
rect 5622 26628 5678 26630
rect 5702 26628 5758 26630
rect 5782 26628 5838 26630
rect 5862 26628 5918 26630
rect 3289 26138 3345 26140
rect 3369 26138 3425 26140
rect 3449 26138 3505 26140
rect 3529 26138 3585 26140
rect 3289 26086 3315 26138
rect 3315 26086 3345 26138
rect 3369 26086 3379 26138
rect 3379 26086 3425 26138
rect 3449 26086 3495 26138
rect 3495 26086 3505 26138
rect 3529 26086 3559 26138
rect 3559 26086 3585 26138
rect 3289 26084 3345 26086
rect 3369 26084 3425 26086
rect 3449 26084 3505 26086
rect 3529 26084 3585 26086
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 7982 26138
rect 7982 26086 8012 26138
rect 8036 26086 8046 26138
rect 8046 26086 8092 26138
rect 8116 26086 8162 26138
rect 8162 26086 8172 26138
rect 8196 26086 8226 26138
rect 8226 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 5622 25594 5678 25596
rect 5702 25594 5758 25596
rect 5782 25594 5838 25596
rect 5862 25594 5918 25596
rect 5622 25542 5648 25594
rect 5648 25542 5678 25594
rect 5702 25542 5712 25594
rect 5712 25542 5758 25594
rect 5782 25542 5828 25594
rect 5828 25542 5838 25594
rect 5862 25542 5892 25594
rect 5892 25542 5918 25594
rect 5622 25540 5678 25542
rect 5702 25540 5758 25542
rect 5782 25540 5838 25542
rect 5862 25540 5918 25542
rect 3289 25050 3345 25052
rect 3369 25050 3425 25052
rect 3449 25050 3505 25052
rect 3529 25050 3585 25052
rect 3289 24998 3315 25050
rect 3315 24998 3345 25050
rect 3369 24998 3379 25050
rect 3379 24998 3425 25050
rect 3449 24998 3495 25050
rect 3495 24998 3505 25050
rect 3529 24998 3559 25050
rect 3559 24998 3585 25050
rect 3289 24996 3345 24998
rect 3369 24996 3425 24998
rect 3449 24996 3505 24998
rect 3529 24996 3585 24998
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 7982 25050
rect 7982 24998 8012 25050
rect 8036 24998 8046 25050
rect 8046 24998 8092 25050
rect 8116 24998 8162 25050
rect 8162 24998 8172 25050
rect 8196 24998 8226 25050
rect 8226 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 5622 24506 5678 24508
rect 5702 24506 5758 24508
rect 5782 24506 5838 24508
rect 5862 24506 5918 24508
rect 5622 24454 5648 24506
rect 5648 24454 5678 24506
rect 5702 24454 5712 24506
rect 5712 24454 5758 24506
rect 5782 24454 5828 24506
rect 5828 24454 5838 24506
rect 5862 24454 5892 24506
rect 5892 24454 5918 24506
rect 5622 24452 5678 24454
rect 5702 24452 5758 24454
rect 5782 24452 5838 24454
rect 5862 24452 5918 24454
rect 3289 23962 3345 23964
rect 3369 23962 3425 23964
rect 3449 23962 3505 23964
rect 3529 23962 3585 23964
rect 3289 23910 3315 23962
rect 3315 23910 3345 23962
rect 3369 23910 3379 23962
rect 3379 23910 3425 23962
rect 3449 23910 3495 23962
rect 3495 23910 3505 23962
rect 3529 23910 3559 23962
rect 3559 23910 3585 23962
rect 3289 23908 3345 23910
rect 3369 23908 3425 23910
rect 3449 23908 3505 23910
rect 3529 23908 3585 23910
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 7982 23962
rect 7982 23910 8012 23962
rect 8036 23910 8046 23962
rect 8046 23910 8092 23962
rect 8116 23910 8162 23962
rect 8162 23910 8172 23962
rect 8196 23910 8226 23962
rect 8226 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 5622 23418 5678 23420
rect 5702 23418 5758 23420
rect 5782 23418 5838 23420
rect 5862 23418 5918 23420
rect 5622 23366 5648 23418
rect 5648 23366 5678 23418
rect 5702 23366 5712 23418
rect 5712 23366 5758 23418
rect 5782 23366 5828 23418
rect 5828 23366 5838 23418
rect 5862 23366 5892 23418
rect 5892 23366 5918 23418
rect 5622 23364 5678 23366
rect 5702 23364 5758 23366
rect 5782 23364 5838 23366
rect 5862 23364 5918 23366
rect 3289 22874 3345 22876
rect 3369 22874 3425 22876
rect 3449 22874 3505 22876
rect 3529 22874 3585 22876
rect 3289 22822 3315 22874
rect 3315 22822 3345 22874
rect 3369 22822 3379 22874
rect 3379 22822 3425 22874
rect 3449 22822 3495 22874
rect 3495 22822 3505 22874
rect 3529 22822 3559 22874
rect 3559 22822 3585 22874
rect 3289 22820 3345 22822
rect 3369 22820 3425 22822
rect 3449 22820 3505 22822
rect 3529 22820 3585 22822
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 7982 22874
rect 7982 22822 8012 22874
rect 8036 22822 8046 22874
rect 8046 22822 8092 22874
rect 8116 22822 8162 22874
rect 8162 22822 8172 22874
rect 8196 22822 8226 22874
rect 8226 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 5622 22330 5678 22332
rect 5702 22330 5758 22332
rect 5782 22330 5838 22332
rect 5862 22330 5918 22332
rect 5622 22278 5648 22330
rect 5648 22278 5678 22330
rect 5702 22278 5712 22330
rect 5712 22278 5758 22330
rect 5782 22278 5828 22330
rect 5828 22278 5838 22330
rect 5862 22278 5892 22330
rect 5892 22278 5918 22330
rect 5622 22276 5678 22278
rect 5702 22276 5758 22278
rect 5782 22276 5838 22278
rect 5862 22276 5918 22278
rect 3289 21786 3345 21788
rect 3369 21786 3425 21788
rect 3449 21786 3505 21788
rect 3529 21786 3585 21788
rect 3289 21734 3315 21786
rect 3315 21734 3345 21786
rect 3369 21734 3379 21786
rect 3379 21734 3425 21786
rect 3449 21734 3495 21786
rect 3495 21734 3505 21786
rect 3529 21734 3559 21786
rect 3559 21734 3585 21786
rect 3289 21732 3345 21734
rect 3369 21732 3425 21734
rect 3449 21732 3505 21734
rect 3529 21732 3585 21734
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 7982 21786
rect 7982 21734 8012 21786
rect 8036 21734 8046 21786
rect 8046 21734 8092 21786
rect 8116 21734 8162 21786
rect 8162 21734 8172 21786
rect 8196 21734 8226 21786
rect 8226 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 5622 21242 5678 21244
rect 5702 21242 5758 21244
rect 5782 21242 5838 21244
rect 5862 21242 5918 21244
rect 5622 21190 5648 21242
rect 5648 21190 5678 21242
rect 5702 21190 5712 21242
rect 5712 21190 5758 21242
rect 5782 21190 5828 21242
rect 5828 21190 5838 21242
rect 5862 21190 5892 21242
rect 5892 21190 5918 21242
rect 5622 21188 5678 21190
rect 5702 21188 5758 21190
rect 5782 21188 5838 21190
rect 5862 21188 5918 21190
rect 3289 20698 3345 20700
rect 3369 20698 3425 20700
rect 3449 20698 3505 20700
rect 3529 20698 3585 20700
rect 3289 20646 3315 20698
rect 3315 20646 3345 20698
rect 3369 20646 3379 20698
rect 3379 20646 3425 20698
rect 3449 20646 3495 20698
rect 3495 20646 3505 20698
rect 3529 20646 3559 20698
rect 3559 20646 3585 20698
rect 3289 20644 3345 20646
rect 3369 20644 3425 20646
rect 3449 20644 3505 20646
rect 3529 20644 3585 20646
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 7982 20698
rect 7982 20646 8012 20698
rect 8036 20646 8046 20698
rect 8046 20646 8092 20698
rect 8116 20646 8162 20698
rect 8162 20646 8172 20698
rect 8196 20646 8226 20698
rect 8226 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 110 20440 166 20496
rect 5622 20154 5678 20156
rect 5702 20154 5758 20156
rect 5782 20154 5838 20156
rect 5862 20154 5918 20156
rect 5622 20102 5648 20154
rect 5648 20102 5678 20154
rect 5702 20102 5712 20154
rect 5712 20102 5758 20154
rect 5782 20102 5828 20154
rect 5828 20102 5838 20154
rect 5862 20102 5892 20154
rect 5892 20102 5918 20154
rect 5622 20100 5678 20102
rect 5702 20100 5758 20102
rect 5782 20100 5838 20102
rect 5862 20100 5918 20102
rect 3289 19610 3345 19612
rect 3369 19610 3425 19612
rect 3449 19610 3505 19612
rect 3529 19610 3585 19612
rect 3289 19558 3315 19610
rect 3315 19558 3345 19610
rect 3369 19558 3379 19610
rect 3379 19558 3425 19610
rect 3449 19558 3495 19610
rect 3495 19558 3505 19610
rect 3529 19558 3559 19610
rect 3559 19558 3585 19610
rect 3289 19556 3345 19558
rect 3369 19556 3425 19558
rect 3449 19556 3505 19558
rect 3529 19556 3585 19558
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 7982 19610
rect 7982 19558 8012 19610
rect 8036 19558 8046 19610
rect 8046 19558 8092 19610
rect 8116 19558 8162 19610
rect 8162 19558 8172 19610
rect 8196 19558 8226 19610
rect 8226 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 5622 19066 5678 19068
rect 5702 19066 5758 19068
rect 5782 19066 5838 19068
rect 5862 19066 5918 19068
rect 5622 19014 5648 19066
rect 5648 19014 5678 19066
rect 5702 19014 5712 19066
rect 5712 19014 5758 19066
rect 5782 19014 5828 19066
rect 5828 19014 5838 19066
rect 5862 19014 5892 19066
rect 5892 19014 5918 19066
rect 5622 19012 5678 19014
rect 5702 19012 5758 19014
rect 5782 19012 5838 19014
rect 5862 19012 5918 19014
rect 3289 18522 3345 18524
rect 3369 18522 3425 18524
rect 3449 18522 3505 18524
rect 3529 18522 3585 18524
rect 3289 18470 3315 18522
rect 3315 18470 3345 18522
rect 3369 18470 3379 18522
rect 3379 18470 3425 18522
rect 3449 18470 3495 18522
rect 3495 18470 3505 18522
rect 3529 18470 3559 18522
rect 3559 18470 3585 18522
rect 3289 18468 3345 18470
rect 3369 18468 3425 18470
rect 3449 18468 3505 18470
rect 3529 18468 3585 18470
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 7982 18522
rect 7982 18470 8012 18522
rect 8036 18470 8046 18522
rect 8046 18470 8092 18522
rect 8116 18470 8162 18522
rect 8162 18470 8172 18522
rect 8196 18470 8226 18522
rect 8226 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 5622 17978 5678 17980
rect 5702 17978 5758 17980
rect 5782 17978 5838 17980
rect 5862 17978 5918 17980
rect 5622 17926 5648 17978
rect 5648 17926 5678 17978
rect 5702 17926 5712 17978
rect 5712 17926 5758 17978
rect 5782 17926 5828 17978
rect 5828 17926 5838 17978
rect 5862 17926 5892 17978
rect 5892 17926 5918 17978
rect 5622 17924 5678 17926
rect 5702 17924 5758 17926
rect 5782 17924 5838 17926
rect 5862 17924 5918 17926
rect 3289 17434 3345 17436
rect 3369 17434 3425 17436
rect 3449 17434 3505 17436
rect 3529 17434 3585 17436
rect 3289 17382 3315 17434
rect 3315 17382 3345 17434
rect 3369 17382 3379 17434
rect 3379 17382 3425 17434
rect 3449 17382 3495 17434
rect 3495 17382 3505 17434
rect 3529 17382 3559 17434
rect 3559 17382 3585 17434
rect 3289 17380 3345 17382
rect 3369 17380 3425 17382
rect 3449 17380 3505 17382
rect 3529 17380 3585 17382
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 7982 17434
rect 7982 17382 8012 17434
rect 8036 17382 8046 17434
rect 8046 17382 8092 17434
rect 8116 17382 8162 17434
rect 8162 17382 8172 17434
rect 8196 17382 8226 17434
rect 8226 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 110 17176 166 17232
rect 5622 16890 5678 16892
rect 5702 16890 5758 16892
rect 5782 16890 5838 16892
rect 5862 16890 5918 16892
rect 5622 16838 5648 16890
rect 5648 16838 5678 16890
rect 5702 16838 5712 16890
rect 5712 16838 5758 16890
rect 5782 16838 5828 16890
rect 5828 16838 5838 16890
rect 5862 16838 5892 16890
rect 5892 16838 5918 16890
rect 5622 16836 5678 16838
rect 5702 16836 5758 16838
rect 5782 16836 5838 16838
rect 5862 16836 5918 16838
rect 3289 16346 3345 16348
rect 3369 16346 3425 16348
rect 3449 16346 3505 16348
rect 3529 16346 3585 16348
rect 3289 16294 3315 16346
rect 3315 16294 3345 16346
rect 3369 16294 3379 16346
rect 3379 16294 3425 16346
rect 3449 16294 3495 16346
rect 3495 16294 3505 16346
rect 3529 16294 3559 16346
rect 3559 16294 3585 16346
rect 3289 16292 3345 16294
rect 3369 16292 3425 16294
rect 3449 16292 3505 16294
rect 3529 16292 3585 16294
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 7982 16346
rect 7982 16294 8012 16346
rect 8036 16294 8046 16346
rect 8046 16294 8092 16346
rect 8116 16294 8162 16346
rect 8162 16294 8172 16346
rect 8196 16294 8226 16346
rect 8226 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 5622 15802 5678 15804
rect 5702 15802 5758 15804
rect 5782 15802 5838 15804
rect 5862 15802 5918 15804
rect 5622 15750 5648 15802
rect 5648 15750 5678 15802
rect 5702 15750 5712 15802
rect 5712 15750 5758 15802
rect 5782 15750 5828 15802
rect 5828 15750 5838 15802
rect 5862 15750 5892 15802
rect 5892 15750 5918 15802
rect 5622 15748 5678 15750
rect 5702 15748 5758 15750
rect 5782 15748 5838 15750
rect 5862 15748 5918 15750
rect 3289 15258 3345 15260
rect 3369 15258 3425 15260
rect 3449 15258 3505 15260
rect 3529 15258 3585 15260
rect 3289 15206 3315 15258
rect 3315 15206 3345 15258
rect 3369 15206 3379 15258
rect 3379 15206 3425 15258
rect 3449 15206 3495 15258
rect 3495 15206 3505 15258
rect 3529 15206 3559 15258
rect 3559 15206 3585 15258
rect 3289 15204 3345 15206
rect 3369 15204 3425 15206
rect 3449 15204 3505 15206
rect 3529 15204 3585 15206
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 7982 15258
rect 7982 15206 8012 15258
rect 8036 15206 8046 15258
rect 8046 15206 8092 15258
rect 8116 15206 8162 15258
rect 8162 15206 8172 15258
rect 8196 15206 8226 15258
rect 8226 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 5622 14714 5678 14716
rect 5702 14714 5758 14716
rect 5782 14714 5838 14716
rect 5862 14714 5918 14716
rect 5622 14662 5648 14714
rect 5648 14662 5678 14714
rect 5702 14662 5712 14714
rect 5712 14662 5758 14714
rect 5782 14662 5828 14714
rect 5828 14662 5838 14714
rect 5862 14662 5892 14714
rect 5892 14662 5918 14714
rect 5622 14660 5678 14662
rect 5702 14660 5758 14662
rect 5782 14660 5838 14662
rect 5862 14660 5918 14662
rect 10289 65850 10345 65852
rect 10369 65850 10425 65852
rect 10449 65850 10505 65852
rect 10529 65850 10585 65852
rect 10289 65798 10315 65850
rect 10315 65798 10345 65850
rect 10369 65798 10379 65850
rect 10379 65798 10425 65850
rect 10449 65798 10495 65850
rect 10495 65798 10505 65850
rect 10529 65798 10559 65850
rect 10559 65798 10585 65850
rect 10289 65796 10345 65798
rect 10369 65796 10425 65798
rect 10449 65796 10505 65798
rect 10529 65796 10585 65798
rect 10289 64762 10345 64764
rect 10369 64762 10425 64764
rect 10449 64762 10505 64764
rect 10529 64762 10585 64764
rect 10289 64710 10315 64762
rect 10315 64710 10345 64762
rect 10369 64710 10379 64762
rect 10379 64710 10425 64762
rect 10449 64710 10495 64762
rect 10495 64710 10505 64762
rect 10529 64710 10559 64762
rect 10559 64710 10585 64762
rect 10289 64708 10345 64710
rect 10369 64708 10425 64710
rect 10449 64708 10505 64710
rect 10529 64708 10585 64710
rect 10289 63674 10345 63676
rect 10369 63674 10425 63676
rect 10449 63674 10505 63676
rect 10529 63674 10585 63676
rect 10289 63622 10315 63674
rect 10315 63622 10345 63674
rect 10369 63622 10379 63674
rect 10379 63622 10425 63674
rect 10449 63622 10495 63674
rect 10495 63622 10505 63674
rect 10529 63622 10559 63674
rect 10559 63622 10585 63674
rect 10289 63620 10345 63622
rect 10369 63620 10425 63622
rect 10449 63620 10505 63622
rect 10529 63620 10585 63622
rect 10289 62586 10345 62588
rect 10369 62586 10425 62588
rect 10449 62586 10505 62588
rect 10529 62586 10585 62588
rect 10289 62534 10315 62586
rect 10315 62534 10345 62586
rect 10369 62534 10379 62586
rect 10379 62534 10425 62586
rect 10449 62534 10495 62586
rect 10495 62534 10505 62586
rect 10529 62534 10559 62586
rect 10559 62534 10585 62586
rect 10289 62532 10345 62534
rect 10369 62532 10425 62534
rect 10449 62532 10505 62534
rect 10529 62532 10585 62534
rect 10289 61498 10345 61500
rect 10369 61498 10425 61500
rect 10449 61498 10505 61500
rect 10529 61498 10585 61500
rect 10289 61446 10315 61498
rect 10315 61446 10345 61498
rect 10369 61446 10379 61498
rect 10379 61446 10425 61498
rect 10449 61446 10495 61498
rect 10495 61446 10505 61498
rect 10529 61446 10559 61498
rect 10559 61446 10585 61498
rect 10289 61444 10345 61446
rect 10369 61444 10425 61446
rect 10449 61444 10505 61446
rect 10529 61444 10585 61446
rect 10289 60410 10345 60412
rect 10369 60410 10425 60412
rect 10449 60410 10505 60412
rect 10529 60410 10585 60412
rect 10289 60358 10315 60410
rect 10315 60358 10345 60410
rect 10369 60358 10379 60410
rect 10379 60358 10425 60410
rect 10449 60358 10495 60410
rect 10495 60358 10505 60410
rect 10529 60358 10559 60410
rect 10559 60358 10585 60410
rect 10289 60356 10345 60358
rect 10369 60356 10425 60358
rect 10449 60356 10505 60358
rect 10529 60356 10585 60358
rect 10289 59322 10345 59324
rect 10369 59322 10425 59324
rect 10449 59322 10505 59324
rect 10529 59322 10585 59324
rect 10289 59270 10315 59322
rect 10315 59270 10345 59322
rect 10369 59270 10379 59322
rect 10379 59270 10425 59322
rect 10449 59270 10495 59322
rect 10495 59270 10505 59322
rect 10529 59270 10559 59322
rect 10559 59270 10585 59322
rect 10289 59268 10345 59270
rect 10369 59268 10425 59270
rect 10449 59268 10505 59270
rect 10529 59268 10585 59270
rect 10289 58234 10345 58236
rect 10369 58234 10425 58236
rect 10449 58234 10505 58236
rect 10529 58234 10585 58236
rect 10289 58182 10315 58234
rect 10315 58182 10345 58234
rect 10369 58182 10379 58234
rect 10379 58182 10425 58234
rect 10449 58182 10495 58234
rect 10495 58182 10505 58234
rect 10529 58182 10559 58234
rect 10559 58182 10585 58234
rect 10289 58180 10345 58182
rect 10369 58180 10425 58182
rect 10449 58180 10505 58182
rect 10529 58180 10585 58182
rect 10289 57146 10345 57148
rect 10369 57146 10425 57148
rect 10449 57146 10505 57148
rect 10529 57146 10585 57148
rect 10289 57094 10315 57146
rect 10315 57094 10345 57146
rect 10369 57094 10379 57146
rect 10379 57094 10425 57146
rect 10449 57094 10495 57146
rect 10495 57094 10505 57146
rect 10529 57094 10559 57146
rect 10559 57094 10585 57146
rect 10289 57092 10345 57094
rect 10369 57092 10425 57094
rect 10449 57092 10505 57094
rect 10529 57092 10585 57094
rect 10289 56058 10345 56060
rect 10369 56058 10425 56060
rect 10449 56058 10505 56060
rect 10529 56058 10585 56060
rect 10289 56006 10315 56058
rect 10315 56006 10345 56058
rect 10369 56006 10379 56058
rect 10379 56006 10425 56058
rect 10449 56006 10495 56058
rect 10495 56006 10505 56058
rect 10529 56006 10559 56058
rect 10559 56006 10585 56058
rect 10289 56004 10345 56006
rect 10369 56004 10425 56006
rect 10449 56004 10505 56006
rect 10529 56004 10585 56006
rect 10289 54970 10345 54972
rect 10369 54970 10425 54972
rect 10449 54970 10505 54972
rect 10529 54970 10585 54972
rect 10289 54918 10315 54970
rect 10315 54918 10345 54970
rect 10369 54918 10379 54970
rect 10379 54918 10425 54970
rect 10449 54918 10495 54970
rect 10495 54918 10505 54970
rect 10529 54918 10559 54970
rect 10559 54918 10585 54970
rect 10289 54916 10345 54918
rect 10369 54916 10425 54918
rect 10449 54916 10505 54918
rect 10529 54916 10585 54918
rect 10289 53882 10345 53884
rect 10369 53882 10425 53884
rect 10449 53882 10505 53884
rect 10529 53882 10585 53884
rect 10289 53830 10315 53882
rect 10315 53830 10345 53882
rect 10369 53830 10379 53882
rect 10379 53830 10425 53882
rect 10449 53830 10495 53882
rect 10495 53830 10505 53882
rect 10529 53830 10559 53882
rect 10559 53830 10585 53882
rect 10289 53828 10345 53830
rect 10369 53828 10425 53830
rect 10449 53828 10505 53830
rect 10529 53828 10585 53830
rect 10289 52794 10345 52796
rect 10369 52794 10425 52796
rect 10449 52794 10505 52796
rect 10529 52794 10585 52796
rect 10289 52742 10315 52794
rect 10315 52742 10345 52794
rect 10369 52742 10379 52794
rect 10379 52742 10425 52794
rect 10449 52742 10495 52794
rect 10495 52742 10505 52794
rect 10529 52742 10559 52794
rect 10559 52742 10585 52794
rect 10289 52740 10345 52742
rect 10369 52740 10425 52742
rect 10449 52740 10505 52742
rect 10529 52740 10585 52742
rect 10289 51706 10345 51708
rect 10369 51706 10425 51708
rect 10449 51706 10505 51708
rect 10529 51706 10585 51708
rect 10289 51654 10315 51706
rect 10315 51654 10345 51706
rect 10369 51654 10379 51706
rect 10379 51654 10425 51706
rect 10449 51654 10495 51706
rect 10495 51654 10505 51706
rect 10529 51654 10559 51706
rect 10559 51654 10585 51706
rect 10289 51652 10345 51654
rect 10369 51652 10425 51654
rect 10449 51652 10505 51654
rect 10529 51652 10585 51654
rect 10289 50618 10345 50620
rect 10369 50618 10425 50620
rect 10449 50618 10505 50620
rect 10529 50618 10585 50620
rect 10289 50566 10315 50618
rect 10315 50566 10345 50618
rect 10369 50566 10379 50618
rect 10379 50566 10425 50618
rect 10449 50566 10495 50618
rect 10495 50566 10505 50618
rect 10529 50566 10559 50618
rect 10559 50566 10585 50618
rect 10289 50564 10345 50566
rect 10369 50564 10425 50566
rect 10449 50564 10505 50566
rect 10529 50564 10585 50566
rect 10289 49530 10345 49532
rect 10369 49530 10425 49532
rect 10449 49530 10505 49532
rect 10529 49530 10585 49532
rect 10289 49478 10315 49530
rect 10315 49478 10345 49530
rect 10369 49478 10379 49530
rect 10379 49478 10425 49530
rect 10449 49478 10495 49530
rect 10495 49478 10505 49530
rect 10529 49478 10559 49530
rect 10559 49478 10585 49530
rect 10289 49476 10345 49478
rect 10369 49476 10425 49478
rect 10449 49476 10505 49478
rect 10529 49476 10585 49478
rect 10289 48442 10345 48444
rect 10369 48442 10425 48444
rect 10449 48442 10505 48444
rect 10529 48442 10585 48444
rect 10289 48390 10315 48442
rect 10315 48390 10345 48442
rect 10369 48390 10379 48442
rect 10379 48390 10425 48442
rect 10449 48390 10495 48442
rect 10495 48390 10505 48442
rect 10529 48390 10559 48442
rect 10559 48390 10585 48442
rect 10289 48388 10345 48390
rect 10369 48388 10425 48390
rect 10449 48388 10505 48390
rect 10529 48388 10585 48390
rect 10289 47354 10345 47356
rect 10369 47354 10425 47356
rect 10449 47354 10505 47356
rect 10529 47354 10585 47356
rect 10289 47302 10315 47354
rect 10315 47302 10345 47354
rect 10369 47302 10379 47354
rect 10379 47302 10425 47354
rect 10449 47302 10495 47354
rect 10495 47302 10505 47354
rect 10529 47302 10559 47354
rect 10559 47302 10585 47354
rect 10289 47300 10345 47302
rect 10369 47300 10425 47302
rect 10449 47300 10505 47302
rect 10529 47300 10585 47302
rect 10289 46266 10345 46268
rect 10369 46266 10425 46268
rect 10449 46266 10505 46268
rect 10529 46266 10585 46268
rect 10289 46214 10315 46266
rect 10315 46214 10345 46266
rect 10369 46214 10379 46266
rect 10379 46214 10425 46266
rect 10449 46214 10495 46266
rect 10495 46214 10505 46266
rect 10529 46214 10559 46266
rect 10559 46214 10585 46266
rect 10289 46212 10345 46214
rect 10369 46212 10425 46214
rect 10449 46212 10505 46214
rect 10529 46212 10585 46214
rect 10289 45178 10345 45180
rect 10369 45178 10425 45180
rect 10449 45178 10505 45180
rect 10529 45178 10585 45180
rect 10289 45126 10315 45178
rect 10315 45126 10345 45178
rect 10369 45126 10379 45178
rect 10379 45126 10425 45178
rect 10449 45126 10495 45178
rect 10495 45126 10505 45178
rect 10529 45126 10559 45178
rect 10559 45126 10585 45178
rect 10289 45124 10345 45126
rect 10369 45124 10425 45126
rect 10449 45124 10505 45126
rect 10529 45124 10585 45126
rect 10782 44240 10838 44296
rect 10289 44090 10345 44092
rect 10369 44090 10425 44092
rect 10449 44090 10505 44092
rect 10529 44090 10585 44092
rect 10289 44038 10315 44090
rect 10315 44038 10345 44090
rect 10369 44038 10379 44090
rect 10379 44038 10425 44090
rect 10449 44038 10495 44090
rect 10495 44038 10505 44090
rect 10529 44038 10559 44090
rect 10559 44038 10585 44090
rect 10289 44036 10345 44038
rect 10369 44036 10425 44038
rect 10449 44036 10505 44038
rect 10529 44036 10585 44038
rect 10289 43002 10345 43004
rect 10369 43002 10425 43004
rect 10449 43002 10505 43004
rect 10529 43002 10585 43004
rect 10289 42950 10315 43002
rect 10315 42950 10345 43002
rect 10369 42950 10379 43002
rect 10379 42950 10425 43002
rect 10449 42950 10495 43002
rect 10495 42950 10505 43002
rect 10529 42950 10559 43002
rect 10559 42950 10585 43002
rect 10289 42948 10345 42950
rect 10369 42948 10425 42950
rect 10449 42948 10505 42950
rect 10529 42948 10585 42950
rect 10289 41914 10345 41916
rect 10369 41914 10425 41916
rect 10449 41914 10505 41916
rect 10529 41914 10585 41916
rect 10289 41862 10315 41914
rect 10315 41862 10345 41914
rect 10369 41862 10379 41914
rect 10379 41862 10425 41914
rect 10449 41862 10495 41914
rect 10495 41862 10505 41914
rect 10529 41862 10559 41914
rect 10559 41862 10585 41914
rect 10289 41860 10345 41862
rect 10369 41860 10425 41862
rect 10449 41860 10505 41862
rect 10529 41860 10585 41862
rect 10289 40826 10345 40828
rect 10369 40826 10425 40828
rect 10449 40826 10505 40828
rect 10529 40826 10585 40828
rect 10289 40774 10315 40826
rect 10315 40774 10345 40826
rect 10369 40774 10379 40826
rect 10379 40774 10425 40826
rect 10449 40774 10495 40826
rect 10495 40774 10505 40826
rect 10529 40774 10559 40826
rect 10559 40774 10585 40826
rect 10289 40772 10345 40774
rect 10369 40772 10425 40774
rect 10449 40772 10505 40774
rect 10529 40772 10585 40774
rect 10289 39738 10345 39740
rect 10369 39738 10425 39740
rect 10449 39738 10505 39740
rect 10529 39738 10585 39740
rect 10289 39686 10315 39738
rect 10315 39686 10345 39738
rect 10369 39686 10379 39738
rect 10379 39686 10425 39738
rect 10449 39686 10495 39738
rect 10495 39686 10505 39738
rect 10529 39686 10559 39738
rect 10559 39686 10585 39738
rect 10289 39684 10345 39686
rect 10369 39684 10425 39686
rect 10449 39684 10505 39686
rect 10529 39684 10585 39686
rect 10289 38650 10345 38652
rect 10369 38650 10425 38652
rect 10449 38650 10505 38652
rect 10529 38650 10585 38652
rect 10289 38598 10315 38650
rect 10315 38598 10345 38650
rect 10369 38598 10379 38650
rect 10379 38598 10425 38650
rect 10449 38598 10495 38650
rect 10495 38598 10505 38650
rect 10529 38598 10559 38650
rect 10559 38598 10585 38650
rect 10289 38596 10345 38598
rect 10369 38596 10425 38598
rect 10449 38596 10505 38598
rect 10529 38596 10585 38598
rect 10289 37562 10345 37564
rect 10369 37562 10425 37564
rect 10449 37562 10505 37564
rect 10529 37562 10585 37564
rect 10289 37510 10315 37562
rect 10315 37510 10345 37562
rect 10369 37510 10379 37562
rect 10379 37510 10425 37562
rect 10449 37510 10495 37562
rect 10495 37510 10505 37562
rect 10529 37510 10559 37562
rect 10559 37510 10585 37562
rect 10289 37508 10345 37510
rect 10369 37508 10425 37510
rect 10449 37508 10505 37510
rect 10529 37508 10585 37510
rect 10289 36474 10345 36476
rect 10369 36474 10425 36476
rect 10449 36474 10505 36476
rect 10529 36474 10585 36476
rect 10289 36422 10315 36474
rect 10315 36422 10345 36474
rect 10369 36422 10379 36474
rect 10379 36422 10425 36474
rect 10449 36422 10495 36474
rect 10495 36422 10505 36474
rect 10529 36422 10559 36474
rect 10559 36422 10585 36474
rect 10289 36420 10345 36422
rect 10369 36420 10425 36422
rect 10449 36420 10505 36422
rect 10529 36420 10585 36422
rect 10289 35386 10345 35388
rect 10369 35386 10425 35388
rect 10449 35386 10505 35388
rect 10529 35386 10585 35388
rect 10289 35334 10315 35386
rect 10315 35334 10345 35386
rect 10369 35334 10379 35386
rect 10379 35334 10425 35386
rect 10449 35334 10495 35386
rect 10495 35334 10505 35386
rect 10529 35334 10559 35386
rect 10559 35334 10585 35386
rect 10289 35332 10345 35334
rect 10369 35332 10425 35334
rect 10449 35332 10505 35334
rect 10529 35332 10585 35334
rect 10289 34298 10345 34300
rect 10369 34298 10425 34300
rect 10449 34298 10505 34300
rect 10529 34298 10585 34300
rect 10289 34246 10315 34298
rect 10315 34246 10345 34298
rect 10369 34246 10379 34298
rect 10379 34246 10425 34298
rect 10449 34246 10495 34298
rect 10495 34246 10505 34298
rect 10529 34246 10559 34298
rect 10559 34246 10585 34298
rect 10289 34244 10345 34246
rect 10369 34244 10425 34246
rect 10449 34244 10505 34246
rect 10529 34244 10585 34246
rect 10289 33210 10345 33212
rect 10369 33210 10425 33212
rect 10449 33210 10505 33212
rect 10529 33210 10585 33212
rect 10289 33158 10315 33210
rect 10315 33158 10345 33210
rect 10369 33158 10379 33210
rect 10379 33158 10425 33210
rect 10449 33158 10495 33210
rect 10495 33158 10505 33210
rect 10529 33158 10559 33210
rect 10559 33158 10585 33210
rect 10289 33156 10345 33158
rect 10369 33156 10425 33158
rect 10449 33156 10505 33158
rect 10529 33156 10585 33158
rect 10289 32122 10345 32124
rect 10369 32122 10425 32124
rect 10449 32122 10505 32124
rect 10529 32122 10585 32124
rect 10289 32070 10315 32122
rect 10315 32070 10345 32122
rect 10369 32070 10379 32122
rect 10379 32070 10425 32122
rect 10449 32070 10495 32122
rect 10495 32070 10505 32122
rect 10529 32070 10559 32122
rect 10559 32070 10585 32122
rect 10289 32068 10345 32070
rect 10369 32068 10425 32070
rect 10449 32068 10505 32070
rect 10529 32068 10585 32070
rect 10966 31184 11022 31240
rect 10289 31034 10345 31036
rect 10369 31034 10425 31036
rect 10449 31034 10505 31036
rect 10529 31034 10585 31036
rect 10289 30982 10315 31034
rect 10315 30982 10345 31034
rect 10369 30982 10379 31034
rect 10379 30982 10425 31034
rect 10449 30982 10495 31034
rect 10495 30982 10505 31034
rect 10529 30982 10559 31034
rect 10559 30982 10585 31034
rect 10289 30980 10345 30982
rect 10369 30980 10425 30982
rect 10449 30980 10505 30982
rect 10529 30980 10585 30982
rect 10782 30640 10838 30696
rect 10289 29946 10345 29948
rect 10369 29946 10425 29948
rect 10449 29946 10505 29948
rect 10529 29946 10585 29948
rect 10289 29894 10315 29946
rect 10315 29894 10345 29946
rect 10369 29894 10379 29946
rect 10379 29894 10425 29946
rect 10449 29894 10495 29946
rect 10495 29894 10505 29946
rect 10529 29894 10559 29946
rect 10559 29894 10585 29946
rect 10289 29892 10345 29894
rect 10369 29892 10425 29894
rect 10449 29892 10505 29894
rect 10529 29892 10585 29894
rect 10289 28858 10345 28860
rect 10369 28858 10425 28860
rect 10449 28858 10505 28860
rect 10529 28858 10585 28860
rect 10289 28806 10315 28858
rect 10315 28806 10345 28858
rect 10369 28806 10379 28858
rect 10379 28806 10425 28858
rect 10449 28806 10495 28858
rect 10495 28806 10505 28858
rect 10529 28806 10559 28858
rect 10559 28806 10585 28858
rect 10289 28804 10345 28806
rect 10369 28804 10425 28806
rect 10449 28804 10505 28806
rect 10529 28804 10585 28806
rect 10289 27770 10345 27772
rect 10369 27770 10425 27772
rect 10449 27770 10505 27772
rect 10529 27770 10585 27772
rect 10289 27718 10315 27770
rect 10315 27718 10345 27770
rect 10369 27718 10379 27770
rect 10379 27718 10425 27770
rect 10449 27718 10495 27770
rect 10495 27718 10505 27770
rect 10529 27718 10559 27770
rect 10559 27718 10585 27770
rect 10289 27716 10345 27718
rect 10369 27716 10425 27718
rect 10449 27716 10505 27718
rect 10529 27716 10585 27718
rect 10289 26682 10345 26684
rect 10369 26682 10425 26684
rect 10449 26682 10505 26684
rect 10529 26682 10585 26684
rect 10289 26630 10315 26682
rect 10315 26630 10345 26682
rect 10369 26630 10379 26682
rect 10379 26630 10425 26682
rect 10449 26630 10495 26682
rect 10495 26630 10505 26682
rect 10529 26630 10559 26682
rect 10559 26630 10585 26682
rect 10289 26628 10345 26630
rect 10369 26628 10425 26630
rect 10449 26628 10505 26630
rect 10529 26628 10585 26630
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10690 23840 10746 23896
rect 3289 14170 3345 14172
rect 3369 14170 3425 14172
rect 3449 14170 3505 14172
rect 3529 14170 3585 14172
rect 3289 14118 3315 14170
rect 3315 14118 3345 14170
rect 3369 14118 3379 14170
rect 3379 14118 3425 14170
rect 3449 14118 3495 14170
rect 3495 14118 3505 14170
rect 3529 14118 3559 14170
rect 3559 14118 3585 14170
rect 3289 14116 3345 14118
rect 3369 14116 3425 14118
rect 3449 14116 3505 14118
rect 3529 14116 3585 14118
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 7982 14170
rect 7982 14118 8012 14170
rect 8036 14118 8046 14170
rect 8046 14118 8092 14170
rect 8116 14118 8162 14170
rect 8162 14118 8172 14170
rect 8196 14118 8226 14170
rect 8226 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 5622 13626 5678 13628
rect 5702 13626 5758 13628
rect 5782 13626 5838 13628
rect 5862 13626 5918 13628
rect 5622 13574 5648 13626
rect 5648 13574 5678 13626
rect 5702 13574 5712 13626
rect 5712 13574 5758 13626
rect 5782 13574 5828 13626
rect 5828 13574 5838 13626
rect 5862 13574 5892 13626
rect 5892 13574 5918 13626
rect 5622 13572 5678 13574
rect 5702 13572 5758 13574
rect 5782 13572 5838 13574
rect 5862 13572 5918 13574
rect 3289 13082 3345 13084
rect 3369 13082 3425 13084
rect 3449 13082 3505 13084
rect 3529 13082 3585 13084
rect 3289 13030 3315 13082
rect 3315 13030 3345 13082
rect 3369 13030 3379 13082
rect 3379 13030 3425 13082
rect 3449 13030 3495 13082
rect 3495 13030 3505 13082
rect 3529 13030 3559 13082
rect 3559 13030 3585 13082
rect 3289 13028 3345 13030
rect 3369 13028 3425 13030
rect 3449 13028 3505 13030
rect 3529 13028 3585 13030
rect 110 6840 166 6896
rect 110 5616 166 5672
rect 5622 12538 5678 12540
rect 5702 12538 5758 12540
rect 5782 12538 5838 12540
rect 5862 12538 5918 12540
rect 5622 12486 5648 12538
rect 5648 12486 5678 12538
rect 5702 12486 5712 12538
rect 5712 12486 5758 12538
rect 5782 12486 5828 12538
rect 5828 12486 5838 12538
rect 5862 12486 5892 12538
rect 5892 12486 5918 12538
rect 5622 12484 5678 12486
rect 5702 12484 5758 12486
rect 5782 12484 5838 12486
rect 5862 12484 5918 12486
rect 3289 11994 3345 11996
rect 3369 11994 3425 11996
rect 3449 11994 3505 11996
rect 3529 11994 3585 11996
rect 3289 11942 3315 11994
rect 3315 11942 3345 11994
rect 3369 11942 3379 11994
rect 3379 11942 3425 11994
rect 3449 11942 3495 11994
rect 3495 11942 3505 11994
rect 3529 11942 3559 11994
rect 3559 11942 3585 11994
rect 3289 11940 3345 11942
rect 3369 11940 3425 11942
rect 3449 11940 3505 11942
rect 3529 11940 3585 11942
rect 5622 11450 5678 11452
rect 5702 11450 5758 11452
rect 5782 11450 5838 11452
rect 5862 11450 5918 11452
rect 5622 11398 5648 11450
rect 5648 11398 5678 11450
rect 5702 11398 5712 11450
rect 5712 11398 5758 11450
rect 5782 11398 5828 11450
rect 5828 11398 5838 11450
rect 5862 11398 5892 11450
rect 5892 11398 5918 11450
rect 5622 11396 5678 11398
rect 5702 11396 5758 11398
rect 5782 11396 5838 11398
rect 5862 11396 5918 11398
rect 3289 10906 3345 10908
rect 3369 10906 3425 10908
rect 3449 10906 3505 10908
rect 3529 10906 3585 10908
rect 3289 10854 3315 10906
rect 3315 10854 3345 10906
rect 3369 10854 3379 10906
rect 3379 10854 3425 10906
rect 3449 10854 3495 10906
rect 3495 10854 3505 10906
rect 3529 10854 3559 10906
rect 3559 10854 3585 10906
rect 3289 10852 3345 10854
rect 3369 10852 3425 10854
rect 3449 10852 3505 10854
rect 3529 10852 3585 10854
rect 5622 10362 5678 10364
rect 5702 10362 5758 10364
rect 5782 10362 5838 10364
rect 5862 10362 5918 10364
rect 5622 10310 5648 10362
rect 5648 10310 5678 10362
rect 5702 10310 5712 10362
rect 5712 10310 5758 10362
rect 5782 10310 5828 10362
rect 5828 10310 5838 10362
rect 5862 10310 5892 10362
rect 5892 10310 5918 10362
rect 5622 10308 5678 10310
rect 5702 10308 5758 10310
rect 5782 10308 5838 10310
rect 5862 10308 5918 10310
rect 3289 9818 3345 9820
rect 3369 9818 3425 9820
rect 3449 9818 3505 9820
rect 3529 9818 3585 9820
rect 3289 9766 3315 9818
rect 3315 9766 3345 9818
rect 3369 9766 3379 9818
rect 3379 9766 3425 9818
rect 3449 9766 3495 9818
rect 3495 9766 3505 9818
rect 3529 9766 3559 9818
rect 3559 9766 3585 9818
rect 3289 9764 3345 9766
rect 3369 9764 3425 9766
rect 3449 9764 3505 9766
rect 3529 9764 3585 9766
rect 5622 9274 5678 9276
rect 5702 9274 5758 9276
rect 5782 9274 5838 9276
rect 5862 9274 5918 9276
rect 5622 9222 5648 9274
rect 5648 9222 5678 9274
rect 5702 9222 5712 9274
rect 5712 9222 5758 9274
rect 5782 9222 5828 9274
rect 5828 9222 5838 9274
rect 5862 9222 5892 9274
rect 5892 9222 5918 9274
rect 5622 9220 5678 9222
rect 5702 9220 5758 9222
rect 5782 9220 5838 9222
rect 5862 9220 5918 9222
rect 3289 8730 3345 8732
rect 3369 8730 3425 8732
rect 3449 8730 3505 8732
rect 3529 8730 3585 8732
rect 3289 8678 3315 8730
rect 3315 8678 3345 8730
rect 3369 8678 3379 8730
rect 3379 8678 3425 8730
rect 3449 8678 3495 8730
rect 3495 8678 3505 8730
rect 3529 8678 3559 8730
rect 3559 8678 3585 8730
rect 3289 8676 3345 8678
rect 3369 8676 3425 8678
rect 3449 8676 3505 8678
rect 3529 8676 3585 8678
rect 5622 8186 5678 8188
rect 5702 8186 5758 8188
rect 5782 8186 5838 8188
rect 5862 8186 5918 8188
rect 5622 8134 5648 8186
rect 5648 8134 5678 8186
rect 5702 8134 5712 8186
rect 5712 8134 5758 8186
rect 5782 8134 5828 8186
rect 5828 8134 5838 8186
rect 5862 8134 5892 8186
rect 5892 8134 5918 8186
rect 5622 8132 5678 8134
rect 5702 8132 5758 8134
rect 5782 8132 5838 8134
rect 5862 8132 5918 8134
rect 3289 7642 3345 7644
rect 3369 7642 3425 7644
rect 3449 7642 3505 7644
rect 3529 7642 3585 7644
rect 3289 7590 3315 7642
rect 3315 7590 3345 7642
rect 3369 7590 3379 7642
rect 3379 7590 3425 7642
rect 3449 7590 3495 7642
rect 3495 7590 3505 7642
rect 3529 7590 3559 7642
rect 3559 7590 3585 7642
rect 3289 7588 3345 7590
rect 3369 7588 3425 7590
rect 3449 7588 3505 7590
rect 3529 7588 3585 7590
rect 5622 7098 5678 7100
rect 5702 7098 5758 7100
rect 5782 7098 5838 7100
rect 5862 7098 5918 7100
rect 5622 7046 5648 7098
rect 5648 7046 5678 7098
rect 5702 7046 5712 7098
rect 5712 7046 5758 7098
rect 5782 7046 5828 7098
rect 5828 7046 5838 7098
rect 5862 7046 5892 7098
rect 5892 7046 5918 7098
rect 5622 7044 5678 7046
rect 5702 7044 5758 7046
rect 5782 7044 5838 7046
rect 5862 7044 5918 7046
rect 3289 6554 3345 6556
rect 3369 6554 3425 6556
rect 3449 6554 3505 6556
rect 3529 6554 3585 6556
rect 3289 6502 3315 6554
rect 3315 6502 3345 6554
rect 3369 6502 3379 6554
rect 3379 6502 3425 6554
rect 3449 6502 3495 6554
rect 3495 6502 3505 6554
rect 3529 6502 3559 6554
rect 3559 6502 3585 6554
rect 3289 6500 3345 6502
rect 3369 6500 3425 6502
rect 3449 6500 3505 6502
rect 3529 6500 3585 6502
rect 5622 6010 5678 6012
rect 5702 6010 5758 6012
rect 5782 6010 5838 6012
rect 5862 6010 5918 6012
rect 5622 5958 5648 6010
rect 5648 5958 5678 6010
rect 5702 5958 5712 6010
rect 5712 5958 5758 6010
rect 5782 5958 5828 6010
rect 5828 5958 5838 6010
rect 5862 5958 5892 6010
rect 5892 5958 5918 6010
rect 5622 5956 5678 5958
rect 5702 5956 5758 5958
rect 5782 5956 5838 5958
rect 5862 5956 5918 5958
rect 3289 5466 3345 5468
rect 3369 5466 3425 5468
rect 3449 5466 3505 5468
rect 3529 5466 3585 5468
rect 3289 5414 3315 5466
rect 3315 5414 3345 5466
rect 3369 5414 3379 5466
rect 3379 5414 3425 5466
rect 3449 5414 3495 5466
rect 3495 5414 3505 5466
rect 3529 5414 3559 5466
rect 3559 5414 3585 5466
rect 3289 5412 3345 5414
rect 3369 5412 3425 5414
rect 3449 5412 3505 5414
rect 3529 5412 3585 5414
rect 5622 4922 5678 4924
rect 5702 4922 5758 4924
rect 5782 4922 5838 4924
rect 5862 4922 5918 4924
rect 5622 4870 5648 4922
rect 5648 4870 5678 4922
rect 5702 4870 5712 4922
rect 5712 4870 5758 4922
rect 5782 4870 5828 4922
rect 5828 4870 5838 4922
rect 5862 4870 5892 4922
rect 5892 4870 5918 4922
rect 5622 4868 5678 4870
rect 5702 4868 5758 4870
rect 5782 4868 5838 4870
rect 5862 4868 5918 4870
rect 3289 4378 3345 4380
rect 3369 4378 3425 4380
rect 3449 4378 3505 4380
rect 3529 4378 3585 4380
rect 3289 4326 3315 4378
rect 3315 4326 3345 4378
rect 3369 4326 3379 4378
rect 3379 4326 3425 4378
rect 3449 4326 3495 4378
rect 3495 4326 3505 4378
rect 3529 4326 3559 4378
rect 3559 4326 3585 4378
rect 3289 4324 3345 4326
rect 3369 4324 3425 4326
rect 3449 4324 3505 4326
rect 3529 4324 3585 4326
rect 5622 3834 5678 3836
rect 5702 3834 5758 3836
rect 5782 3834 5838 3836
rect 5862 3834 5918 3836
rect 5622 3782 5648 3834
rect 5648 3782 5678 3834
rect 5702 3782 5712 3834
rect 5712 3782 5758 3834
rect 5782 3782 5828 3834
rect 5828 3782 5838 3834
rect 5862 3782 5892 3834
rect 5892 3782 5918 3834
rect 5622 3780 5678 3782
rect 5702 3780 5758 3782
rect 5782 3780 5838 3782
rect 5862 3780 5918 3782
rect 3289 3290 3345 3292
rect 3369 3290 3425 3292
rect 3449 3290 3505 3292
rect 3529 3290 3585 3292
rect 3289 3238 3315 3290
rect 3315 3238 3345 3290
rect 3369 3238 3379 3290
rect 3379 3238 3425 3290
rect 3449 3238 3495 3290
rect 3495 3238 3505 3290
rect 3529 3238 3559 3290
rect 3559 3238 3585 3290
rect 3289 3236 3345 3238
rect 3369 3236 3425 3238
rect 3449 3236 3505 3238
rect 3529 3236 3585 3238
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 7982 13082
rect 7982 13030 8012 13082
rect 8036 13030 8046 13082
rect 8046 13030 8092 13082
rect 8116 13030 8162 13082
rect 8162 13030 8172 13082
rect 8196 13030 8226 13082
rect 8226 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 11518 85196 11574 85232
rect 11518 85176 11520 85196
rect 11520 85176 11572 85196
rect 11572 85176 11574 85196
rect 11150 85040 11206 85096
rect 11242 71576 11298 71632
rect 11426 71440 11482 71496
rect 11426 64640 11482 64696
rect 11242 58520 11298 58576
rect 11426 57840 11482 57896
rect 11518 44784 11574 44840
rect 11426 37440 11482 37496
rect 11702 51040 11758 51096
rect 11242 17176 11298 17232
rect 11150 17040 11206 17096
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 7982 11994
rect 7982 11942 8012 11994
rect 8036 11942 8046 11994
rect 8046 11942 8092 11994
rect 8116 11942 8162 11994
rect 8162 11942 8172 11994
rect 8196 11942 8226 11994
rect 8226 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 7982 10906
rect 7982 10854 8012 10906
rect 8036 10854 8046 10906
rect 8046 10854 8092 10906
rect 8116 10854 8162 10906
rect 8162 10854 8172 10906
rect 8196 10854 8226 10906
rect 8226 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 7982 9818
rect 7982 9766 8012 9818
rect 8036 9766 8046 9818
rect 8046 9766 8092 9818
rect 8116 9766 8162 9818
rect 8162 9766 8172 9818
rect 8196 9766 8226 9818
rect 8226 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 7982 8730
rect 7982 8678 8012 8730
rect 8036 8678 8046 8730
rect 8046 8678 8092 8730
rect 8116 8678 8162 8730
rect 8162 8678 8172 8730
rect 8196 8678 8226 8730
rect 8226 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 7982 7642
rect 7982 7590 8012 7642
rect 8036 7590 8046 7642
rect 8046 7590 8092 7642
rect 8116 7590 8162 7642
rect 8162 7590 8172 7642
rect 8196 7590 8226 7642
rect 8226 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 7982 6554
rect 7982 6502 8012 6554
rect 8036 6502 8046 6554
rect 8046 6502 8092 6554
rect 8116 6502 8162 6554
rect 8162 6502 8172 6554
rect 8196 6502 8226 6554
rect 8226 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 7982 5466
rect 7982 5414 8012 5466
rect 8036 5414 8046 5466
rect 8046 5414 8092 5466
rect 8116 5414 8162 5466
rect 8162 5414 8172 5466
rect 8196 5414 8226 5466
rect 8226 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 7982 4378
rect 7982 4326 8012 4378
rect 8036 4326 8046 4378
rect 8046 4326 8092 4378
rect 8116 4326 8162 4378
rect 8162 4326 8172 4378
rect 8196 4326 8226 4378
rect 8226 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 7982 3290
rect 7982 3238 8012 3290
rect 8036 3238 8046 3290
rect 8046 3238 8092 3290
rect 8116 3238 8162 3290
rect 8162 3238 8172 3290
rect 8196 3238 8226 3290
rect 8226 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 11426 10240 11482 10296
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11242 5616 11298 5672
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 5622 2746 5678 2748
rect 5702 2746 5758 2748
rect 5782 2746 5838 2748
rect 5862 2746 5918 2748
rect 5622 2694 5648 2746
rect 5648 2694 5678 2746
rect 5702 2694 5712 2746
rect 5712 2694 5758 2746
rect 5782 2694 5828 2746
rect 5828 2694 5838 2746
rect 5862 2694 5892 2746
rect 5892 2694 5918 2746
rect 5622 2692 5678 2694
rect 5702 2692 5758 2694
rect 5782 2692 5838 2694
rect 5862 2692 5918 2694
rect 3289 2202 3345 2204
rect 3369 2202 3425 2204
rect 3449 2202 3505 2204
rect 3529 2202 3585 2204
rect 3289 2150 3315 2202
rect 3315 2150 3345 2202
rect 3369 2150 3379 2202
rect 3379 2150 3425 2202
rect 3449 2150 3495 2202
rect 3495 2150 3505 2202
rect 3529 2150 3559 2202
rect 3559 2150 3585 2202
rect 3289 2148 3345 2150
rect 3369 2148 3425 2150
rect 3449 2148 3505 2150
rect 3529 2148 3585 2150
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 7982 2202
rect 7982 2150 8012 2202
rect 8036 2150 8046 2202
rect 8046 2150 8092 2202
rect 8116 2150 8162 2202
rect 8162 2150 8172 2202
rect 8196 2150 8226 2202
rect 8226 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10966 3440 11022 3496
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
<< metal3 >>
rect 3277 106656 3597 106657
rect 3277 106592 3285 106656
rect 3349 106592 3365 106656
rect 3429 106592 3445 106656
rect 3509 106592 3525 106656
rect 3589 106592 3597 106656
rect 3277 106591 3597 106592
rect 7944 106656 8264 106657
rect 7944 106592 7952 106656
rect 8016 106592 8032 106656
rect 8096 106592 8112 106656
rect 8176 106592 8192 106656
rect 8256 106592 8264 106656
rect 7944 106591 8264 106592
rect 5610 106112 5930 106113
rect 5610 106048 5618 106112
rect 5682 106048 5698 106112
rect 5762 106048 5778 106112
rect 5842 106048 5858 106112
rect 5922 106048 5930 106112
rect 5610 106047 5930 106048
rect 10277 106112 10597 106113
rect 10277 106048 10285 106112
rect 10349 106048 10365 106112
rect 10429 106048 10445 106112
rect 10509 106048 10525 106112
rect 10589 106048 10597 106112
rect 10277 106047 10597 106048
rect 3277 105568 3597 105569
rect 3277 105504 3285 105568
rect 3349 105504 3365 105568
rect 3429 105504 3445 105568
rect 3509 105504 3525 105568
rect 3589 105504 3597 105568
rect 3277 105503 3597 105504
rect 7944 105568 8264 105569
rect 7944 105504 7952 105568
rect 8016 105504 8032 105568
rect 8096 105504 8112 105568
rect 8176 105504 8192 105568
rect 8256 105504 8264 105568
rect 7944 105503 8264 105504
rect 11421 105498 11487 105501
rect 13520 105498 14000 105528
rect 11421 105496 14000 105498
rect 11421 105440 11426 105496
rect 11482 105440 14000 105496
rect 11421 105438 14000 105440
rect 11421 105435 11487 105438
rect 13520 105408 14000 105438
rect 5610 105024 5930 105025
rect 5610 104960 5618 105024
rect 5682 104960 5698 105024
rect 5762 104960 5778 105024
rect 5842 104960 5858 105024
rect 5922 104960 5930 105024
rect 5610 104959 5930 104960
rect 10277 105024 10597 105025
rect 10277 104960 10285 105024
rect 10349 104960 10365 105024
rect 10429 104960 10445 105024
rect 10509 104960 10525 105024
rect 10589 104960 10597 105024
rect 10277 104959 10597 104960
rect 3277 104480 3597 104481
rect 3277 104416 3285 104480
rect 3349 104416 3365 104480
rect 3429 104416 3445 104480
rect 3509 104416 3525 104480
rect 3589 104416 3597 104480
rect 3277 104415 3597 104416
rect 7944 104480 8264 104481
rect 7944 104416 7952 104480
rect 8016 104416 8032 104480
rect 8096 104416 8112 104480
rect 8176 104416 8192 104480
rect 8256 104416 8264 104480
rect 7944 104415 8264 104416
rect 5610 103936 5930 103937
rect 5610 103872 5618 103936
rect 5682 103872 5698 103936
rect 5762 103872 5778 103936
rect 5842 103872 5858 103936
rect 5922 103872 5930 103936
rect 5610 103871 5930 103872
rect 10277 103936 10597 103937
rect 10277 103872 10285 103936
rect 10349 103872 10365 103936
rect 10429 103872 10445 103936
rect 10509 103872 10525 103936
rect 10589 103872 10597 103936
rect 10277 103871 10597 103872
rect 3277 103392 3597 103393
rect 3277 103328 3285 103392
rect 3349 103328 3365 103392
rect 3429 103328 3445 103392
rect 3509 103328 3525 103392
rect 3589 103328 3597 103392
rect 3277 103327 3597 103328
rect 7944 103392 8264 103393
rect 7944 103328 7952 103392
rect 8016 103328 8032 103392
rect 8096 103328 8112 103392
rect 8176 103328 8192 103392
rect 8256 103328 8264 103392
rect 7944 103327 8264 103328
rect 5610 102848 5930 102849
rect 5610 102784 5618 102848
rect 5682 102784 5698 102848
rect 5762 102784 5778 102848
rect 5842 102784 5858 102848
rect 5922 102784 5930 102848
rect 5610 102783 5930 102784
rect 10277 102848 10597 102849
rect 10277 102784 10285 102848
rect 10349 102784 10365 102848
rect 10429 102784 10445 102848
rect 10509 102784 10525 102848
rect 10589 102784 10597 102848
rect 10277 102783 10597 102784
rect 3277 102304 3597 102305
rect 3277 102240 3285 102304
rect 3349 102240 3365 102304
rect 3429 102240 3445 102304
rect 3509 102240 3525 102304
rect 3589 102240 3597 102304
rect 3277 102239 3597 102240
rect 7944 102304 8264 102305
rect 7944 102240 7952 102304
rect 8016 102240 8032 102304
rect 8096 102240 8112 102304
rect 8176 102240 8192 102304
rect 8256 102240 8264 102304
rect 7944 102239 8264 102240
rect 0 102096 480 102128
rect 0 102040 110 102096
rect 166 102040 480 102096
rect 0 102008 480 102040
rect 5610 101760 5930 101761
rect 5610 101696 5618 101760
rect 5682 101696 5698 101760
rect 5762 101696 5778 101760
rect 5842 101696 5858 101760
rect 5922 101696 5930 101760
rect 5610 101695 5930 101696
rect 10277 101760 10597 101761
rect 10277 101696 10285 101760
rect 10349 101696 10365 101760
rect 10429 101696 10445 101760
rect 10509 101696 10525 101760
rect 10589 101696 10597 101760
rect 10277 101695 10597 101696
rect 3277 101216 3597 101217
rect 3277 101152 3285 101216
rect 3349 101152 3365 101216
rect 3429 101152 3445 101216
rect 3509 101152 3525 101216
rect 3589 101152 3597 101216
rect 3277 101151 3597 101152
rect 7944 101216 8264 101217
rect 7944 101152 7952 101216
rect 8016 101152 8032 101216
rect 8096 101152 8112 101216
rect 8176 101152 8192 101216
rect 8256 101152 8264 101216
rect 7944 101151 8264 101152
rect 5610 100672 5930 100673
rect 5610 100608 5618 100672
rect 5682 100608 5698 100672
rect 5762 100608 5778 100672
rect 5842 100608 5858 100672
rect 5922 100608 5930 100672
rect 5610 100607 5930 100608
rect 10277 100672 10597 100673
rect 10277 100608 10285 100672
rect 10349 100608 10365 100672
rect 10429 100608 10445 100672
rect 10509 100608 10525 100672
rect 10589 100608 10597 100672
rect 10277 100607 10597 100608
rect 3277 100128 3597 100129
rect 3277 100064 3285 100128
rect 3349 100064 3365 100128
rect 3429 100064 3445 100128
rect 3509 100064 3525 100128
rect 3589 100064 3597 100128
rect 3277 100063 3597 100064
rect 7944 100128 8264 100129
rect 7944 100064 7952 100128
rect 8016 100064 8032 100128
rect 8096 100064 8112 100128
rect 8176 100064 8192 100128
rect 8256 100064 8264 100128
rect 7944 100063 8264 100064
rect 5610 99584 5930 99585
rect 5610 99520 5618 99584
rect 5682 99520 5698 99584
rect 5762 99520 5778 99584
rect 5842 99520 5858 99584
rect 5922 99520 5930 99584
rect 5610 99519 5930 99520
rect 10277 99584 10597 99585
rect 10277 99520 10285 99584
rect 10349 99520 10365 99584
rect 10429 99520 10445 99584
rect 10509 99520 10525 99584
rect 10589 99520 10597 99584
rect 10277 99519 10597 99520
rect 3277 99040 3597 99041
rect 3277 98976 3285 99040
rect 3349 98976 3365 99040
rect 3429 98976 3445 99040
rect 3509 98976 3525 99040
rect 3589 98976 3597 99040
rect 3277 98975 3597 98976
rect 7944 99040 8264 99041
rect 7944 98976 7952 99040
rect 8016 98976 8032 99040
rect 8096 98976 8112 99040
rect 8176 98976 8192 99040
rect 8256 98976 8264 99040
rect 7944 98975 8264 98976
rect 11145 98698 11211 98701
rect 13520 98698 14000 98728
rect 11145 98696 14000 98698
rect 11145 98640 11150 98696
rect 11206 98640 14000 98696
rect 11145 98638 14000 98640
rect 11145 98635 11211 98638
rect 13520 98608 14000 98638
rect 5610 98496 5930 98497
rect 5610 98432 5618 98496
rect 5682 98432 5698 98496
rect 5762 98432 5778 98496
rect 5842 98432 5858 98496
rect 5922 98432 5930 98496
rect 5610 98431 5930 98432
rect 10277 98496 10597 98497
rect 10277 98432 10285 98496
rect 10349 98432 10365 98496
rect 10429 98432 10445 98496
rect 10509 98432 10525 98496
rect 10589 98432 10597 98496
rect 10277 98431 10597 98432
rect 3277 97952 3597 97953
rect 3277 97888 3285 97952
rect 3349 97888 3365 97952
rect 3429 97888 3445 97952
rect 3509 97888 3525 97952
rect 3589 97888 3597 97952
rect 3277 97887 3597 97888
rect 7944 97952 8264 97953
rect 7944 97888 7952 97952
rect 8016 97888 8032 97952
rect 8096 97888 8112 97952
rect 8176 97888 8192 97952
rect 8256 97888 8264 97952
rect 7944 97887 8264 97888
rect 5610 97408 5930 97409
rect 5610 97344 5618 97408
rect 5682 97344 5698 97408
rect 5762 97344 5778 97408
rect 5842 97344 5858 97408
rect 5922 97344 5930 97408
rect 5610 97343 5930 97344
rect 10277 97408 10597 97409
rect 10277 97344 10285 97408
rect 10349 97344 10365 97408
rect 10429 97344 10445 97408
rect 10509 97344 10525 97408
rect 10589 97344 10597 97408
rect 10277 97343 10597 97344
rect 105 97202 171 97205
rect 11237 97202 11303 97205
rect 105 97200 11303 97202
rect 105 97144 110 97200
rect 166 97144 11242 97200
rect 11298 97144 11303 97200
rect 105 97142 11303 97144
rect 105 97139 171 97142
rect 11237 97139 11303 97142
rect 3277 96864 3597 96865
rect 3277 96800 3285 96864
rect 3349 96800 3365 96864
rect 3429 96800 3445 96864
rect 3509 96800 3525 96864
rect 3589 96800 3597 96864
rect 3277 96799 3597 96800
rect 7944 96864 8264 96865
rect 7944 96800 7952 96864
rect 8016 96800 8032 96864
rect 8096 96800 8112 96864
rect 8176 96800 8192 96864
rect 8256 96800 8264 96864
rect 7944 96799 8264 96800
rect 5610 96320 5930 96321
rect 5610 96256 5618 96320
rect 5682 96256 5698 96320
rect 5762 96256 5778 96320
rect 5842 96256 5858 96320
rect 5922 96256 5930 96320
rect 5610 96255 5930 96256
rect 10277 96320 10597 96321
rect 10277 96256 10285 96320
rect 10349 96256 10365 96320
rect 10429 96256 10445 96320
rect 10509 96256 10525 96320
rect 10589 96256 10597 96320
rect 10277 96255 10597 96256
rect 3277 95776 3597 95777
rect 3277 95712 3285 95776
rect 3349 95712 3365 95776
rect 3429 95712 3445 95776
rect 3509 95712 3525 95776
rect 3589 95712 3597 95776
rect 3277 95711 3597 95712
rect 7944 95776 8264 95777
rect 7944 95712 7952 95776
rect 8016 95712 8032 95776
rect 8096 95712 8112 95776
rect 8176 95712 8192 95776
rect 8256 95712 8264 95776
rect 7944 95711 8264 95712
rect 5610 95232 5930 95233
rect 5610 95168 5618 95232
rect 5682 95168 5698 95232
rect 5762 95168 5778 95232
rect 5842 95168 5858 95232
rect 5922 95168 5930 95232
rect 5610 95167 5930 95168
rect 10277 95232 10597 95233
rect 10277 95168 10285 95232
rect 10349 95168 10365 95232
rect 10429 95168 10445 95232
rect 10509 95168 10525 95232
rect 10589 95168 10597 95232
rect 10277 95167 10597 95168
rect 3277 94688 3597 94689
rect 3277 94624 3285 94688
rect 3349 94624 3365 94688
rect 3429 94624 3445 94688
rect 3509 94624 3525 94688
rect 3589 94624 3597 94688
rect 3277 94623 3597 94624
rect 7944 94688 8264 94689
rect 7944 94624 7952 94688
rect 8016 94624 8032 94688
rect 8096 94624 8112 94688
rect 8176 94624 8192 94688
rect 8256 94624 8264 94688
rect 7944 94623 8264 94624
rect 5610 94144 5930 94145
rect 5610 94080 5618 94144
rect 5682 94080 5698 94144
rect 5762 94080 5778 94144
rect 5842 94080 5858 94144
rect 5922 94080 5930 94144
rect 5610 94079 5930 94080
rect 10277 94144 10597 94145
rect 10277 94080 10285 94144
rect 10349 94080 10365 94144
rect 10429 94080 10445 94144
rect 10509 94080 10525 94144
rect 10589 94080 10597 94144
rect 10277 94079 10597 94080
rect 3277 93600 3597 93601
rect 3277 93536 3285 93600
rect 3349 93536 3365 93600
rect 3429 93536 3445 93600
rect 3509 93536 3525 93600
rect 3589 93536 3597 93600
rect 3277 93535 3597 93536
rect 7944 93600 8264 93601
rect 7944 93536 7952 93600
rect 8016 93536 8032 93600
rect 8096 93536 8112 93600
rect 8176 93536 8192 93600
rect 8256 93536 8264 93600
rect 7944 93535 8264 93536
rect 5610 93056 5930 93057
rect 5610 92992 5618 93056
rect 5682 92992 5698 93056
rect 5762 92992 5778 93056
rect 5842 92992 5858 93056
rect 5922 92992 5930 93056
rect 5610 92991 5930 92992
rect 10277 93056 10597 93057
rect 10277 92992 10285 93056
rect 10349 92992 10365 93056
rect 10429 92992 10445 93056
rect 10509 92992 10525 93056
rect 10589 92992 10597 93056
rect 10277 92991 10597 92992
rect 3277 92512 3597 92513
rect 3277 92448 3285 92512
rect 3349 92448 3365 92512
rect 3429 92448 3445 92512
rect 3509 92448 3525 92512
rect 3589 92448 3597 92512
rect 3277 92447 3597 92448
rect 7944 92512 8264 92513
rect 7944 92448 7952 92512
rect 8016 92448 8032 92512
rect 8096 92448 8112 92512
rect 8176 92448 8192 92512
rect 8256 92448 8264 92512
rect 7944 92447 8264 92448
rect 5610 91968 5930 91969
rect 5610 91904 5618 91968
rect 5682 91904 5698 91968
rect 5762 91904 5778 91968
rect 5842 91904 5858 91968
rect 5922 91904 5930 91968
rect 5610 91903 5930 91904
rect 10277 91968 10597 91969
rect 10277 91904 10285 91968
rect 10349 91904 10365 91968
rect 10429 91904 10445 91968
rect 10509 91904 10525 91968
rect 10589 91904 10597 91968
rect 10277 91903 10597 91904
rect 10685 91898 10751 91901
rect 13520 91898 14000 91928
rect 10685 91896 14000 91898
rect 10685 91840 10690 91896
rect 10746 91840 14000 91896
rect 10685 91838 14000 91840
rect 10685 91835 10751 91838
rect 13520 91808 14000 91838
rect 3277 91424 3597 91425
rect 3277 91360 3285 91424
rect 3349 91360 3365 91424
rect 3429 91360 3445 91424
rect 3509 91360 3525 91424
rect 3589 91360 3597 91424
rect 3277 91359 3597 91360
rect 7944 91424 8264 91425
rect 7944 91360 7952 91424
rect 8016 91360 8032 91424
rect 8096 91360 8112 91424
rect 8176 91360 8192 91424
rect 8256 91360 8264 91424
rect 7944 91359 8264 91360
rect 5610 90880 5930 90881
rect 5610 90816 5618 90880
rect 5682 90816 5698 90880
rect 5762 90816 5778 90880
rect 5842 90816 5858 90880
rect 5922 90816 5930 90880
rect 5610 90815 5930 90816
rect 10277 90880 10597 90881
rect 10277 90816 10285 90880
rect 10349 90816 10365 90880
rect 10429 90816 10445 90880
rect 10509 90816 10525 90880
rect 10589 90816 10597 90880
rect 10277 90815 10597 90816
rect 3277 90336 3597 90337
rect 3277 90272 3285 90336
rect 3349 90272 3365 90336
rect 3429 90272 3445 90336
rect 3509 90272 3525 90336
rect 3589 90272 3597 90336
rect 3277 90271 3597 90272
rect 7944 90336 8264 90337
rect 7944 90272 7952 90336
rect 8016 90272 8032 90336
rect 8096 90272 8112 90336
rect 8176 90272 8192 90336
rect 8256 90272 8264 90336
rect 7944 90271 8264 90272
rect 5610 89792 5930 89793
rect 5610 89728 5618 89792
rect 5682 89728 5698 89792
rect 5762 89728 5778 89792
rect 5842 89728 5858 89792
rect 5922 89728 5930 89792
rect 5610 89727 5930 89728
rect 10277 89792 10597 89793
rect 10277 89728 10285 89792
rect 10349 89728 10365 89792
rect 10429 89728 10445 89792
rect 10509 89728 10525 89792
rect 10589 89728 10597 89792
rect 10277 89727 10597 89728
rect 3277 89248 3597 89249
rect 3277 89184 3285 89248
rect 3349 89184 3365 89248
rect 3429 89184 3445 89248
rect 3509 89184 3525 89248
rect 3589 89184 3597 89248
rect 3277 89183 3597 89184
rect 7944 89248 8264 89249
rect 7944 89184 7952 89248
rect 8016 89184 8032 89248
rect 8096 89184 8112 89248
rect 8176 89184 8192 89248
rect 8256 89184 8264 89248
rect 7944 89183 8264 89184
rect 5610 88704 5930 88705
rect 5610 88640 5618 88704
rect 5682 88640 5698 88704
rect 5762 88640 5778 88704
rect 5842 88640 5858 88704
rect 5922 88640 5930 88704
rect 5610 88639 5930 88640
rect 10277 88704 10597 88705
rect 10277 88640 10285 88704
rect 10349 88640 10365 88704
rect 10429 88640 10445 88704
rect 10509 88640 10525 88704
rect 10589 88640 10597 88704
rect 10277 88639 10597 88640
rect 0 88496 480 88528
rect 0 88440 110 88496
rect 166 88440 480 88496
rect 0 88408 480 88440
rect 3277 88160 3597 88161
rect 3277 88096 3285 88160
rect 3349 88096 3365 88160
rect 3429 88096 3445 88160
rect 3509 88096 3525 88160
rect 3589 88096 3597 88160
rect 3277 88095 3597 88096
rect 7944 88160 8264 88161
rect 7944 88096 7952 88160
rect 8016 88096 8032 88160
rect 8096 88096 8112 88160
rect 8176 88096 8192 88160
rect 8256 88096 8264 88160
rect 7944 88095 8264 88096
rect 5610 87616 5930 87617
rect 5610 87552 5618 87616
rect 5682 87552 5698 87616
rect 5762 87552 5778 87616
rect 5842 87552 5858 87616
rect 5922 87552 5930 87616
rect 5610 87551 5930 87552
rect 10277 87616 10597 87617
rect 10277 87552 10285 87616
rect 10349 87552 10365 87616
rect 10429 87552 10445 87616
rect 10509 87552 10525 87616
rect 10589 87552 10597 87616
rect 10277 87551 10597 87552
rect 3277 87072 3597 87073
rect 3277 87008 3285 87072
rect 3349 87008 3365 87072
rect 3429 87008 3445 87072
rect 3509 87008 3525 87072
rect 3589 87008 3597 87072
rect 3277 87007 3597 87008
rect 7944 87072 8264 87073
rect 7944 87008 7952 87072
rect 8016 87008 8032 87072
rect 8096 87008 8112 87072
rect 8176 87008 8192 87072
rect 8256 87008 8264 87072
rect 7944 87007 8264 87008
rect 5610 86528 5930 86529
rect 5610 86464 5618 86528
rect 5682 86464 5698 86528
rect 5762 86464 5778 86528
rect 5842 86464 5858 86528
rect 5922 86464 5930 86528
rect 5610 86463 5930 86464
rect 10277 86528 10597 86529
rect 10277 86464 10285 86528
rect 10349 86464 10365 86528
rect 10429 86464 10445 86528
rect 10509 86464 10525 86528
rect 10589 86464 10597 86528
rect 10277 86463 10597 86464
rect 3277 85984 3597 85985
rect 3277 85920 3285 85984
rect 3349 85920 3365 85984
rect 3429 85920 3445 85984
rect 3509 85920 3525 85984
rect 3589 85920 3597 85984
rect 3277 85919 3597 85920
rect 7944 85984 8264 85985
rect 7944 85920 7952 85984
rect 8016 85920 8032 85984
rect 8096 85920 8112 85984
rect 8176 85920 8192 85984
rect 8256 85920 8264 85984
rect 7944 85919 8264 85920
rect 5610 85440 5930 85441
rect 5610 85376 5618 85440
rect 5682 85376 5698 85440
rect 5762 85376 5778 85440
rect 5842 85376 5858 85440
rect 5922 85376 5930 85440
rect 5610 85375 5930 85376
rect 10277 85440 10597 85441
rect 10277 85376 10285 85440
rect 10349 85376 10365 85440
rect 10429 85376 10445 85440
rect 10509 85376 10525 85440
rect 10589 85376 10597 85440
rect 10277 85375 10597 85376
rect 105 85234 171 85237
rect 11513 85234 11579 85237
rect 105 85232 11579 85234
rect 105 85176 110 85232
rect 166 85176 11518 85232
rect 11574 85176 11579 85232
rect 105 85174 11579 85176
rect 105 85171 171 85174
rect 11513 85171 11579 85174
rect 11145 85098 11211 85101
rect 13520 85098 14000 85128
rect 11145 85096 14000 85098
rect 11145 85040 11150 85096
rect 11206 85040 14000 85096
rect 11145 85038 14000 85040
rect 11145 85035 11211 85038
rect 13520 85008 14000 85038
rect 3277 84896 3597 84897
rect 3277 84832 3285 84896
rect 3349 84832 3365 84896
rect 3429 84832 3445 84896
rect 3509 84832 3525 84896
rect 3589 84832 3597 84896
rect 3277 84831 3597 84832
rect 7944 84896 8264 84897
rect 7944 84832 7952 84896
rect 8016 84832 8032 84896
rect 8096 84832 8112 84896
rect 8176 84832 8192 84896
rect 8256 84832 8264 84896
rect 7944 84831 8264 84832
rect 5610 84352 5930 84353
rect 5610 84288 5618 84352
rect 5682 84288 5698 84352
rect 5762 84288 5778 84352
rect 5842 84288 5858 84352
rect 5922 84288 5930 84352
rect 5610 84287 5930 84288
rect 10277 84352 10597 84353
rect 10277 84288 10285 84352
rect 10349 84288 10365 84352
rect 10429 84288 10445 84352
rect 10509 84288 10525 84352
rect 10589 84288 10597 84352
rect 10277 84287 10597 84288
rect 3277 83808 3597 83809
rect 3277 83744 3285 83808
rect 3349 83744 3365 83808
rect 3429 83744 3445 83808
rect 3509 83744 3525 83808
rect 3589 83744 3597 83808
rect 3277 83743 3597 83744
rect 7944 83808 8264 83809
rect 7944 83744 7952 83808
rect 8016 83744 8032 83808
rect 8096 83744 8112 83808
rect 8176 83744 8192 83808
rect 8256 83744 8264 83808
rect 7944 83743 8264 83744
rect 5610 83264 5930 83265
rect 5610 83200 5618 83264
rect 5682 83200 5698 83264
rect 5762 83200 5778 83264
rect 5842 83200 5858 83264
rect 5922 83200 5930 83264
rect 5610 83199 5930 83200
rect 10277 83264 10597 83265
rect 10277 83200 10285 83264
rect 10349 83200 10365 83264
rect 10429 83200 10445 83264
rect 10509 83200 10525 83264
rect 10589 83200 10597 83264
rect 10277 83199 10597 83200
rect 3277 82720 3597 82721
rect 3277 82656 3285 82720
rect 3349 82656 3365 82720
rect 3429 82656 3445 82720
rect 3509 82656 3525 82720
rect 3589 82656 3597 82720
rect 3277 82655 3597 82656
rect 7944 82720 8264 82721
rect 7944 82656 7952 82720
rect 8016 82656 8032 82720
rect 8096 82656 8112 82720
rect 8176 82656 8192 82720
rect 8256 82656 8264 82720
rect 7944 82655 8264 82656
rect 5610 82176 5930 82177
rect 5610 82112 5618 82176
rect 5682 82112 5698 82176
rect 5762 82112 5778 82176
rect 5842 82112 5858 82176
rect 5922 82112 5930 82176
rect 5610 82111 5930 82112
rect 10277 82176 10597 82177
rect 10277 82112 10285 82176
rect 10349 82112 10365 82176
rect 10429 82112 10445 82176
rect 10509 82112 10525 82176
rect 10589 82112 10597 82176
rect 10277 82111 10597 82112
rect 3277 81632 3597 81633
rect 3277 81568 3285 81632
rect 3349 81568 3365 81632
rect 3429 81568 3445 81632
rect 3509 81568 3525 81632
rect 3589 81568 3597 81632
rect 3277 81567 3597 81568
rect 7944 81632 8264 81633
rect 7944 81568 7952 81632
rect 8016 81568 8032 81632
rect 8096 81568 8112 81632
rect 8176 81568 8192 81632
rect 8256 81568 8264 81632
rect 7944 81567 8264 81568
rect 5610 81088 5930 81089
rect 5610 81024 5618 81088
rect 5682 81024 5698 81088
rect 5762 81024 5778 81088
rect 5842 81024 5858 81088
rect 5922 81024 5930 81088
rect 5610 81023 5930 81024
rect 10277 81088 10597 81089
rect 10277 81024 10285 81088
rect 10349 81024 10365 81088
rect 10429 81024 10445 81088
rect 10509 81024 10525 81088
rect 10589 81024 10597 81088
rect 10277 81023 10597 81024
rect 3277 80544 3597 80545
rect 3277 80480 3285 80544
rect 3349 80480 3365 80544
rect 3429 80480 3445 80544
rect 3509 80480 3525 80544
rect 3589 80480 3597 80544
rect 3277 80479 3597 80480
rect 7944 80544 8264 80545
rect 7944 80480 7952 80544
rect 8016 80480 8032 80544
rect 8096 80480 8112 80544
rect 8176 80480 8192 80544
rect 8256 80480 8264 80544
rect 7944 80479 8264 80480
rect 5610 80000 5930 80001
rect 5610 79936 5618 80000
rect 5682 79936 5698 80000
rect 5762 79936 5778 80000
rect 5842 79936 5858 80000
rect 5922 79936 5930 80000
rect 5610 79935 5930 79936
rect 10277 80000 10597 80001
rect 10277 79936 10285 80000
rect 10349 79936 10365 80000
rect 10429 79936 10445 80000
rect 10509 79936 10525 80000
rect 10589 79936 10597 80000
rect 10277 79935 10597 79936
rect 3277 79456 3597 79457
rect 3277 79392 3285 79456
rect 3349 79392 3365 79456
rect 3429 79392 3445 79456
rect 3509 79392 3525 79456
rect 3589 79392 3597 79456
rect 3277 79391 3597 79392
rect 7944 79456 8264 79457
rect 7944 79392 7952 79456
rect 8016 79392 8032 79456
rect 8096 79392 8112 79456
rect 8176 79392 8192 79456
rect 8256 79392 8264 79456
rect 7944 79391 8264 79392
rect 5610 78912 5930 78913
rect 5610 78848 5618 78912
rect 5682 78848 5698 78912
rect 5762 78848 5778 78912
rect 5842 78848 5858 78912
rect 5922 78848 5930 78912
rect 5610 78847 5930 78848
rect 10277 78912 10597 78913
rect 10277 78848 10285 78912
rect 10349 78848 10365 78912
rect 10429 78848 10445 78912
rect 10509 78848 10525 78912
rect 10589 78848 10597 78912
rect 10277 78847 10597 78848
rect 3277 78368 3597 78369
rect 3277 78304 3285 78368
rect 3349 78304 3365 78368
rect 3429 78304 3445 78368
rect 3509 78304 3525 78368
rect 3589 78304 3597 78368
rect 3277 78303 3597 78304
rect 7944 78368 8264 78369
rect 7944 78304 7952 78368
rect 8016 78304 8032 78368
rect 8096 78304 8112 78368
rect 8176 78304 8192 78368
rect 8256 78304 8264 78368
rect 7944 78303 8264 78304
rect 10961 78298 11027 78301
rect 13520 78298 14000 78328
rect 10961 78296 14000 78298
rect 10961 78240 10966 78296
rect 11022 78240 14000 78296
rect 10961 78238 14000 78240
rect 10961 78235 11027 78238
rect 13520 78208 14000 78238
rect 5610 77824 5930 77825
rect 5610 77760 5618 77824
rect 5682 77760 5698 77824
rect 5762 77760 5778 77824
rect 5842 77760 5858 77824
rect 5922 77760 5930 77824
rect 5610 77759 5930 77760
rect 10277 77824 10597 77825
rect 10277 77760 10285 77824
rect 10349 77760 10365 77824
rect 10429 77760 10445 77824
rect 10509 77760 10525 77824
rect 10589 77760 10597 77824
rect 10277 77759 10597 77760
rect 3277 77280 3597 77281
rect 3277 77216 3285 77280
rect 3349 77216 3365 77280
rect 3429 77216 3445 77280
rect 3509 77216 3525 77280
rect 3589 77216 3597 77280
rect 3277 77215 3597 77216
rect 7944 77280 8264 77281
rect 7944 77216 7952 77280
rect 8016 77216 8032 77280
rect 8096 77216 8112 77280
rect 8176 77216 8192 77280
rect 8256 77216 8264 77280
rect 7944 77215 8264 77216
rect 5610 76736 5930 76737
rect 5610 76672 5618 76736
rect 5682 76672 5698 76736
rect 5762 76672 5778 76736
rect 5842 76672 5858 76736
rect 5922 76672 5930 76736
rect 5610 76671 5930 76672
rect 10277 76736 10597 76737
rect 10277 76672 10285 76736
rect 10349 76672 10365 76736
rect 10429 76672 10445 76736
rect 10509 76672 10525 76736
rect 10589 76672 10597 76736
rect 10277 76671 10597 76672
rect 3277 76192 3597 76193
rect 3277 76128 3285 76192
rect 3349 76128 3365 76192
rect 3429 76128 3445 76192
rect 3509 76128 3525 76192
rect 3589 76128 3597 76192
rect 3277 76127 3597 76128
rect 7944 76192 8264 76193
rect 7944 76128 7952 76192
rect 8016 76128 8032 76192
rect 8096 76128 8112 76192
rect 8176 76128 8192 76192
rect 8256 76128 8264 76192
rect 7944 76127 8264 76128
rect 5610 75648 5930 75649
rect 5610 75584 5618 75648
rect 5682 75584 5698 75648
rect 5762 75584 5778 75648
rect 5842 75584 5858 75648
rect 5922 75584 5930 75648
rect 5610 75583 5930 75584
rect 10277 75648 10597 75649
rect 10277 75584 10285 75648
rect 10349 75584 10365 75648
rect 10429 75584 10445 75648
rect 10509 75584 10525 75648
rect 10589 75584 10597 75648
rect 10277 75583 10597 75584
rect 3277 75104 3597 75105
rect 3277 75040 3285 75104
rect 3349 75040 3365 75104
rect 3429 75040 3445 75104
rect 3509 75040 3525 75104
rect 3589 75040 3597 75104
rect 3277 75039 3597 75040
rect 7944 75104 8264 75105
rect 7944 75040 7952 75104
rect 8016 75040 8032 75104
rect 8096 75040 8112 75104
rect 8176 75040 8192 75104
rect 8256 75040 8264 75104
rect 7944 75039 8264 75040
rect 0 74896 480 74928
rect 0 74840 110 74896
rect 166 74840 480 74896
rect 0 74808 480 74840
rect 5610 74560 5930 74561
rect 5610 74496 5618 74560
rect 5682 74496 5698 74560
rect 5762 74496 5778 74560
rect 5842 74496 5858 74560
rect 5922 74496 5930 74560
rect 5610 74495 5930 74496
rect 10277 74560 10597 74561
rect 10277 74496 10285 74560
rect 10349 74496 10365 74560
rect 10429 74496 10445 74560
rect 10509 74496 10525 74560
rect 10589 74496 10597 74560
rect 10277 74495 10597 74496
rect 3277 74016 3597 74017
rect 3277 73952 3285 74016
rect 3349 73952 3365 74016
rect 3429 73952 3445 74016
rect 3509 73952 3525 74016
rect 3589 73952 3597 74016
rect 3277 73951 3597 73952
rect 7944 74016 8264 74017
rect 7944 73952 7952 74016
rect 8016 73952 8032 74016
rect 8096 73952 8112 74016
rect 8176 73952 8192 74016
rect 8256 73952 8264 74016
rect 7944 73951 8264 73952
rect 5610 73472 5930 73473
rect 5610 73408 5618 73472
rect 5682 73408 5698 73472
rect 5762 73408 5778 73472
rect 5842 73408 5858 73472
rect 5922 73408 5930 73472
rect 5610 73407 5930 73408
rect 10277 73472 10597 73473
rect 10277 73408 10285 73472
rect 10349 73408 10365 73472
rect 10429 73408 10445 73472
rect 10509 73408 10525 73472
rect 10589 73408 10597 73472
rect 10277 73407 10597 73408
rect 3277 72928 3597 72929
rect 3277 72864 3285 72928
rect 3349 72864 3365 72928
rect 3429 72864 3445 72928
rect 3509 72864 3525 72928
rect 3589 72864 3597 72928
rect 3277 72863 3597 72864
rect 7944 72928 8264 72929
rect 7944 72864 7952 72928
rect 8016 72864 8032 72928
rect 8096 72864 8112 72928
rect 8176 72864 8192 72928
rect 8256 72864 8264 72928
rect 7944 72863 8264 72864
rect 5610 72384 5930 72385
rect 5610 72320 5618 72384
rect 5682 72320 5698 72384
rect 5762 72320 5778 72384
rect 5842 72320 5858 72384
rect 5922 72320 5930 72384
rect 5610 72319 5930 72320
rect 10277 72384 10597 72385
rect 10277 72320 10285 72384
rect 10349 72320 10365 72384
rect 10429 72320 10445 72384
rect 10509 72320 10525 72384
rect 10589 72320 10597 72384
rect 10277 72319 10597 72320
rect 3277 71840 3597 71841
rect 3277 71776 3285 71840
rect 3349 71776 3365 71840
rect 3429 71776 3445 71840
rect 3509 71776 3525 71840
rect 3589 71776 3597 71840
rect 3277 71775 3597 71776
rect 7944 71840 8264 71841
rect 7944 71776 7952 71840
rect 8016 71776 8032 71840
rect 8096 71776 8112 71840
rect 8176 71776 8192 71840
rect 8256 71776 8264 71840
rect 7944 71775 8264 71776
rect 105 71634 171 71637
rect 11237 71634 11303 71637
rect 105 71632 11303 71634
rect 105 71576 110 71632
rect 166 71576 11242 71632
rect 11298 71576 11303 71632
rect 105 71574 11303 71576
rect 105 71571 171 71574
rect 11237 71571 11303 71574
rect 11421 71498 11487 71501
rect 13520 71498 14000 71528
rect 11421 71496 14000 71498
rect 11421 71440 11426 71496
rect 11482 71440 14000 71496
rect 11421 71438 14000 71440
rect 11421 71435 11487 71438
rect 13520 71408 14000 71438
rect 5610 71296 5930 71297
rect 5610 71232 5618 71296
rect 5682 71232 5698 71296
rect 5762 71232 5778 71296
rect 5842 71232 5858 71296
rect 5922 71232 5930 71296
rect 5610 71231 5930 71232
rect 10277 71296 10597 71297
rect 10277 71232 10285 71296
rect 10349 71232 10365 71296
rect 10429 71232 10445 71296
rect 10509 71232 10525 71296
rect 10589 71232 10597 71296
rect 10277 71231 10597 71232
rect 3277 70752 3597 70753
rect 3277 70688 3285 70752
rect 3349 70688 3365 70752
rect 3429 70688 3445 70752
rect 3509 70688 3525 70752
rect 3589 70688 3597 70752
rect 3277 70687 3597 70688
rect 7944 70752 8264 70753
rect 7944 70688 7952 70752
rect 8016 70688 8032 70752
rect 8096 70688 8112 70752
rect 8176 70688 8192 70752
rect 8256 70688 8264 70752
rect 7944 70687 8264 70688
rect 5610 70208 5930 70209
rect 5610 70144 5618 70208
rect 5682 70144 5698 70208
rect 5762 70144 5778 70208
rect 5842 70144 5858 70208
rect 5922 70144 5930 70208
rect 5610 70143 5930 70144
rect 10277 70208 10597 70209
rect 10277 70144 10285 70208
rect 10349 70144 10365 70208
rect 10429 70144 10445 70208
rect 10509 70144 10525 70208
rect 10589 70144 10597 70208
rect 10277 70143 10597 70144
rect 3277 69664 3597 69665
rect 3277 69600 3285 69664
rect 3349 69600 3365 69664
rect 3429 69600 3445 69664
rect 3509 69600 3525 69664
rect 3589 69600 3597 69664
rect 3277 69599 3597 69600
rect 7944 69664 8264 69665
rect 7944 69600 7952 69664
rect 8016 69600 8032 69664
rect 8096 69600 8112 69664
rect 8176 69600 8192 69664
rect 8256 69600 8264 69664
rect 7944 69599 8264 69600
rect 5610 69120 5930 69121
rect 5610 69056 5618 69120
rect 5682 69056 5698 69120
rect 5762 69056 5778 69120
rect 5842 69056 5858 69120
rect 5922 69056 5930 69120
rect 5610 69055 5930 69056
rect 10277 69120 10597 69121
rect 10277 69056 10285 69120
rect 10349 69056 10365 69120
rect 10429 69056 10445 69120
rect 10509 69056 10525 69120
rect 10589 69056 10597 69120
rect 10277 69055 10597 69056
rect 3277 68576 3597 68577
rect 3277 68512 3285 68576
rect 3349 68512 3365 68576
rect 3429 68512 3445 68576
rect 3509 68512 3525 68576
rect 3589 68512 3597 68576
rect 3277 68511 3597 68512
rect 7944 68576 8264 68577
rect 7944 68512 7952 68576
rect 8016 68512 8032 68576
rect 8096 68512 8112 68576
rect 8176 68512 8192 68576
rect 8256 68512 8264 68576
rect 7944 68511 8264 68512
rect 5610 68032 5930 68033
rect 5610 67968 5618 68032
rect 5682 67968 5698 68032
rect 5762 67968 5778 68032
rect 5842 67968 5858 68032
rect 5922 67968 5930 68032
rect 5610 67967 5930 67968
rect 10277 68032 10597 68033
rect 10277 67968 10285 68032
rect 10349 67968 10365 68032
rect 10429 67968 10445 68032
rect 10509 67968 10525 68032
rect 10589 67968 10597 68032
rect 10277 67967 10597 67968
rect 3277 67488 3597 67489
rect 3277 67424 3285 67488
rect 3349 67424 3365 67488
rect 3429 67424 3445 67488
rect 3509 67424 3525 67488
rect 3589 67424 3597 67488
rect 3277 67423 3597 67424
rect 7944 67488 8264 67489
rect 7944 67424 7952 67488
rect 8016 67424 8032 67488
rect 8096 67424 8112 67488
rect 8176 67424 8192 67488
rect 8256 67424 8264 67488
rect 7944 67423 8264 67424
rect 5610 66944 5930 66945
rect 5610 66880 5618 66944
rect 5682 66880 5698 66944
rect 5762 66880 5778 66944
rect 5842 66880 5858 66944
rect 5922 66880 5930 66944
rect 5610 66879 5930 66880
rect 10277 66944 10597 66945
rect 10277 66880 10285 66944
rect 10349 66880 10365 66944
rect 10429 66880 10445 66944
rect 10509 66880 10525 66944
rect 10589 66880 10597 66944
rect 10277 66879 10597 66880
rect 3277 66400 3597 66401
rect 3277 66336 3285 66400
rect 3349 66336 3365 66400
rect 3429 66336 3445 66400
rect 3509 66336 3525 66400
rect 3589 66336 3597 66400
rect 3277 66335 3597 66336
rect 7944 66400 8264 66401
rect 7944 66336 7952 66400
rect 8016 66336 8032 66400
rect 8096 66336 8112 66400
rect 8176 66336 8192 66400
rect 8256 66336 8264 66400
rect 7944 66335 8264 66336
rect 5610 65856 5930 65857
rect 5610 65792 5618 65856
rect 5682 65792 5698 65856
rect 5762 65792 5778 65856
rect 5842 65792 5858 65856
rect 5922 65792 5930 65856
rect 5610 65791 5930 65792
rect 10277 65856 10597 65857
rect 10277 65792 10285 65856
rect 10349 65792 10365 65856
rect 10429 65792 10445 65856
rect 10509 65792 10525 65856
rect 10589 65792 10597 65856
rect 10277 65791 10597 65792
rect 3277 65312 3597 65313
rect 3277 65248 3285 65312
rect 3349 65248 3365 65312
rect 3429 65248 3445 65312
rect 3509 65248 3525 65312
rect 3589 65248 3597 65312
rect 3277 65247 3597 65248
rect 7944 65312 8264 65313
rect 7944 65248 7952 65312
rect 8016 65248 8032 65312
rect 8096 65248 8112 65312
rect 8176 65248 8192 65312
rect 8256 65248 8264 65312
rect 7944 65247 8264 65248
rect 5610 64768 5930 64769
rect 5610 64704 5618 64768
rect 5682 64704 5698 64768
rect 5762 64704 5778 64768
rect 5842 64704 5858 64768
rect 5922 64704 5930 64768
rect 5610 64703 5930 64704
rect 10277 64768 10597 64769
rect 10277 64704 10285 64768
rect 10349 64704 10365 64768
rect 10429 64704 10445 64768
rect 10509 64704 10525 64768
rect 10589 64704 10597 64768
rect 10277 64703 10597 64704
rect 11421 64698 11487 64701
rect 13520 64698 14000 64728
rect 11421 64696 14000 64698
rect 11421 64640 11426 64696
rect 11482 64640 14000 64696
rect 11421 64638 14000 64640
rect 11421 64635 11487 64638
rect 13520 64608 14000 64638
rect 3277 64224 3597 64225
rect 3277 64160 3285 64224
rect 3349 64160 3365 64224
rect 3429 64160 3445 64224
rect 3509 64160 3525 64224
rect 3589 64160 3597 64224
rect 3277 64159 3597 64160
rect 7944 64224 8264 64225
rect 7944 64160 7952 64224
rect 8016 64160 8032 64224
rect 8096 64160 8112 64224
rect 8176 64160 8192 64224
rect 8256 64160 8264 64224
rect 7944 64159 8264 64160
rect 5610 63680 5930 63681
rect 5610 63616 5618 63680
rect 5682 63616 5698 63680
rect 5762 63616 5778 63680
rect 5842 63616 5858 63680
rect 5922 63616 5930 63680
rect 5610 63615 5930 63616
rect 10277 63680 10597 63681
rect 10277 63616 10285 63680
rect 10349 63616 10365 63680
rect 10429 63616 10445 63680
rect 10509 63616 10525 63680
rect 10589 63616 10597 63680
rect 10277 63615 10597 63616
rect 3277 63136 3597 63137
rect 3277 63072 3285 63136
rect 3349 63072 3365 63136
rect 3429 63072 3445 63136
rect 3509 63072 3525 63136
rect 3589 63072 3597 63136
rect 3277 63071 3597 63072
rect 7944 63136 8264 63137
rect 7944 63072 7952 63136
rect 8016 63072 8032 63136
rect 8096 63072 8112 63136
rect 8176 63072 8192 63136
rect 8256 63072 8264 63136
rect 7944 63071 8264 63072
rect 5610 62592 5930 62593
rect 5610 62528 5618 62592
rect 5682 62528 5698 62592
rect 5762 62528 5778 62592
rect 5842 62528 5858 62592
rect 5922 62528 5930 62592
rect 5610 62527 5930 62528
rect 10277 62592 10597 62593
rect 10277 62528 10285 62592
rect 10349 62528 10365 62592
rect 10429 62528 10445 62592
rect 10509 62528 10525 62592
rect 10589 62528 10597 62592
rect 10277 62527 10597 62528
rect 3277 62048 3597 62049
rect 3277 61984 3285 62048
rect 3349 61984 3365 62048
rect 3429 61984 3445 62048
rect 3509 61984 3525 62048
rect 3589 61984 3597 62048
rect 3277 61983 3597 61984
rect 7944 62048 8264 62049
rect 7944 61984 7952 62048
rect 8016 61984 8032 62048
rect 8096 61984 8112 62048
rect 8176 61984 8192 62048
rect 8256 61984 8264 62048
rect 7944 61983 8264 61984
rect 5610 61504 5930 61505
rect 5610 61440 5618 61504
rect 5682 61440 5698 61504
rect 5762 61440 5778 61504
rect 5842 61440 5858 61504
rect 5922 61440 5930 61504
rect 5610 61439 5930 61440
rect 10277 61504 10597 61505
rect 10277 61440 10285 61504
rect 10349 61440 10365 61504
rect 10429 61440 10445 61504
rect 10509 61440 10525 61504
rect 10589 61440 10597 61504
rect 10277 61439 10597 61440
rect 0 61296 480 61328
rect 0 61240 110 61296
rect 166 61240 480 61296
rect 0 61208 480 61240
rect 3277 60960 3597 60961
rect 3277 60896 3285 60960
rect 3349 60896 3365 60960
rect 3429 60896 3445 60960
rect 3509 60896 3525 60960
rect 3589 60896 3597 60960
rect 3277 60895 3597 60896
rect 7944 60960 8264 60961
rect 7944 60896 7952 60960
rect 8016 60896 8032 60960
rect 8096 60896 8112 60960
rect 8176 60896 8192 60960
rect 8256 60896 8264 60960
rect 7944 60895 8264 60896
rect 5610 60416 5930 60417
rect 5610 60352 5618 60416
rect 5682 60352 5698 60416
rect 5762 60352 5778 60416
rect 5842 60352 5858 60416
rect 5922 60352 5930 60416
rect 5610 60351 5930 60352
rect 10277 60416 10597 60417
rect 10277 60352 10285 60416
rect 10349 60352 10365 60416
rect 10429 60352 10445 60416
rect 10509 60352 10525 60416
rect 10589 60352 10597 60416
rect 10277 60351 10597 60352
rect 3277 59872 3597 59873
rect 3277 59808 3285 59872
rect 3349 59808 3365 59872
rect 3429 59808 3445 59872
rect 3509 59808 3525 59872
rect 3589 59808 3597 59872
rect 3277 59807 3597 59808
rect 7944 59872 8264 59873
rect 7944 59808 7952 59872
rect 8016 59808 8032 59872
rect 8096 59808 8112 59872
rect 8176 59808 8192 59872
rect 8256 59808 8264 59872
rect 7944 59807 8264 59808
rect 5610 59328 5930 59329
rect 5610 59264 5618 59328
rect 5682 59264 5698 59328
rect 5762 59264 5778 59328
rect 5842 59264 5858 59328
rect 5922 59264 5930 59328
rect 5610 59263 5930 59264
rect 10277 59328 10597 59329
rect 10277 59264 10285 59328
rect 10349 59264 10365 59328
rect 10429 59264 10445 59328
rect 10509 59264 10525 59328
rect 10589 59264 10597 59328
rect 10277 59263 10597 59264
rect 3277 58784 3597 58785
rect 3277 58720 3285 58784
rect 3349 58720 3365 58784
rect 3429 58720 3445 58784
rect 3509 58720 3525 58784
rect 3589 58720 3597 58784
rect 3277 58719 3597 58720
rect 7944 58784 8264 58785
rect 7944 58720 7952 58784
rect 8016 58720 8032 58784
rect 8096 58720 8112 58784
rect 8176 58720 8192 58784
rect 8256 58720 8264 58784
rect 7944 58719 8264 58720
rect 105 58578 171 58581
rect 11237 58578 11303 58581
rect 105 58576 11303 58578
rect 105 58520 110 58576
rect 166 58520 11242 58576
rect 11298 58520 11303 58576
rect 105 58518 11303 58520
rect 105 58515 171 58518
rect 11237 58515 11303 58518
rect 5610 58240 5930 58241
rect 5610 58176 5618 58240
rect 5682 58176 5698 58240
rect 5762 58176 5778 58240
rect 5842 58176 5858 58240
rect 5922 58176 5930 58240
rect 5610 58175 5930 58176
rect 10277 58240 10597 58241
rect 10277 58176 10285 58240
rect 10349 58176 10365 58240
rect 10429 58176 10445 58240
rect 10509 58176 10525 58240
rect 10589 58176 10597 58240
rect 10277 58175 10597 58176
rect 11421 57898 11487 57901
rect 13520 57898 14000 57928
rect 11421 57896 14000 57898
rect 11421 57840 11426 57896
rect 11482 57840 14000 57896
rect 11421 57838 14000 57840
rect 11421 57835 11487 57838
rect 13520 57808 14000 57838
rect 3277 57696 3597 57697
rect 3277 57632 3285 57696
rect 3349 57632 3365 57696
rect 3429 57632 3445 57696
rect 3509 57632 3525 57696
rect 3589 57632 3597 57696
rect 3277 57631 3597 57632
rect 7944 57696 8264 57697
rect 7944 57632 7952 57696
rect 8016 57632 8032 57696
rect 8096 57632 8112 57696
rect 8176 57632 8192 57696
rect 8256 57632 8264 57696
rect 7944 57631 8264 57632
rect 5610 57152 5930 57153
rect 5610 57088 5618 57152
rect 5682 57088 5698 57152
rect 5762 57088 5778 57152
rect 5842 57088 5858 57152
rect 5922 57088 5930 57152
rect 5610 57087 5930 57088
rect 10277 57152 10597 57153
rect 10277 57088 10285 57152
rect 10349 57088 10365 57152
rect 10429 57088 10445 57152
rect 10509 57088 10525 57152
rect 10589 57088 10597 57152
rect 10277 57087 10597 57088
rect 3277 56608 3597 56609
rect 3277 56544 3285 56608
rect 3349 56544 3365 56608
rect 3429 56544 3445 56608
rect 3509 56544 3525 56608
rect 3589 56544 3597 56608
rect 3277 56543 3597 56544
rect 7944 56608 8264 56609
rect 7944 56544 7952 56608
rect 8016 56544 8032 56608
rect 8096 56544 8112 56608
rect 8176 56544 8192 56608
rect 8256 56544 8264 56608
rect 7944 56543 8264 56544
rect 5610 56064 5930 56065
rect 5610 56000 5618 56064
rect 5682 56000 5698 56064
rect 5762 56000 5778 56064
rect 5842 56000 5858 56064
rect 5922 56000 5930 56064
rect 5610 55999 5930 56000
rect 10277 56064 10597 56065
rect 10277 56000 10285 56064
rect 10349 56000 10365 56064
rect 10429 56000 10445 56064
rect 10509 56000 10525 56064
rect 10589 56000 10597 56064
rect 10277 55999 10597 56000
rect 3277 55520 3597 55521
rect 3277 55456 3285 55520
rect 3349 55456 3365 55520
rect 3429 55456 3445 55520
rect 3509 55456 3525 55520
rect 3589 55456 3597 55520
rect 3277 55455 3597 55456
rect 7944 55520 8264 55521
rect 7944 55456 7952 55520
rect 8016 55456 8032 55520
rect 8096 55456 8112 55520
rect 8176 55456 8192 55520
rect 8256 55456 8264 55520
rect 7944 55455 8264 55456
rect 5610 54976 5930 54977
rect 5610 54912 5618 54976
rect 5682 54912 5698 54976
rect 5762 54912 5778 54976
rect 5842 54912 5858 54976
rect 5922 54912 5930 54976
rect 5610 54911 5930 54912
rect 10277 54976 10597 54977
rect 10277 54912 10285 54976
rect 10349 54912 10365 54976
rect 10429 54912 10445 54976
rect 10509 54912 10525 54976
rect 10589 54912 10597 54976
rect 10277 54911 10597 54912
rect 3277 54432 3597 54433
rect 3277 54368 3285 54432
rect 3349 54368 3365 54432
rect 3429 54368 3445 54432
rect 3509 54368 3525 54432
rect 3589 54368 3597 54432
rect 3277 54367 3597 54368
rect 7944 54432 8264 54433
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 54367 8264 54368
rect 5610 53888 5930 53889
rect 5610 53824 5618 53888
rect 5682 53824 5698 53888
rect 5762 53824 5778 53888
rect 5842 53824 5858 53888
rect 5922 53824 5930 53888
rect 5610 53823 5930 53824
rect 10277 53888 10597 53889
rect 10277 53824 10285 53888
rect 10349 53824 10365 53888
rect 10429 53824 10445 53888
rect 10509 53824 10525 53888
rect 10589 53824 10597 53888
rect 10277 53823 10597 53824
rect 3277 53344 3597 53345
rect 3277 53280 3285 53344
rect 3349 53280 3365 53344
rect 3429 53280 3445 53344
rect 3509 53280 3525 53344
rect 3589 53280 3597 53344
rect 3277 53279 3597 53280
rect 7944 53344 8264 53345
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 53279 8264 53280
rect 5610 52800 5930 52801
rect 5610 52736 5618 52800
rect 5682 52736 5698 52800
rect 5762 52736 5778 52800
rect 5842 52736 5858 52800
rect 5922 52736 5930 52800
rect 5610 52735 5930 52736
rect 10277 52800 10597 52801
rect 10277 52736 10285 52800
rect 10349 52736 10365 52800
rect 10429 52736 10445 52800
rect 10509 52736 10525 52800
rect 10589 52736 10597 52800
rect 10277 52735 10597 52736
rect 3277 52256 3597 52257
rect 3277 52192 3285 52256
rect 3349 52192 3365 52256
rect 3429 52192 3445 52256
rect 3509 52192 3525 52256
rect 3589 52192 3597 52256
rect 3277 52191 3597 52192
rect 7944 52256 8264 52257
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 52191 8264 52192
rect 5610 51712 5930 51713
rect 5610 51648 5618 51712
rect 5682 51648 5698 51712
rect 5762 51648 5778 51712
rect 5842 51648 5858 51712
rect 5922 51648 5930 51712
rect 5610 51647 5930 51648
rect 10277 51712 10597 51713
rect 10277 51648 10285 51712
rect 10349 51648 10365 51712
rect 10429 51648 10445 51712
rect 10509 51648 10525 51712
rect 10589 51648 10597 51712
rect 10277 51647 10597 51648
rect 3277 51168 3597 51169
rect 3277 51104 3285 51168
rect 3349 51104 3365 51168
rect 3429 51104 3445 51168
rect 3509 51104 3525 51168
rect 3589 51104 3597 51168
rect 3277 51103 3597 51104
rect 7944 51168 8264 51169
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 51103 8264 51104
rect 11697 51098 11763 51101
rect 13520 51098 14000 51128
rect 11697 51096 14000 51098
rect 11697 51040 11702 51096
rect 11758 51040 14000 51096
rect 11697 51038 14000 51040
rect 11697 51035 11763 51038
rect 13520 51008 14000 51038
rect 5610 50624 5930 50625
rect 5610 50560 5618 50624
rect 5682 50560 5698 50624
rect 5762 50560 5778 50624
rect 5842 50560 5858 50624
rect 5922 50560 5930 50624
rect 5610 50559 5930 50560
rect 10277 50624 10597 50625
rect 10277 50560 10285 50624
rect 10349 50560 10365 50624
rect 10429 50560 10445 50624
rect 10509 50560 10525 50624
rect 10589 50560 10597 50624
rect 10277 50559 10597 50560
rect 3277 50080 3597 50081
rect 3277 50016 3285 50080
rect 3349 50016 3365 50080
rect 3429 50016 3445 50080
rect 3509 50016 3525 50080
rect 3589 50016 3597 50080
rect 3277 50015 3597 50016
rect 7944 50080 8264 50081
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 50015 8264 50016
rect 5610 49536 5930 49537
rect 5610 49472 5618 49536
rect 5682 49472 5698 49536
rect 5762 49472 5778 49536
rect 5842 49472 5858 49536
rect 5922 49472 5930 49536
rect 5610 49471 5930 49472
rect 10277 49536 10597 49537
rect 10277 49472 10285 49536
rect 10349 49472 10365 49536
rect 10429 49472 10445 49536
rect 10509 49472 10525 49536
rect 10589 49472 10597 49536
rect 10277 49471 10597 49472
rect 3277 48992 3597 48993
rect 3277 48928 3285 48992
rect 3349 48928 3365 48992
rect 3429 48928 3445 48992
rect 3509 48928 3525 48992
rect 3589 48928 3597 48992
rect 3277 48927 3597 48928
rect 7944 48992 8264 48993
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 48927 8264 48928
rect 5610 48448 5930 48449
rect 5610 48384 5618 48448
rect 5682 48384 5698 48448
rect 5762 48384 5778 48448
rect 5842 48384 5858 48448
rect 5922 48384 5930 48448
rect 5610 48383 5930 48384
rect 10277 48448 10597 48449
rect 10277 48384 10285 48448
rect 10349 48384 10365 48448
rect 10429 48384 10445 48448
rect 10509 48384 10525 48448
rect 10589 48384 10597 48448
rect 10277 48383 10597 48384
rect 3277 47904 3597 47905
rect 3277 47840 3285 47904
rect 3349 47840 3365 47904
rect 3429 47840 3445 47904
rect 3509 47840 3525 47904
rect 3589 47840 3597 47904
rect 3277 47839 3597 47840
rect 7944 47904 8264 47905
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 47839 8264 47840
rect 0 47696 480 47728
rect 0 47640 110 47696
rect 166 47640 480 47696
rect 0 47608 480 47640
rect 5610 47360 5930 47361
rect 5610 47296 5618 47360
rect 5682 47296 5698 47360
rect 5762 47296 5778 47360
rect 5842 47296 5858 47360
rect 5922 47296 5930 47360
rect 5610 47295 5930 47296
rect 10277 47360 10597 47361
rect 10277 47296 10285 47360
rect 10349 47296 10365 47360
rect 10429 47296 10445 47360
rect 10509 47296 10525 47360
rect 10589 47296 10597 47360
rect 10277 47295 10597 47296
rect 3277 46816 3597 46817
rect 3277 46752 3285 46816
rect 3349 46752 3365 46816
rect 3429 46752 3445 46816
rect 3509 46752 3525 46816
rect 3589 46752 3597 46816
rect 3277 46751 3597 46752
rect 7944 46816 8264 46817
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 46751 8264 46752
rect 5610 46272 5930 46273
rect 5610 46208 5618 46272
rect 5682 46208 5698 46272
rect 5762 46208 5778 46272
rect 5842 46208 5858 46272
rect 5922 46208 5930 46272
rect 5610 46207 5930 46208
rect 10277 46272 10597 46273
rect 10277 46208 10285 46272
rect 10349 46208 10365 46272
rect 10429 46208 10445 46272
rect 10509 46208 10525 46272
rect 10589 46208 10597 46272
rect 10277 46207 10597 46208
rect 3277 45728 3597 45729
rect 3277 45664 3285 45728
rect 3349 45664 3365 45728
rect 3429 45664 3445 45728
rect 3509 45664 3525 45728
rect 3589 45664 3597 45728
rect 3277 45663 3597 45664
rect 7944 45728 8264 45729
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 45663 8264 45664
rect 5610 45184 5930 45185
rect 5610 45120 5618 45184
rect 5682 45120 5698 45184
rect 5762 45120 5778 45184
rect 5842 45120 5858 45184
rect 5922 45120 5930 45184
rect 5610 45119 5930 45120
rect 10277 45184 10597 45185
rect 10277 45120 10285 45184
rect 10349 45120 10365 45184
rect 10429 45120 10445 45184
rect 10509 45120 10525 45184
rect 10589 45120 10597 45184
rect 10277 45119 10597 45120
rect 105 44842 171 44845
rect 11513 44842 11579 44845
rect 105 44840 11579 44842
rect 105 44784 110 44840
rect 166 44784 11518 44840
rect 11574 44784 11579 44840
rect 105 44782 11579 44784
rect 105 44779 171 44782
rect 11513 44779 11579 44782
rect 3277 44640 3597 44641
rect 3277 44576 3285 44640
rect 3349 44576 3365 44640
rect 3429 44576 3445 44640
rect 3509 44576 3525 44640
rect 3589 44576 3597 44640
rect 3277 44575 3597 44576
rect 7944 44640 8264 44641
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 44575 8264 44576
rect 10777 44298 10843 44301
rect 13520 44298 14000 44328
rect 10777 44296 14000 44298
rect 10777 44240 10782 44296
rect 10838 44240 14000 44296
rect 10777 44238 14000 44240
rect 10777 44235 10843 44238
rect 13520 44208 14000 44238
rect 5610 44096 5930 44097
rect 5610 44032 5618 44096
rect 5682 44032 5698 44096
rect 5762 44032 5778 44096
rect 5842 44032 5858 44096
rect 5922 44032 5930 44096
rect 5610 44031 5930 44032
rect 10277 44096 10597 44097
rect 10277 44032 10285 44096
rect 10349 44032 10365 44096
rect 10429 44032 10445 44096
rect 10509 44032 10525 44096
rect 10589 44032 10597 44096
rect 10277 44031 10597 44032
rect 3277 43552 3597 43553
rect 3277 43488 3285 43552
rect 3349 43488 3365 43552
rect 3429 43488 3445 43552
rect 3509 43488 3525 43552
rect 3589 43488 3597 43552
rect 3277 43487 3597 43488
rect 7944 43552 8264 43553
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 43487 8264 43488
rect 5610 43008 5930 43009
rect 5610 42944 5618 43008
rect 5682 42944 5698 43008
rect 5762 42944 5778 43008
rect 5842 42944 5858 43008
rect 5922 42944 5930 43008
rect 5610 42943 5930 42944
rect 10277 43008 10597 43009
rect 10277 42944 10285 43008
rect 10349 42944 10365 43008
rect 10429 42944 10445 43008
rect 10509 42944 10525 43008
rect 10589 42944 10597 43008
rect 10277 42943 10597 42944
rect 3277 42464 3597 42465
rect 3277 42400 3285 42464
rect 3349 42400 3365 42464
rect 3429 42400 3445 42464
rect 3509 42400 3525 42464
rect 3589 42400 3597 42464
rect 3277 42399 3597 42400
rect 7944 42464 8264 42465
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 42399 8264 42400
rect 5610 41920 5930 41921
rect 5610 41856 5618 41920
rect 5682 41856 5698 41920
rect 5762 41856 5778 41920
rect 5842 41856 5858 41920
rect 5922 41856 5930 41920
rect 5610 41855 5930 41856
rect 10277 41920 10597 41921
rect 10277 41856 10285 41920
rect 10349 41856 10365 41920
rect 10429 41856 10445 41920
rect 10509 41856 10525 41920
rect 10589 41856 10597 41920
rect 10277 41855 10597 41856
rect 3277 41376 3597 41377
rect 3277 41312 3285 41376
rect 3349 41312 3365 41376
rect 3429 41312 3445 41376
rect 3509 41312 3525 41376
rect 3589 41312 3597 41376
rect 3277 41311 3597 41312
rect 7944 41376 8264 41377
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 41311 8264 41312
rect 5610 40832 5930 40833
rect 5610 40768 5618 40832
rect 5682 40768 5698 40832
rect 5762 40768 5778 40832
rect 5842 40768 5858 40832
rect 5922 40768 5930 40832
rect 5610 40767 5930 40768
rect 10277 40832 10597 40833
rect 10277 40768 10285 40832
rect 10349 40768 10365 40832
rect 10429 40768 10445 40832
rect 10509 40768 10525 40832
rect 10589 40768 10597 40832
rect 10277 40767 10597 40768
rect 3277 40288 3597 40289
rect 3277 40224 3285 40288
rect 3349 40224 3365 40288
rect 3429 40224 3445 40288
rect 3509 40224 3525 40288
rect 3589 40224 3597 40288
rect 3277 40223 3597 40224
rect 7944 40288 8264 40289
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 40223 8264 40224
rect 5610 39744 5930 39745
rect 5610 39680 5618 39744
rect 5682 39680 5698 39744
rect 5762 39680 5778 39744
rect 5842 39680 5858 39744
rect 5922 39680 5930 39744
rect 5610 39679 5930 39680
rect 10277 39744 10597 39745
rect 10277 39680 10285 39744
rect 10349 39680 10365 39744
rect 10429 39680 10445 39744
rect 10509 39680 10525 39744
rect 10589 39680 10597 39744
rect 10277 39679 10597 39680
rect 3277 39200 3597 39201
rect 3277 39136 3285 39200
rect 3349 39136 3365 39200
rect 3429 39136 3445 39200
rect 3509 39136 3525 39200
rect 3589 39136 3597 39200
rect 3277 39135 3597 39136
rect 7944 39200 8264 39201
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 39135 8264 39136
rect 5610 38656 5930 38657
rect 5610 38592 5618 38656
rect 5682 38592 5698 38656
rect 5762 38592 5778 38656
rect 5842 38592 5858 38656
rect 5922 38592 5930 38656
rect 5610 38591 5930 38592
rect 10277 38656 10597 38657
rect 10277 38592 10285 38656
rect 10349 38592 10365 38656
rect 10429 38592 10445 38656
rect 10509 38592 10525 38656
rect 10589 38592 10597 38656
rect 10277 38591 10597 38592
rect 3277 38112 3597 38113
rect 3277 38048 3285 38112
rect 3349 38048 3365 38112
rect 3429 38048 3445 38112
rect 3509 38048 3525 38112
rect 3589 38048 3597 38112
rect 3277 38047 3597 38048
rect 7944 38112 8264 38113
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 38047 8264 38048
rect 5610 37568 5930 37569
rect 5610 37504 5618 37568
rect 5682 37504 5698 37568
rect 5762 37504 5778 37568
rect 5842 37504 5858 37568
rect 5922 37504 5930 37568
rect 5610 37503 5930 37504
rect 10277 37568 10597 37569
rect 10277 37504 10285 37568
rect 10349 37504 10365 37568
rect 10429 37504 10445 37568
rect 10509 37504 10525 37568
rect 10589 37504 10597 37568
rect 10277 37503 10597 37504
rect 11421 37498 11487 37501
rect 13520 37498 14000 37528
rect 11421 37496 14000 37498
rect 11421 37440 11426 37496
rect 11482 37440 14000 37496
rect 11421 37438 14000 37440
rect 11421 37435 11487 37438
rect 13520 37408 14000 37438
rect 3277 37024 3597 37025
rect 3277 36960 3285 37024
rect 3349 36960 3365 37024
rect 3429 36960 3445 37024
rect 3509 36960 3525 37024
rect 3589 36960 3597 37024
rect 3277 36959 3597 36960
rect 7944 37024 8264 37025
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 36959 8264 36960
rect 5610 36480 5930 36481
rect 5610 36416 5618 36480
rect 5682 36416 5698 36480
rect 5762 36416 5778 36480
rect 5842 36416 5858 36480
rect 5922 36416 5930 36480
rect 5610 36415 5930 36416
rect 10277 36480 10597 36481
rect 10277 36416 10285 36480
rect 10349 36416 10365 36480
rect 10429 36416 10445 36480
rect 10509 36416 10525 36480
rect 10589 36416 10597 36480
rect 10277 36415 10597 36416
rect 3277 35936 3597 35937
rect 3277 35872 3285 35936
rect 3349 35872 3365 35936
rect 3429 35872 3445 35936
rect 3509 35872 3525 35936
rect 3589 35872 3597 35936
rect 3277 35871 3597 35872
rect 7944 35936 8264 35937
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 35871 8264 35872
rect 5610 35392 5930 35393
rect 5610 35328 5618 35392
rect 5682 35328 5698 35392
rect 5762 35328 5778 35392
rect 5842 35328 5858 35392
rect 5922 35328 5930 35392
rect 5610 35327 5930 35328
rect 10277 35392 10597 35393
rect 10277 35328 10285 35392
rect 10349 35328 10365 35392
rect 10429 35328 10445 35392
rect 10509 35328 10525 35392
rect 10589 35328 10597 35392
rect 10277 35327 10597 35328
rect 3277 34848 3597 34849
rect 3277 34784 3285 34848
rect 3349 34784 3365 34848
rect 3429 34784 3445 34848
rect 3509 34784 3525 34848
rect 3589 34784 3597 34848
rect 3277 34783 3597 34784
rect 7944 34848 8264 34849
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 34783 8264 34784
rect 5610 34304 5930 34305
rect 5610 34240 5618 34304
rect 5682 34240 5698 34304
rect 5762 34240 5778 34304
rect 5842 34240 5858 34304
rect 5922 34240 5930 34304
rect 5610 34239 5930 34240
rect 10277 34304 10597 34305
rect 10277 34240 10285 34304
rect 10349 34240 10365 34304
rect 10429 34240 10445 34304
rect 10509 34240 10525 34304
rect 10589 34240 10597 34304
rect 10277 34239 10597 34240
rect 0 34096 480 34128
rect 0 34040 110 34096
rect 166 34040 480 34096
rect 0 34008 480 34040
rect 3277 33760 3597 33761
rect 3277 33696 3285 33760
rect 3349 33696 3365 33760
rect 3429 33696 3445 33760
rect 3509 33696 3525 33760
rect 3589 33696 3597 33760
rect 3277 33695 3597 33696
rect 7944 33760 8264 33761
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 33695 8264 33696
rect 5610 33216 5930 33217
rect 5610 33152 5618 33216
rect 5682 33152 5698 33216
rect 5762 33152 5778 33216
rect 5842 33152 5858 33216
rect 5922 33152 5930 33216
rect 5610 33151 5930 33152
rect 10277 33216 10597 33217
rect 10277 33152 10285 33216
rect 10349 33152 10365 33216
rect 10429 33152 10445 33216
rect 10509 33152 10525 33216
rect 10589 33152 10597 33216
rect 10277 33151 10597 33152
rect 3277 32672 3597 32673
rect 3277 32608 3285 32672
rect 3349 32608 3365 32672
rect 3429 32608 3445 32672
rect 3509 32608 3525 32672
rect 3589 32608 3597 32672
rect 3277 32607 3597 32608
rect 7944 32672 8264 32673
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 32607 8264 32608
rect 5610 32128 5930 32129
rect 5610 32064 5618 32128
rect 5682 32064 5698 32128
rect 5762 32064 5778 32128
rect 5842 32064 5858 32128
rect 5922 32064 5930 32128
rect 5610 32063 5930 32064
rect 10277 32128 10597 32129
rect 10277 32064 10285 32128
rect 10349 32064 10365 32128
rect 10429 32064 10445 32128
rect 10509 32064 10525 32128
rect 10589 32064 10597 32128
rect 10277 32063 10597 32064
rect 3277 31584 3597 31585
rect 3277 31520 3285 31584
rect 3349 31520 3365 31584
rect 3429 31520 3445 31584
rect 3509 31520 3525 31584
rect 3589 31520 3597 31584
rect 3277 31519 3597 31520
rect 7944 31584 8264 31585
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 31519 8264 31520
rect 105 31242 171 31245
rect 10961 31242 11027 31245
rect 105 31240 11027 31242
rect 105 31184 110 31240
rect 166 31184 10966 31240
rect 11022 31184 11027 31240
rect 105 31182 11027 31184
rect 105 31179 171 31182
rect 10961 31179 11027 31182
rect 5610 31040 5930 31041
rect 5610 30976 5618 31040
rect 5682 30976 5698 31040
rect 5762 30976 5778 31040
rect 5842 30976 5858 31040
rect 5922 30976 5930 31040
rect 5610 30975 5930 30976
rect 10277 31040 10597 31041
rect 10277 30976 10285 31040
rect 10349 30976 10365 31040
rect 10429 30976 10445 31040
rect 10509 30976 10525 31040
rect 10589 30976 10597 31040
rect 10277 30975 10597 30976
rect 10777 30698 10843 30701
rect 13520 30698 14000 30728
rect 10777 30696 14000 30698
rect 10777 30640 10782 30696
rect 10838 30640 14000 30696
rect 10777 30638 14000 30640
rect 10777 30635 10843 30638
rect 13520 30608 14000 30638
rect 3277 30496 3597 30497
rect 3277 30432 3285 30496
rect 3349 30432 3365 30496
rect 3429 30432 3445 30496
rect 3509 30432 3525 30496
rect 3589 30432 3597 30496
rect 3277 30431 3597 30432
rect 7944 30496 8264 30497
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 30431 8264 30432
rect 5610 29952 5930 29953
rect 5610 29888 5618 29952
rect 5682 29888 5698 29952
rect 5762 29888 5778 29952
rect 5842 29888 5858 29952
rect 5922 29888 5930 29952
rect 5610 29887 5930 29888
rect 10277 29952 10597 29953
rect 10277 29888 10285 29952
rect 10349 29888 10365 29952
rect 10429 29888 10445 29952
rect 10509 29888 10525 29952
rect 10589 29888 10597 29952
rect 10277 29887 10597 29888
rect 3277 29408 3597 29409
rect 3277 29344 3285 29408
rect 3349 29344 3365 29408
rect 3429 29344 3445 29408
rect 3509 29344 3525 29408
rect 3589 29344 3597 29408
rect 3277 29343 3597 29344
rect 7944 29408 8264 29409
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 29343 8264 29344
rect 5610 28864 5930 28865
rect 5610 28800 5618 28864
rect 5682 28800 5698 28864
rect 5762 28800 5778 28864
rect 5842 28800 5858 28864
rect 5922 28800 5930 28864
rect 5610 28799 5930 28800
rect 10277 28864 10597 28865
rect 10277 28800 10285 28864
rect 10349 28800 10365 28864
rect 10429 28800 10445 28864
rect 10509 28800 10525 28864
rect 10589 28800 10597 28864
rect 10277 28799 10597 28800
rect 3277 28320 3597 28321
rect 3277 28256 3285 28320
rect 3349 28256 3365 28320
rect 3429 28256 3445 28320
rect 3509 28256 3525 28320
rect 3589 28256 3597 28320
rect 3277 28255 3597 28256
rect 7944 28320 8264 28321
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 28255 8264 28256
rect 5610 27776 5930 27777
rect 5610 27712 5618 27776
rect 5682 27712 5698 27776
rect 5762 27712 5778 27776
rect 5842 27712 5858 27776
rect 5922 27712 5930 27776
rect 5610 27711 5930 27712
rect 10277 27776 10597 27777
rect 10277 27712 10285 27776
rect 10349 27712 10365 27776
rect 10429 27712 10445 27776
rect 10509 27712 10525 27776
rect 10589 27712 10597 27776
rect 10277 27711 10597 27712
rect 3277 27232 3597 27233
rect 3277 27168 3285 27232
rect 3349 27168 3365 27232
rect 3429 27168 3445 27232
rect 3509 27168 3525 27232
rect 3589 27168 3597 27232
rect 3277 27167 3597 27168
rect 7944 27232 8264 27233
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 27167 8264 27168
rect 5610 26688 5930 26689
rect 5610 26624 5618 26688
rect 5682 26624 5698 26688
rect 5762 26624 5778 26688
rect 5842 26624 5858 26688
rect 5922 26624 5930 26688
rect 5610 26623 5930 26624
rect 10277 26688 10597 26689
rect 10277 26624 10285 26688
rect 10349 26624 10365 26688
rect 10429 26624 10445 26688
rect 10509 26624 10525 26688
rect 10589 26624 10597 26688
rect 10277 26623 10597 26624
rect 3277 26144 3597 26145
rect 3277 26080 3285 26144
rect 3349 26080 3365 26144
rect 3429 26080 3445 26144
rect 3509 26080 3525 26144
rect 3589 26080 3597 26144
rect 3277 26079 3597 26080
rect 7944 26144 8264 26145
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 26079 8264 26080
rect 5610 25600 5930 25601
rect 5610 25536 5618 25600
rect 5682 25536 5698 25600
rect 5762 25536 5778 25600
rect 5842 25536 5858 25600
rect 5922 25536 5930 25600
rect 5610 25535 5930 25536
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 3277 25056 3597 25057
rect 3277 24992 3285 25056
rect 3349 24992 3365 25056
rect 3429 24992 3445 25056
rect 3509 24992 3525 25056
rect 3589 24992 3597 25056
rect 3277 24991 3597 24992
rect 7944 25056 8264 25057
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 24991 8264 24992
rect 5610 24512 5930 24513
rect 5610 24448 5618 24512
rect 5682 24448 5698 24512
rect 5762 24448 5778 24512
rect 5842 24448 5858 24512
rect 5922 24448 5930 24512
rect 5610 24447 5930 24448
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 3277 23968 3597 23969
rect 3277 23904 3285 23968
rect 3349 23904 3365 23968
rect 3429 23904 3445 23968
rect 3509 23904 3525 23968
rect 3589 23904 3597 23968
rect 3277 23903 3597 23904
rect 7944 23968 8264 23969
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 23903 8264 23904
rect 10685 23898 10751 23901
rect 13520 23898 14000 23928
rect 10685 23896 14000 23898
rect 10685 23840 10690 23896
rect 10746 23840 14000 23896
rect 10685 23838 14000 23840
rect 10685 23835 10751 23838
rect 13520 23808 14000 23838
rect 5610 23424 5930 23425
rect 5610 23360 5618 23424
rect 5682 23360 5698 23424
rect 5762 23360 5778 23424
rect 5842 23360 5858 23424
rect 5922 23360 5930 23424
rect 5610 23359 5930 23360
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 3277 22880 3597 22881
rect 3277 22816 3285 22880
rect 3349 22816 3365 22880
rect 3429 22816 3445 22880
rect 3509 22816 3525 22880
rect 3589 22816 3597 22880
rect 3277 22815 3597 22816
rect 7944 22880 8264 22881
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 22815 8264 22816
rect 5610 22336 5930 22337
rect 5610 22272 5618 22336
rect 5682 22272 5698 22336
rect 5762 22272 5778 22336
rect 5842 22272 5858 22336
rect 5922 22272 5930 22336
rect 5610 22271 5930 22272
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 3277 21792 3597 21793
rect 3277 21728 3285 21792
rect 3349 21728 3365 21792
rect 3429 21728 3445 21792
rect 3509 21728 3525 21792
rect 3589 21728 3597 21792
rect 3277 21727 3597 21728
rect 7944 21792 8264 21793
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 21727 8264 21728
rect 5610 21248 5930 21249
rect 5610 21184 5618 21248
rect 5682 21184 5698 21248
rect 5762 21184 5778 21248
rect 5842 21184 5858 21248
rect 5922 21184 5930 21248
rect 5610 21183 5930 21184
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 3277 20704 3597 20705
rect 3277 20640 3285 20704
rect 3349 20640 3365 20704
rect 3429 20640 3445 20704
rect 3509 20640 3525 20704
rect 3589 20640 3597 20704
rect 3277 20639 3597 20640
rect 7944 20704 8264 20705
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 20639 8264 20640
rect 0 20496 480 20528
rect 0 20440 110 20496
rect 166 20440 480 20496
rect 0 20408 480 20440
rect 5610 20160 5930 20161
rect 5610 20096 5618 20160
rect 5682 20096 5698 20160
rect 5762 20096 5778 20160
rect 5842 20096 5858 20160
rect 5922 20096 5930 20160
rect 5610 20095 5930 20096
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 3277 19616 3597 19617
rect 3277 19552 3285 19616
rect 3349 19552 3365 19616
rect 3429 19552 3445 19616
rect 3509 19552 3525 19616
rect 3589 19552 3597 19616
rect 3277 19551 3597 19552
rect 7944 19616 8264 19617
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 19551 8264 19552
rect 5610 19072 5930 19073
rect 5610 19008 5618 19072
rect 5682 19008 5698 19072
rect 5762 19008 5778 19072
rect 5842 19008 5858 19072
rect 5922 19008 5930 19072
rect 5610 19007 5930 19008
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 3277 18528 3597 18529
rect 3277 18464 3285 18528
rect 3349 18464 3365 18528
rect 3429 18464 3445 18528
rect 3509 18464 3525 18528
rect 3589 18464 3597 18528
rect 3277 18463 3597 18464
rect 7944 18528 8264 18529
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 18463 8264 18464
rect 5610 17984 5930 17985
rect 5610 17920 5618 17984
rect 5682 17920 5698 17984
rect 5762 17920 5778 17984
rect 5842 17920 5858 17984
rect 5922 17920 5930 17984
rect 5610 17919 5930 17920
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 3277 17440 3597 17441
rect 3277 17376 3285 17440
rect 3349 17376 3365 17440
rect 3429 17376 3445 17440
rect 3509 17376 3525 17440
rect 3589 17376 3597 17440
rect 3277 17375 3597 17376
rect 7944 17440 8264 17441
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 17375 8264 17376
rect 105 17234 171 17237
rect 11237 17234 11303 17237
rect 105 17232 11303 17234
rect 105 17176 110 17232
rect 166 17176 11242 17232
rect 11298 17176 11303 17232
rect 105 17174 11303 17176
rect 105 17171 171 17174
rect 11237 17171 11303 17174
rect 11145 17098 11211 17101
rect 13520 17098 14000 17128
rect 11145 17096 14000 17098
rect 11145 17040 11150 17096
rect 11206 17040 14000 17096
rect 11145 17038 14000 17040
rect 11145 17035 11211 17038
rect 13520 17008 14000 17038
rect 5610 16896 5930 16897
rect 5610 16832 5618 16896
rect 5682 16832 5698 16896
rect 5762 16832 5778 16896
rect 5842 16832 5858 16896
rect 5922 16832 5930 16896
rect 5610 16831 5930 16832
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 3277 16352 3597 16353
rect 3277 16288 3285 16352
rect 3349 16288 3365 16352
rect 3429 16288 3445 16352
rect 3509 16288 3525 16352
rect 3589 16288 3597 16352
rect 3277 16287 3597 16288
rect 7944 16352 8264 16353
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 16287 8264 16288
rect 5610 15808 5930 15809
rect 5610 15744 5618 15808
rect 5682 15744 5698 15808
rect 5762 15744 5778 15808
rect 5842 15744 5858 15808
rect 5922 15744 5930 15808
rect 5610 15743 5930 15744
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 3277 15264 3597 15265
rect 3277 15200 3285 15264
rect 3349 15200 3365 15264
rect 3429 15200 3445 15264
rect 3509 15200 3525 15264
rect 3589 15200 3597 15264
rect 3277 15199 3597 15200
rect 7944 15264 8264 15265
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 15199 8264 15200
rect 5610 14720 5930 14721
rect 5610 14656 5618 14720
rect 5682 14656 5698 14720
rect 5762 14656 5778 14720
rect 5842 14656 5858 14720
rect 5922 14656 5930 14720
rect 5610 14655 5930 14656
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 3277 14176 3597 14177
rect 3277 14112 3285 14176
rect 3349 14112 3365 14176
rect 3429 14112 3445 14176
rect 3509 14112 3525 14176
rect 3589 14112 3597 14176
rect 3277 14111 3597 14112
rect 7944 14176 8264 14177
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 14111 8264 14112
rect 5610 13632 5930 13633
rect 5610 13568 5618 13632
rect 5682 13568 5698 13632
rect 5762 13568 5778 13632
rect 5842 13568 5858 13632
rect 5922 13568 5930 13632
rect 5610 13567 5930 13568
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 3277 13088 3597 13089
rect 3277 13024 3285 13088
rect 3349 13024 3365 13088
rect 3429 13024 3445 13088
rect 3509 13024 3525 13088
rect 3589 13024 3597 13088
rect 3277 13023 3597 13024
rect 7944 13088 8264 13089
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 13023 8264 13024
rect 5610 12544 5930 12545
rect 5610 12480 5618 12544
rect 5682 12480 5698 12544
rect 5762 12480 5778 12544
rect 5842 12480 5858 12544
rect 5922 12480 5930 12544
rect 5610 12479 5930 12480
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 3277 12000 3597 12001
rect 3277 11936 3285 12000
rect 3349 11936 3365 12000
rect 3429 11936 3445 12000
rect 3509 11936 3525 12000
rect 3589 11936 3597 12000
rect 3277 11935 3597 11936
rect 7944 12000 8264 12001
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 11935 8264 11936
rect 5610 11456 5930 11457
rect 5610 11392 5618 11456
rect 5682 11392 5698 11456
rect 5762 11392 5778 11456
rect 5842 11392 5858 11456
rect 5922 11392 5930 11456
rect 5610 11391 5930 11392
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 3277 10912 3597 10913
rect 3277 10848 3285 10912
rect 3349 10848 3365 10912
rect 3429 10848 3445 10912
rect 3509 10848 3525 10912
rect 3589 10848 3597 10912
rect 3277 10847 3597 10848
rect 7944 10912 8264 10913
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 10847 8264 10848
rect 5610 10368 5930 10369
rect 5610 10304 5618 10368
rect 5682 10304 5698 10368
rect 5762 10304 5778 10368
rect 5842 10304 5858 10368
rect 5922 10304 5930 10368
rect 5610 10303 5930 10304
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 11421 10298 11487 10301
rect 13520 10298 14000 10328
rect 11421 10296 14000 10298
rect 11421 10240 11426 10296
rect 11482 10240 14000 10296
rect 11421 10238 14000 10240
rect 11421 10235 11487 10238
rect 13520 10208 14000 10238
rect 3277 9824 3597 9825
rect 3277 9760 3285 9824
rect 3349 9760 3365 9824
rect 3429 9760 3445 9824
rect 3509 9760 3525 9824
rect 3589 9760 3597 9824
rect 3277 9759 3597 9760
rect 7944 9824 8264 9825
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 9759 8264 9760
rect 5610 9280 5930 9281
rect 5610 9216 5618 9280
rect 5682 9216 5698 9280
rect 5762 9216 5778 9280
rect 5842 9216 5858 9280
rect 5922 9216 5930 9280
rect 5610 9215 5930 9216
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 3277 8736 3597 8737
rect 3277 8672 3285 8736
rect 3349 8672 3365 8736
rect 3429 8672 3445 8736
rect 3509 8672 3525 8736
rect 3589 8672 3597 8736
rect 3277 8671 3597 8672
rect 7944 8736 8264 8737
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 8671 8264 8672
rect 5610 8192 5930 8193
rect 5610 8128 5618 8192
rect 5682 8128 5698 8192
rect 5762 8128 5778 8192
rect 5842 8128 5858 8192
rect 5922 8128 5930 8192
rect 5610 8127 5930 8128
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 3277 7648 3597 7649
rect 3277 7584 3285 7648
rect 3349 7584 3365 7648
rect 3429 7584 3445 7648
rect 3509 7584 3525 7648
rect 3589 7584 3597 7648
rect 3277 7583 3597 7584
rect 7944 7648 8264 7649
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 7583 8264 7584
rect 5610 7104 5930 7105
rect 5610 7040 5618 7104
rect 5682 7040 5698 7104
rect 5762 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5930 7104
rect 5610 7039 5930 7040
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 0 6896 480 6928
rect 0 6840 110 6896
rect 166 6840 480 6896
rect 0 6808 480 6840
rect 3277 6560 3597 6561
rect 3277 6496 3285 6560
rect 3349 6496 3365 6560
rect 3429 6496 3445 6560
rect 3509 6496 3525 6560
rect 3589 6496 3597 6560
rect 3277 6495 3597 6496
rect 7944 6560 8264 6561
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 6495 8264 6496
rect 5610 6016 5930 6017
rect 5610 5952 5618 6016
rect 5682 5952 5698 6016
rect 5762 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5930 6016
rect 5610 5951 5930 5952
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 105 5674 171 5677
rect 11237 5674 11303 5677
rect 105 5672 11303 5674
rect 105 5616 110 5672
rect 166 5616 11242 5672
rect 11298 5616 11303 5672
rect 105 5614 11303 5616
rect 105 5611 171 5614
rect 11237 5611 11303 5614
rect 3277 5472 3597 5473
rect 3277 5408 3285 5472
rect 3349 5408 3365 5472
rect 3429 5408 3445 5472
rect 3509 5408 3525 5472
rect 3589 5408 3597 5472
rect 3277 5407 3597 5408
rect 7944 5472 8264 5473
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 5407 8264 5408
rect 5610 4928 5930 4929
rect 5610 4864 5618 4928
rect 5682 4864 5698 4928
rect 5762 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5930 4928
rect 5610 4863 5930 4864
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 3277 4384 3597 4385
rect 3277 4320 3285 4384
rect 3349 4320 3365 4384
rect 3429 4320 3445 4384
rect 3509 4320 3525 4384
rect 3589 4320 3597 4384
rect 3277 4319 3597 4320
rect 7944 4384 8264 4385
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 4319 8264 4320
rect 5610 3840 5930 3841
rect 5610 3776 5618 3840
rect 5682 3776 5698 3840
rect 5762 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5930 3840
rect 5610 3775 5930 3776
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 10961 3498 11027 3501
rect 13520 3498 14000 3528
rect 10961 3496 14000 3498
rect 10961 3440 10966 3496
rect 11022 3440 14000 3496
rect 10961 3438 14000 3440
rect 10961 3435 11027 3438
rect 13520 3408 14000 3438
rect 3277 3296 3597 3297
rect 3277 3232 3285 3296
rect 3349 3232 3365 3296
rect 3429 3232 3445 3296
rect 3509 3232 3525 3296
rect 3589 3232 3597 3296
rect 3277 3231 3597 3232
rect 7944 3296 8264 3297
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 3231 8264 3232
rect 5610 2752 5930 2753
rect 5610 2688 5618 2752
rect 5682 2688 5698 2752
rect 5762 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5930 2752
rect 5610 2687 5930 2688
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 3277 2208 3597 2209
rect 3277 2144 3285 2208
rect 3349 2144 3365 2208
rect 3429 2144 3445 2208
rect 3509 2144 3525 2208
rect 3589 2144 3597 2208
rect 3277 2143 3597 2144
rect 7944 2208 8264 2209
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2143 8264 2144
<< via3 >>
rect 3285 106652 3349 106656
rect 3285 106596 3289 106652
rect 3289 106596 3345 106652
rect 3345 106596 3349 106652
rect 3285 106592 3349 106596
rect 3365 106652 3429 106656
rect 3365 106596 3369 106652
rect 3369 106596 3425 106652
rect 3425 106596 3429 106652
rect 3365 106592 3429 106596
rect 3445 106652 3509 106656
rect 3445 106596 3449 106652
rect 3449 106596 3505 106652
rect 3505 106596 3509 106652
rect 3445 106592 3509 106596
rect 3525 106652 3589 106656
rect 3525 106596 3529 106652
rect 3529 106596 3585 106652
rect 3585 106596 3589 106652
rect 3525 106592 3589 106596
rect 7952 106652 8016 106656
rect 7952 106596 7956 106652
rect 7956 106596 8012 106652
rect 8012 106596 8016 106652
rect 7952 106592 8016 106596
rect 8032 106652 8096 106656
rect 8032 106596 8036 106652
rect 8036 106596 8092 106652
rect 8092 106596 8096 106652
rect 8032 106592 8096 106596
rect 8112 106652 8176 106656
rect 8112 106596 8116 106652
rect 8116 106596 8172 106652
rect 8172 106596 8176 106652
rect 8112 106592 8176 106596
rect 8192 106652 8256 106656
rect 8192 106596 8196 106652
rect 8196 106596 8252 106652
rect 8252 106596 8256 106652
rect 8192 106592 8256 106596
rect 5618 106108 5682 106112
rect 5618 106052 5622 106108
rect 5622 106052 5678 106108
rect 5678 106052 5682 106108
rect 5618 106048 5682 106052
rect 5698 106108 5762 106112
rect 5698 106052 5702 106108
rect 5702 106052 5758 106108
rect 5758 106052 5762 106108
rect 5698 106048 5762 106052
rect 5778 106108 5842 106112
rect 5778 106052 5782 106108
rect 5782 106052 5838 106108
rect 5838 106052 5842 106108
rect 5778 106048 5842 106052
rect 5858 106108 5922 106112
rect 5858 106052 5862 106108
rect 5862 106052 5918 106108
rect 5918 106052 5922 106108
rect 5858 106048 5922 106052
rect 10285 106108 10349 106112
rect 10285 106052 10289 106108
rect 10289 106052 10345 106108
rect 10345 106052 10349 106108
rect 10285 106048 10349 106052
rect 10365 106108 10429 106112
rect 10365 106052 10369 106108
rect 10369 106052 10425 106108
rect 10425 106052 10429 106108
rect 10365 106048 10429 106052
rect 10445 106108 10509 106112
rect 10445 106052 10449 106108
rect 10449 106052 10505 106108
rect 10505 106052 10509 106108
rect 10445 106048 10509 106052
rect 10525 106108 10589 106112
rect 10525 106052 10529 106108
rect 10529 106052 10585 106108
rect 10585 106052 10589 106108
rect 10525 106048 10589 106052
rect 3285 105564 3349 105568
rect 3285 105508 3289 105564
rect 3289 105508 3345 105564
rect 3345 105508 3349 105564
rect 3285 105504 3349 105508
rect 3365 105564 3429 105568
rect 3365 105508 3369 105564
rect 3369 105508 3425 105564
rect 3425 105508 3429 105564
rect 3365 105504 3429 105508
rect 3445 105564 3509 105568
rect 3445 105508 3449 105564
rect 3449 105508 3505 105564
rect 3505 105508 3509 105564
rect 3445 105504 3509 105508
rect 3525 105564 3589 105568
rect 3525 105508 3529 105564
rect 3529 105508 3585 105564
rect 3585 105508 3589 105564
rect 3525 105504 3589 105508
rect 7952 105564 8016 105568
rect 7952 105508 7956 105564
rect 7956 105508 8012 105564
rect 8012 105508 8016 105564
rect 7952 105504 8016 105508
rect 8032 105564 8096 105568
rect 8032 105508 8036 105564
rect 8036 105508 8092 105564
rect 8092 105508 8096 105564
rect 8032 105504 8096 105508
rect 8112 105564 8176 105568
rect 8112 105508 8116 105564
rect 8116 105508 8172 105564
rect 8172 105508 8176 105564
rect 8112 105504 8176 105508
rect 8192 105564 8256 105568
rect 8192 105508 8196 105564
rect 8196 105508 8252 105564
rect 8252 105508 8256 105564
rect 8192 105504 8256 105508
rect 5618 105020 5682 105024
rect 5618 104964 5622 105020
rect 5622 104964 5678 105020
rect 5678 104964 5682 105020
rect 5618 104960 5682 104964
rect 5698 105020 5762 105024
rect 5698 104964 5702 105020
rect 5702 104964 5758 105020
rect 5758 104964 5762 105020
rect 5698 104960 5762 104964
rect 5778 105020 5842 105024
rect 5778 104964 5782 105020
rect 5782 104964 5838 105020
rect 5838 104964 5842 105020
rect 5778 104960 5842 104964
rect 5858 105020 5922 105024
rect 5858 104964 5862 105020
rect 5862 104964 5918 105020
rect 5918 104964 5922 105020
rect 5858 104960 5922 104964
rect 10285 105020 10349 105024
rect 10285 104964 10289 105020
rect 10289 104964 10345 105020
rect 10345 104964 10349 105020
rect 10285 104960 10349 104964
rect 10365 105020 10429 105024
rect 10365 104964 10369 105020
rect 10369 104964 10425 105020
rect 10425 104964 10429 105020
rect 10365 104960 10429 104964
rect 10445 105020 10509 105024
rect 10445 104964 10449 105020
rect 10449 104964 10505 105020
rect 10505 104964 10509 105020
rect 10445 104960 10509 104964
rect 10525 105020 10589 105024
rect 10525 104964 10529 105020
rect 10529 104964 10585 105020
rect 10585 104964 10589 105020
rect 10525 104960 10589 104964
rect 3285 104476 3349 104480
rect 3285 104420 3289 104476
rect 3289 104420 3345 104476
rect 3345 104420 3349 104476
rect 3285 104416 3349 104420
rect 3365 104476 3429 104480
rect 3365 104420 3369 104476
rect 3369 104420 3425 104476
rect 3425 104420 3429 104476
rect 3365 104416 3429 104420
rect 3445 104476 3509 104480
rect 3445 104420 3449 104476
rect 3449 104420 3505 104476
rect 3505 104420 3509 104476
rect 3445 104416 3509 104420
rect 3525 104476 3589 104480
rect 3525 104420 3529 104476
rect 3529 104420 3585 104476
rect 3585 104420 3589 104476
rect 3525 104416 3589 104420
rect 7952 104476 8016 104480
rect 7952 104420 7956 104476
rect 7956 104420 8012 104476
rect 8012 104420 8016 104476
rect 7952 104416 8016 104420
rect 8032 104476 8096 104480
rect 8032 104420 8036 104476
rect 8036 104420 8092 104476
rect 8092 104420 8096 104476
rect 8032 104416 8096 104420
rect 8112 104476 8176 104480
rect 8112 104420 8116 104476
rect 8116 104420 8172 104476
rect 8172 104420 8176 104476
rect 8112 104416 8176 104420
rect 8192 104476 8256 104480
rect 8192 104420 8196 104476
rect 8196 104420 8252 104476
rect 8252 104420 8256 104476
rect 8192 104416 8256 104420
rect 5618 103932 5682 103936
rect 5618 103876 5622 103932
rect 5622 103876 5678 103932
rect 5678 103876 5682 103932
rect 5618 103872 5682 103876
rect 5698 103932 5762 103936
rect 5698 103876 5702 103932
rect 5702 103876 5758 103932
rect 5758 103876 5762 103932
rect 5698 103872 5762 103876
rect 5778 103932 5842 103936
rect 5778 103876 5782 103932
rect 5782 103876 5838 103932
rect 5838 103876 5842 103932
rect 5778 103872 5842 103876
rect 5858 103932 5922 103936
rect 5858 103876 5862 103932
rect 5862 103876 5918 103932
rect 5918 103876 5922 103932
rect 5858 103872 5922 103876
rect 10285 103932 10349 103936
rect 10285 103876 10289 103932
rect 10289 103876 10345 103932
rect 10345 103876 10349 103932
rect 10285 103872 10349 103876
rect 10365 103932 10429 103936
rect 10365 103876 10369 103932
rect 10369 103876 10425 103932
rect 10425 103876 10429 103932
rect 10365 103872 10429 103876
rect 10445 103932 10509 103936
rect 10445 103876 10449 103932
rect 10449 103876 10505 103932
rect 10505 103876 10509 103932
rect 10445 103872 10509 103876
rect 10525 103932 10589 103936
rect 10525 103876 10529 103932
rect 10529 103876 10585 103932
rect 10585 103876 10589 103932
rect 10525 103872 10589 103876
rect 3285 103388 3349 103392
rect 3285 103332 3289 103388
rect 3289 103332 3345 103388
rect 3345 103332 3349 103388
rect 3285 103328 3349 103332
rect 3365 103388 3429 103392
rect 3365 103332 3369 103388
rect 3369 103332 3425 103388
rect 3425 103332 3429 103388
rect 3365 103328 3429 103332
rect 3445 103388 3509 103392
rect 3445 103332 3449 103388
rect 3449 103332 3505 103388
rect 3505 103332 3509 103388
rect 3445 103328 3509 103332
rect 3525 103388 3589 103392
rect 3525 103332 3529 103388
rect 3529 103332 3585 103388
rect 3585 103332 3589 103388
rect 3525 103328 3589 103332
rect 7952 103388 8016 103392
rect 7952 103332 7956 103388
rect 7956 103332 8012 103388
rect 8012 103332 8016 103388
rect 7952 103328 8016 103332
rect 8032 103388 8096 103392
rect 8032 103332 8036 103388
rect 8036 103332 8092 103388
rect 8092 103332 8096 103388
rect 8032 103328 8096 103332
rect 8112 103388 8176 103392
rect 8112 103332 8116 103388
rect 8116 103332 8172 103388
rect 8172 103332 8176 103388
rect 8112 103328 8176 103332
rect 8192 103388 8256 103392
rect 8192 103332 8196 103388
rect 8196 103332 8252 103388
rect 8252 103332 8256 103388
rect 8192 103328 8256 103332
rect 5618 102844 5682 102848
rect 5618 102788 5622 102844
rect 5622 102788 5678 102844
rect 5678 102788 5682 102844
rect 5618 102784 5682 102788
rect 5698 102844 5762 102848
rect 5698 102788 5702 102844
rect 5702 102788 5758 102844
rect 5758 102788 5762 102844
rect 5698 102784 5762 102788
rect 5778 102844 5842 102848
rect 5778 102788 5782 102844
rect 5782 102788 5838 102844
rect 5838 102788 5842 102844
rect 5778 102784 5842 102788
rect 5858 102844 5922 102848
rect 5858 102788 5862 102844
rect 5862 102788 5918 102844
rect 5918 102788 5922 102844
rect 5858 102784 5922 102788
rect 10285 102844 10349 102848
rect 10285 102788 10289 102844
rect 10289 102788 10345 102844
rect 10345 102788 10349 102844
rect 10285 102784 10349 102788
rect 10365 102844 10429 102848
rect 10365 102788 10369 102844
rect 10369 102788 10425 102844
rect 10425 102788 10429 102844
rect 10365 102784 10429 102788
rect 10445 102844 10509 102848
rect 10445 102788 10449 102844
rect 10449 102788 10505 102844
rect 10505 102788 10509 102844
rect 10445 102784 10509 102788
rect 10525 102844 10589 102848
rect 10525 102788 10529 102844
rect 10529 102788 10585 102844
rect 10585 102788 10589 102844
rect 10525 102784 10589 102788
rect 3285 102300 3349 102304
rect 3285 102244 3289 102300
rect 3289 102244 3345 102300
rect 3345 102244 3349 102300
rect 3285 102240 3349 102244
rect 3365 102300 3429 102304
rect 3365 102244 3369 102300
rect 3369 102244 3425 102300
rect 3425 102244 3429 102300
rect 3365 102240 3429 102244
rect 3445 102300 3509 102304
rect 3445 102244 3449 102300
rect 3449 102244 3505 102300
rect 3505 102244 3509 102300
rect 3445 102240 3509 102244
rect 3525 102300 3589 102304
rect 3525 102244 3529 102300
rect 3529 102244 3585 102300
rect 3585 102244 3589 102300
rect 3525 102240 3589 102244
rect 7952 102300 8016 102304
rect 7952 102244 7956 102300
rect 7956 102244 8012 102300
rect 8012 102244 8016 102300
rect 7952 102240 8016 102244
rect 8032 102300 8096 102304
rect 8032 102244 8036 102300
rect 8036 102244 8092 102300
rect 8092 102244 8096 102300
rect 8032 102240 8096 102244
rect 8112 102300 8176 102304
rect 8112 102244 8116 102300
rect 8116 102244 8172 102300
rect 8172 102244 8176 102300
rect 8112 102240 8176 102244
rect 8192 102300 8256 102304
rect 8192 102244 8196 102300
rect 8196 102244 8252 102300
rect 8252 102244 8256 102300
rect 8192 102240 8256 102244
rect 5618 101756 5682 101760
rect 5618 101700 5622 101756
rect 5622 101700 5678 101756
rect 5678 101700 5682 101756
rect 5618 101696 5682 101700
rect 5698 101756 5762 101760
rect 5698 101700 5702 101756
rect 5702 101700 5758 101756
rect 5758 101700 5762 101756
rect 5698 101696 5762 101700
rect 5778 101756 5842 101760
rect 5778 101700 5782 101756
rect 5782 101700 5838 101756
rect 5838 101700 5842 101756
rect 5778 101696 5842 101700
rect 5858 101756 5922 101760
rect 5858 101700 5862 101756
rect 5862 101700 5918 101756
rect 5918 101700 5922 101756
rect 5858 101696 5922 101700
rect 10285 101756 10349 101760
rect 10285 101700 10289 101756
rect 10289 101700 10345 101756
rect 10345 101700 10349 101756
rect 10285 101696 10349 101700
rect 10365 101756 10429 101760
rect 10365 101700 10369 101756
rect 10369 101700 10425 101756
rect 10425 101700 10429 101756
rect 10365 101696 10429 101700
rect 10445 101756 10509 101760
rect 10445 101700 10449 101756
rect 10449 101700 10505 101756
rect 10505 101700 10509 101756
rect 10445 101696 10509 101700
rect 10525 101756 10589 101760
rect 10525 101700 10529 101756
rect 10529 101700 10585 101756
rect 10585 101700 10589 101756
rect 10525 101696 10589 101700
rect 3285 101212 3349 101216
rect 3285 101156 3289 101212
rect 3289 101156 3345 101212
rect 3345 101156 3349 101212
rect 3285 101152 3349 101156
rect 3365 101212 3429 101216
rect 3365 101156 3369 101212
rect 3369 101156 3425 101212
rect 3425 101156 3429 101212
rect 3365 101152 3429 101156
rect 3445 101212 3509 101216
rect 3445 101156 3449 101212
rect 3449 101156 3505 101212
rect 3505 101156 3509 101212
rect 3445 101152 3509 101156
rect 3525 101212 3589 101216
rect 3525 101156 3529 101212
rect 3529 101156 3585 101212
rect 3585 101156 3589 101212
rect 3525 101152 3589 101156
rect 7952 101212 8016 101216
rect 7952 101156 7956 101212
rect 7956 101156 8012 101212
rect 8012 101156 8016 101212
rect 7952 101152 8016 101156
rect 8032 101212 8096 101216
rect 8032 101156 8036 101212
rect 8036 101156 8092 101212
rect 8092 101156 8096 101212
rect 8032 101152 8096 101156
rect 8112 101212 8176 101216
rect 8112 101156 8116 101212
rect 8116 101156 8172 101212
rect 8172 101156 8176 101212
rect 8112 101152 8176 101156
rect 8192 101212 8256 101216
rect 8192 101156 8196 101212
rect 8196 101156 8252 101212
rect 8252 101156 8256 101212
rect 8192 101152 8256 101156
rect 5618 100668 5682 100672
rect 5618 100612 5622 100668
rect 5622 100612 5678 100668
rect 5678 100612 5682 100668
rect 5618 100608 5682 100612
rect 5698 100668 5762 100672
rect 5698 100612 5702 100668
rect 5702 100612 5758 100668
rect 5758 100612 5762 100668
rect 5698 100608 5762 100612
rect 5778 100668 5842 100672
rect 5778 100612 5782 100668
rect 5782 100612 5838 100668
rect 5838 100612 5842 100668
rect 5778 100608 5842 100612
rect 5858 100668 5922 100672
rect 5858 100612 5862 100668
rect 5862 100612 5918 100668
rect 5918 100612 5922 100668
rect 5858 100608 5922 100612
rect 10285 100668 10349 100672
rect 10285 100612 10289 100668
rect 10289 100612 10345 100668
rect 10345 100612 10349 100668
rect 10285 100608 10349 100612
rect 10365 100668 10429 100672
rect 10365 100612 10369 100668
rect 10369 100612 10425 100668
rect 10425 100612 10429 100668
rect 10365 100608 10429 100612
rect 10445 100668 10509 100672
rect 10445 100612 10449 100668
rect 10449 100612 10505 100668
rect 10505 100612 10509 100668
rect 10445 100608 10509 100612
rect 10525 100668 10589 100672
rect 10525 100612 10529 100668
rect 10529 100612 10585 100668
rect 10585 100612 10589 100668
rect 10525 100608 10589 100612
rect 3285 100124 3349 100128
rect 3285 100068 3289 100124
rect 3289 100068 3345 100124
rect 3345 100068 3349 100124
rect 3285 100064 3349 100068
rect 3365 100124 3429 100128
rect 3365 100068 3369 100124
rect 3369 100068 3425 100124
rect 3425 100068 3429 100124
rect 3365 100064 3429 100068
rect 3445 100124 3509 100128
rect 3445 100068 3449 100124
rect 3449 100068 3505 100124
rect 3505 100068 3509 100124
rect 3445 100064 3509 100068
rect 3525 100124 3589 100128
rect 3525 100068 3529 100124
rect 3529 100068 3585 100124
rect 3585 100068 3589 100124
rect 3525 100064 3589 100068
rect 7952 100124 8016 100128
rect 7952 100068 7956 100124
rect 7956 100068 8012 100124
rect 8012 100068 8016 100124
rect 7952 100064 8016 100068
rect 8032 100124 8096 100128
rect 8032 100068 8036 100124
rect 8036 100068 8092 100124
rect 8092 100068 8096 100124
rect 8032 100064 8096 100068
rect 8112 100124 8176 100128
rect 8112 100068 8116 100124
rect 8116 100068 8172 100124
rect 8172 100068 8176 100124
rect 8112 100064 8176 100068
rect 8192 100124 8256 100128
rect 8192 100068 8196 100124
rect 8196 100068 8252 100124
rect 8252 100068 8256 100124
rect 8192 100064 8256 100068
rect 5618 99580 5682 99584
rect 5618 99524 5622 99580
rect 5622 99524 5678 99580
rect 5678 99524 5682 99580
rect 5618 99520 5682 99524
rect 5698 99580 5762 99584
rect 5698 99524 5702 99580
rect 5702 99524 5758 99580
rect 5758 99524 5762 99580
rect 5698 99520 5762 99524
rect 5778 99580 5842 99584
rect 5778 99524 5782 99580
rect 5782 99524 5838 99580
rect 5838 99524 5842 99580
rect 5778 99520 5842 99524
rect 5858 99580 5922 99584
rect 5858 99524 5862 99580
rect 5862 99524 5918 99580
rect 5918 99524 5922 99580
rect 5858 99520 5922 99524
rect 10285 99580 10349 99584
rect 10285 99524 10289 99580
rect 10289 99524 10345 99580
rect 10345 99524 10349 99580
rect 10285 99520 10349 99524
rect 10365 99580 10429 99584
rect 10365 99524 10369 99580
rect 10369 99524 10425 99580
rect 10425 99524 10429 99580
rect 10365 99520 10429 99524
rect 10445 99580 10509 99584
rect 10445 99524 10449 99580
rect 10449 99524 10505 99580
rect 10505 99524 10509 99580
rect 10445 99520 10509 99524
rect 10525 99580 10589 99584
rect 10525 99524 10529 99580
rect 10529 99524 10585 99580
rect 10585 99524 10589 99580
rect 10525 99520 10589 99524
rect 3285 99036 3349 99040
rect 3285 98980 3289 99036
rect 3289 98980 3345 99036
rect 3345 98980 3349 99036
rect 3285 98976 3349 98980
rect 3365 99036 3429 99040
rect 3365 98980 3369 99036
rect 3369 98980 3425 99036
rect 3425 98980 3429 99036
rect 3365 98976 3429 98980
rect 3445 99036 3509 99040
rect 3445 98980 3449 99036
rect 3449 98980 3505 99036
rect 3505 98980 3509 99036
rect 3445 98976 3509 98980
rect 3525 99036 3589 99040
rect 3525 98980 3529 99036
rect 3529 98980 3585 99036
rect 3585 98980 3589 99036
rect 3525 98976 3589 98980
rect 7952 99036 8016 99040
rect 7952 98980 7956 99036
rect 7956 98980 8012 99036
rect 8012 98980 8016 99036
rect 7952 98976 8016 98980
rect 8032 99036 8096 99040
rect 8032 98980 8036 99036
rect 8036 98980 8092 99036
rect 8092 98980 8096 99036
rect 8032 98976 8096 98980
rect 8112 99036 8176 99040
rect 8112 98980 8116 99036
rect 8116 98980 8172 99036
rect 8172 98980 8176 99036
rect 8112 98976 8176 98980
rect 8192 99036 8256 99040
rect 8192 98980 8196 99036
rect 8196 98980 8252 99036
rect 8252 98980 8256 99036
rect 8192 98976 8256 98980
rect 5618 98492 5682 98496
rect 5618 98436 5622 98492
rect 5622 98436 5678 98492
rect 5678 98436 5682 98492
rect 5618 98432 5682 98436
rect 5698 98492 5762 98496
rect 5698 98436 5702 98492
rect 5702 98436 5758 98492
rect 5758 98436 5762 98492
rect 5698 98432 5762 98436
rect 5778 98492 5842 98496
rect 5778 98436 5782 98492
rect 5782 98436 5838 98492
rect 5838 98436 5842 98492
rect 5778 98432 5842 98436
rect 5858 98492 5922 98496
rect 5858 98436 5862 98492
rect 5862 98436 5918 98492
rect 5918 98436 5922 98492
rect 5858 98432 5922 98436
rect 10285 98492 10349 98496
rect 10285 98436 10289 98492
rect 10289 98436 10345 98492
rect 10345 98436 10349 98492
rect 10285 98432 10349 98436
rect 10365 98492 10429 98496
rect 10365 98436 10369 98492
rect 10369 98436 10425 98492
rect 10425 98436 10429 98492
rect 10365 98432 10429 98436
rect 10445 98492 10509 98496
rect 10445 98436 10449 98492
rect 10449 98436 10505 98492
rect 10505 98436 10509 98492
rect 10445 98432 10509 98436
rect 10525 98492 10589 98496
rect 10525 98436 10529 98492
rect 10529 98436 10585 98492
rect 10585 98436 10589 98492
rect 10525 98432 10589 98436
rect 3285 97948 3349 97952
rect 3285 97892 3289 97948
rect 3289 97892 3345 97948
rect 3345 97892 3349 97948
rect 3285 97888 3349 97892
rect 3365 97948 3429 97952
rect 3365 97892 3369 97948
rect 3369 97892 3425 97948
rect 3425 97892 3429 97948
rect 3365 97888 3429 97892
rect 3445 97948 3509 97952
rect 3445 97892 3449 97948
rect 3449 97892 3505 97948
rect 3505 97892 3509 97948
rect 3445 97888 3509 97892
rect 3525 97948 3589 97952
rect 3525 97892 3529 97948
rect 3529 97892 3585 97948
rect 3585 97892 3589 97948
rect 3525 97888 3589 97892
rect 7952 97948 8016 97952
rect 7952 97892 7956 97948
rect 7956 97892 8012 97948
rect 8012 97892 8016 97948
rect 7952 97888 8016 97892
rect 8032 97948 8096 97952
rect 8032 97892 8036 97948
rect 8036 97892 8092 97948
rect 8092 97892 8096 97948
rect 8032 97888 8096 97892
rect 8112 97948 8176 97952
rect 8112 97892 8116 97948
rect 8116 97892 8172 97948
rect 8172 97892 8176 97948
rect 8112 97888 8176 97892
rect 8192 97948 8256 97952
rect 8192 97892 8196 97948
rect 8196 97892 8252 97948
rect 8252 97892 8256 97948
rect 8192 97888 8256 97892
rect 5618 97404 5682 97408
rect 5618 97348 5622 97404
rect 5622 97348 5678 97404
rect 5678 97348 5682 97404
rect 5618 97344 5682 97348
rect 5698 97404 5762 97408
rect 5698 97348 5702 97404
rect 5702 97348 5758 97404
rect 5758 97348 5762 97404
rect 5698 97344 5762 97348
rect 5778 97404 5842 97408
rect 5778 97348 5782 97404
rect 5782 97348 5838 97404
rect 5838 97348 5842 97404
rect 5778 97344 5842 97348
rect 5858 97404 5922 97408
rect 5858 97348 5862 97404
rect 5862 97348 5918 97404
rect 5918 97348 5922 97404
rect 5858 97344 5922 97348
rect 10285 97404 10349 97408
rect 10285 97348 10289 97404
rect 10289 97348 10345 97404
rect 10345 97348 10349 97404
rect 10285 97344 10349 97348
rect 10365 97404 10429 97408
rect 10365 97348 10369 97404
rect 10369 97348 10425 97404
rect 10425 97348 10429 97404
rect 10365 97344 10429 97348
rect 10445 97404 10509 97408
rect 10445 97348 10449 97404
rect 10449 97348 10505 97404
rect 10505 97348 10509 97404
rect 10445 97344 10509 97348
rect 10525 97404 10589 97408
rect 10525 97348 10529 97404
rect 10529 97348 10585 97404
rect 10585 97348 10589 97404
rect 10525 97344 10589 97348
rect 3285 96860 3349 96864
rect 3285 96804 3289 96860
rect 3289 96804 3345 96860
rect 3345 96804 3349 96860
rect 3285 96800 3349 96804
rect 3365 96860 3429 96864
rect 3365 96804 3369 96860
rect 3369 96804 3425 96860
rect 3425 96804 3429 96860
rect 3365 96800 3429 96804
rect 3445 96860 3509 96864
rect 3445 96804 3449 96860
rect 3449 96804 3505 96860
rect 3505 96804 3509 96860
rect 3445 96800 3509 96804
rect 3525 96860 3589 96864
rect 3525 96804 3529 96860
rect 3529 96804 3585 96860
rect 3585 96804 3589 96860
rect 3525 96800 3589 96804
rect 7952 96860 8016 96864
rect 7952 96804 7956 96860
rect 7956 96804 8012 96860
rect 8012 96804 8016 96860
rect 7952 96800 8016 96804
rect 8032 96860 8096 96864
rect 8032 96804 8036 96860
rect 8036 96804 8092 96860
rect 8092 96804 8096 96860
rect 8032 96800 8096 96804
rect 8112 96860 8176 96864
rect 8112 96804 8116 96860
rect 8116 96804 8172 96860
rect 8172 96804 8176 96860
rect 8112 96800 8176 96804
rect 8192 96860 8256 96864
rect 8192 96804 8196 96860
rect 8196 96804 8252 96860
rect 8252 96804 8256 96860
rect 8192 96800 8256 96804
rect 5618 96316 5682 96320
rect 5618 96260 5622 96316
rect 5622 96260 5678 96316
rect 5678 96260 5682 96316
rect 5618 96256 5682 96260
rect 5698 96316 5762 96320
rect 5698 96260 5702 96316
rect 5702 96260 5758 96316
rect 5758 96260 5762 96316
rect 5698 96256 5762 96260
rect 5778 96316 5842 96320
rect 5778 96260 5782 96316
rect 5782 96260 5838 96316
rect 5838 96260 5842 96316
rect 5778 96256 5842 96260
rect 5858 96316 5922 96320
rect 5858 96260 5862 96316
rect 5862 96260 5918 96316
rect 5918 96260 5922 96316
rect 5858 96256 5922 96260
rect 10285 96316 10349 96320
rect 10285 96260 10289 96316
rect 10289 96260 10345 96316
rect 10345 96260 10349 96316
rect 10285 96256 10349 96260
rect 10365 96316 10429 96320
rect 10365 96260 10369 96316
rect 10369 96260 10425 96316
rect 10425 96260 10429 96316
rect 10365 96256 10429 96260
rect 10445 96316 10509 96320
rect 10445 96260 10449 96316
rect 10449 96260 10505 96316
rect 10505 96260 10509 96316
rect 10445 96256 10509 96260
rect 10525 96316 10589 96320
rect 10525 96260 10529 96316
rect 10529 96260 10585 96316
rect 10585 96260 10589 96316
rect 10525 96256 10589 96260
rect 3285 95772 3349 95776
rect 3285 95716 3289 95772
rect 3289 95716 3345 95772
rect 3345 95716 3349 95772
rect 3285 95712 3349 95716
rect 3365 95772 3429 95776
rect 3365 95716 3369 95772
rect 3369 95716 3425 95772
rect 3425 95716 3429 95772
rect 3365 95712 3429 95716
rect 3445 95772 3509 95776
rect 3445 95716 3449 95772
rect 3449 95716 3505 95772
rect 3505 95716 3509 95772
rect 3445 95712 3509 95716
rect 3525 95772 3589 95776
rect 3525 95716 3529 95772
rect 3529 95716 3585 95772
rect 3585 95716 3589 95772
rect 3525 95712 3589 95716
rect 7952 95772 8016 95776
rect 7952 95716 7956 95772
rect 7956 95716 8012 95772
rect 8012 95716 8016 95772
rect 7952 95712 8016 95716
rect 8032 95772 8096 95776
rect 8032 95716 8036 95772
rect 8036 95716 8092 95772
rect 8092 95716 8096 95772
rect 8032 95712 8096 95716
rect 8112 95772 8176 95776
rect 8112 95716 8116 95772
rect 8116 95716 8172 95772
rect 8172 95716 8176 95772
rect 8112 95712 8176 95716
rect 8192 95772 8256 95776
rect 8192 95716 8196 95772
rect 8196 95716 8252 95772
rect 8252 95716 8256 95772
rect 8192 95712 8256 95716
rect 5618 95228 5682 95232
rect 5618 95172 5622 95228
rect 5622 95172 5678 95228
rect 5678 95172 5682 95228
rect 5618 95168 5682 95172
rect 5698 95228 5762 95232
rect 5698 95172 5702 95228
rect 5702 95172 5758 95228
rect 5758 95172 5762 95228
rect 5698 95168 5762 95172
rect 5778 95228 5842 95232
rect 5778 95172 5782 95228
rect 5782 95172 5838 95228
rect 5838 95172 5842 95228
rect 5778 95168 5842 95172
rect 5858 95228 5922 95232
rect 5858 95172 5862 95228
rect 5862 95172 5918 95228
rect 5918 95172 5922 95228
rect 5858 95168 5922 95172
rect 10285 95228 10349 95232
rect 10285 95172 10289 95228
rect 10289 95172 10345 95228
rect 10345 95172 10349 95228
rect 10285 95168 10349 95172
rect 10365 95228 10429 95232
rect 10365 95172 10369 95228
rect 10369 95172 10425 95228
rect 10425 95172 10429 95228
rect 10365 95168 10429 95172
rect 10445 95228 10509 95232
rect 10445 95172 10449 95228
rect 10449 95172 10505 95228
rect 10505 95172 10509 95228
rect 10445 95168 10509 95172
rect 10525 95228 10589 95232
rect 10525 95172 10529 95228
rect 10529 95172 10585 95228
rect 10585 95172 10589 95228
rect 10525 95168 10589 95172
rect 3285 94684 3349 94688
rect 3285 94628 3289 94684
rect 3289 94628 3345 94684
rect 3345 94628 3349 94684
rect 3285 94624 3349 94628
rect 3365 94684 3429 94688
rect 3365 94628 3369 94684
rect 3369 94628 3425 94684
rect 3425 94628 3429 94684
rect 3365 94624 3429 94628
rect 3445 94684 3509 94688
rect 3445 94628 3449 94684
rect 3449 94628 3505 94684
rect 3505 94628 3509 94684
rect 3445 94624 3509 94628
rect 3525 94684 3589 94688
rect 3525 94628 3529 94684
rect 3529 94628 3585 94684
rect 3585 94628 3589 94684
rect 3525 94624 3589 94628
rect 7952 94684 8016 94688
rect 7952 94628 7956 94684
rect 7956 94628 8012 94684
rect 8012 94628 8016 94684
rect 7952 94624 8016 94628
rect 8032 94684 8096 94688
rect 8032 94628 8036 94684
rect 8036 94628 8092 94684
rect 8092 94628 8096 94684
rect 8032 94624 8096 94628
rect 8112 94684 8176 94688
rect 8112 94628 8116 94684
rect 8116 94628 8172 94684
rect 8172 94628 8176 94684
rect 8112 94624 8176 94628
rect 8192 94684 8256 94688
rect 8192 94628 8196 94684
rect 8196 94628 8252 94684
rect 8252 94628 8256 94684
rect 8192 94624 8256 94628
rect 5618 94140 5682 94144
rect 5618 94084 5622 94140
rect 5622 94084 5678 94140
rect 5678 94084 5682 94140
rect 5618 94080 5682 94084
rect 5698 94140 5762 94144
rect 5698 94084 5702 94140
rect 5702 94084 5758 94140
rect 5758 94084 5762 94140
rect 5698 94080 5762 94084
rect 5778 94140 5842 94144
rect 5778 94084 5782 94140
rect 5782 94084 5838 94140
rect 5838 94084 5842 94140
rect 5778 94080 5842 94084
rect 5858 94140 5922 94144
rect 5858 94084 5862 94140
rect 5862 94084 5918 94140
rect 5918 94084 5922 94140
rect 5858 94080 5922 94084
rect 10285 94140 10349 94144
rect 10285 94084 10289 94140
rect 10289 94084 10345 94140
rect 10345 94084 10349 94140
rect 10285 94080 10349 94084
rect 10365 94140 10429 94144
rect 10365 94084 10369 94140
rect 10369 94084 10425 94140
rect 10425 94084 10429 94140
rect 10365 94080 10429 94084
rect 10445 94140 10509 94144
rect 10445 94084 10449 94140
rect 10449 94084 10505 94140
rect 10505 94084 10509 94140
rect 10445 94080 10509 94084
rect 10525 94140 10589 94144
rect 10525 94084 10529 94140
rect 10529 94084 10585 94140
rect 10585 94084 10589 94140
rect 10525 94080 10589 94084
rect 3285 93596 3349 93600
rect 3285 93540 3289 93596
rect 3289 93540 3345 93596
rect 3345 93540 3349 93596
rect 3285 93536 3349 93540
rect 3365 93596 3429 93600
rect 3365 93540 3369 93596
rect 3369 93540 3425 93596
rect 3425 93540 3429 93596
rect 3365 93536 3429 93540
rect 3445 93596 3509 93600
rect 3445 93540 3449 93596
rect 3449 93540 3505 93596
rect 3505 93540 3509 93596
rect 3445 93536 3509 93540
rect 3525 93596 3589 93600
rect 3525 93540 3529 93596
rect 3529 93540 3585 93596
rect 3585 93540 3589 93596
rect 3525 93536 3589 93540
rect 7952 93596 8016 93600
rect 7952 93540 7956 93596
rect 7956 93540 8012 93596
rect 8012 93540 8016 93596
rect 7952 93536 8016 93540
rect 8032 93596 8096 93600
rect 8032 93540 8036 93596
rect 8036 93540 8092 93596
rect 8092 93540 8096 93596
rect 8032 93536 8096 93540
rect 8112 93596 8176 93600
rect 8112 93540 8116 93596
rect 8116 93540 8172 93596
rect 8172 93540 8176 93596
rect 8112 93536 8176 93540
rect 8192 93596 8256 93600
rect 8192 93540 8196 93596
rect 8196 93540 8252 93596
rect 8252 93540 8256 93596
rect 8192 93536 8256 93540
rect 5618 93052 5682 93056
rect 5618 92996 5622 93052
rect 5622 92996 5678 93052
rect 5678 92996 5682 93052
rect 5618 92992 5682 92996
rect 5698 93052 5762 93056
rect 5698 92996 5702 93052
rect 5702 92996 5758 93052
rect 5758 92996 5762 93052
rect 5698 92992 5762 92996
rect 5778 93052 5842 93056
rect 5778 92996 5782 93052
rect 5782 92996 5838 93052
rect 5838 92996 5842 93052
rect 5778 92992 5842 92996
rect 5858 93052 5922 93056
rect 5858 92996 5862 93052
rect 5862 92996 5918 93052
rect 5918 92996 5922 93052
rect 5858 92992 5922 92996
rect 10285 93052 10349 93056
rect 10285 92996 10289 93052
rect 10289 92996 10345 93052
rect 10345 92996 10349 93052
rect 10285 92992 10349 92996
rect 10365 93052 10429 93056
rect 10365 92996 10369 93052
rect 10369 92996 10425 93052
rect 10425 92996 10429 93052
rect 10365 92992 10429 92996
rect 10445 93052 10509 93056
rect 10445 92996 10449 93052
rect 10449 92996 10505 93052
rect 10505 92996 10509 93052
rect 10445 92992 10509 92996
rect 10525 93052 10589 93056
rect 10525 92996 10529 93052
rect 10529 92996 10585 93052
rect 10585 92996 10589 93052
rect 10525 92992 10589 92996
rect 3285 92508 3349 92512
rect 3285 92452 3289 92508
rect 3289 92452 3345 92508
rect 3345 92452 3349 92508
rect 3285 92448 3349 92452
rect 3365 92508 3429 92512
rect 3365 92452 3369 92508
rect 3369 92452 3425 92508
rect 3425 92452 3429 92508
rect 3365 92448 3429 92452
rect 3445 92508 3509 92512
rect 3445 92452 3449 92508
rect 3449 92452 3505 92508
rect 3505 92452 3509 92508
rect 3445 92448 3509 92452
rect 3525 92508 3589 92512
rect 3525 92452 3529 92508
rect 3529 92452 3585 92508
rect 3585 92452 3589 92508
rect 3525 92448 3589 92452
rect 7952 92508 8016 92512
rect 7952 92452 7956 92508
rect 7956 92452 8012 92508
rect 8012 92452 8016 92508
rect 7952 92448 8016 92452
rect 8032 92508 8096 92512
rect 8032 92452 8036 92508
rect 8036 92452 8092 92508
rect 8092 92452 8096 92508
rect 8032 92448 8096 92452
rect 8112 92508 8176 92512
rect 8112 92452 8116 92508
rect 8116 92452 8172 92508
rect 8172 92452 8176 92508
rect 8112 92448 8176 92452
rect 8192 92508 8256 92512
rect 8192 92452 8196 92508
rect 8196 92452 8252 92508
rect 8252 92452 8256 92508
rect 8192 92448 8256 92452
rect 5618 91964 5682 91968
rect 5618 91908 5622 91964
rect 5622 91908 5678 91964
rect 5678 91908 5682 91964
rect 5618 91904 5682 91908
rect 5698 91964 5762 91968
rect 5698 91908 5702 91964
rect 5702 91908 5758 91964
rect 5758 91908 5762 91964
rect 5698 91904 5762 91908
rect 5778 91964 5842 91968
rect 5778 91908 5782 91964
rect 5782 91908 5838 91964
rect 5838 91908 5842 91964
rect 5778 91904 5842 91908
rect 5858 91964 5922 91968
rect 5858 91908 5862 91964
rect 5862 91908 5918 91964
rect 5918 91908 5922 91964
rect 5858 91904 5922 91908
rect 10285 91964 10349 91968
rect 10285 91908 10289 91964
rect 10289 91908 10345 91964
rect 10345 91908 10349 91964
rect 10285 91904 10349 91908
rect 10365 91964 10429 91968
rect 10365 91908 10369 91964
rect 10369 91908 10425 91964
rect 10425 91908 10429 91964
rect 10365 91904 10429 91908
rect 10445 91964 10509 91968
rect 10445 91908 10449 91964
rect 10449 91908 10505 91964
rect 10505 91908 10509 91964
rect 10445 91904 10509 91908
rect 10525 91964 10589 91968
rect 10525 91908 10529 91964
rect 10529 91908 10585 91964
rect 10585 91908 10589 91964
rect 10525 91904 10589 91908
rect 3285 91420 3349 91424
rect 3285 91364 3289 91420
rect 3289 91364 3345 91420
rect 3345 91364 3349 91420
rect 3285 91360 3349 91364
rect 3365 91420 3429 91424
rect 3365 91364 3369 91420
rect 3369 91364 3425 91420
rect 3425 91364 3429 91420
rect 3365 91360 3429 91364
rect 3445 91420 3509 91424
rect 3445 91364 3449 91420
rect 3449 91364 3505 91420
rect 3505 91364 3509 91420
rect 3445 91360 3509 91364
rect 3525 91420 3589 91424
rect 3525 91364 3529 91420
rect 3529 91364 3585 91420
rect 3585 91364 3589 91420
rect 3525 91360 3589 91364
rect 7952 91420 8016 91424
rect 7952 91364 7956 91420
rect 7956 91364 8012 91420
rect 8012 91364 8016 91420
rect 7952 91360 8016 91364
rect 8032 91420 8096 91424
rect 8032 91364 8036 91420
rect 8036 91364 8092 91420
rect 8092 91364 8096 91420
rect 8032 91360 8096 91364
rect 8112 91420 8176 91424
rect 8112 91364 8116 91420
rect 8116 91364 8172 91420
rect 8172 91364 8176 91420
rect 8112 91360 8176 91364
rect 8192 91420 8256 91424
rect 8192 91364 8196 91420
rect 8196 91364 8252 91420
rect 8252 91364 8256 91420
rect 8192 91360 8256 91364
rect 5618 90876 5682 90880
rect 5618 90820 5622 90876
rect 5622 90820 5678 90876
rect 5678 90820 5682 90876
rect 5618 90816 5682 90820
rect 5698 90876 5762 90880
rect 5698 90820 5702 90876
rect 5702 90820 5758 90876
rect 5758 90820 5762 90876
rect 5698 90816 5762 90820
rect 5778 90876 5842 90880
rect 5778 90820 5782 90876
rect 5782 90820 5838 90876
rect 5838 90820 5842 90876
rect 5778 90816 5842 90820
rect 5858 90876 5922 90880
rect 5858 90820 5862 90876
rect 5862 90820 5918 90876
rect 5918 90820 5922 90876
rect 5858 90816 5922 90820
rect 10285 90876 10349 90880
rect 10285 90820 10289 90876
rect 10289 90820 10345 90876
rect 10345 90820 10349 90876
rect 10285 90816 10349 90820
rect 10365 90876 10429 90880
rect 10365 90820 10369 90876
rect 10369 90820 10425 90876
rect 10425 90820 10429 90876
rect 10365 90816 10429 90820
rect 10445 90876 10509 90880
rect 10445 90820 10449 90876
rect 10449 90820 10505 90876
rect 10505 90820 10509 90876
rect 10445 90816 10509 90820
rect 10525 90876 10589 90880
rect 10525 90820 10529 90876
rect 10529 90820 10585 90876
rect 10585 90820 10589 90876
rect 10525 90816 10589 90820
rect 3285 90332 3349 90336
rect 3285 90276 3289 90332
rect 3289 90276 3345 90332
rect 3345 90276 3349 90332
rect 3285 90272 3349 90276
rect 3365 90332 3429 90336
rect 3365 90276 3369 90332
rect 3369 90276 3425 90332
rect 3425 90276 3429 90332
rect 3365 90272 3429 90276
rect 3445 90332 3509 90336
rect 3445 90276 3449 90332
rect 3449 90276 3505 90332
rect 3505 90276 3509 90332
rect 3445 90272 3509 90276
rect 3525 90332 3589 90336
rect 3525 90276 3529 90332
rect 3529 90276 3585 90332
rect 3585 90276 3589 90332
rect 3525 90272 3589 90276
rect 7952 90332 8016 90336
rect 7952 90276 7956 90332
rect 7956 90276 8012 90332
rect 8012 90276 8016 90332
rect 7952 90272 8016 90276
rect 8032 90332 8096 90336
rect 8032 90276 8036 90332
rect 8036 90276 8092 90332
rect 8092 90276 8096 90332
rect 8032 90272 8096 90276
rect 8112 90332 8176 90336
rect 8112 90276 8116 90332
rect 8116 90276 8172 90332
rect 8172 90276 8176 90332
rect 8112 90272 8176 90276
rect 8192 90332 8256 90336
rect 8192 90276 8196 90332
rect 8196 90276 8252 90332
rect 8252 90276 8256 90332
rect 8192 90272 8256 90276
rect 5618 89788 5682 89792
rect 5618 89732 5622 89788
rect 5622 89732 5678 89788
rect 5678 89732 5682 89788
rect 5618 89728 5682 89732
rect 5698 89788 5762 89792
rect 5698 89732 5702 89788
rect 5702 89732 5758 89788
rect 5758 89732 5762 89788
rect 5698 89728 5762 89732
rect 5778 89788 5842 89792
rect 5778 89732 5782 89788
rect 5782 89732 5838 89788
rect 5838 89732 5842 89788
rect 5778 89728 5842 89732
rect 5858 89788 5922 89792
rect 5858 89732 5862 89788
rect 5862 89732 5918 89788
rect 5918 89732 5922 89788
rect 5858 89728 5922 89732
rect 10285 89788 10349 89792
rect 10285 89732 10289 89788
rect 10289 89732 10345 89788
rect 10345 89732 10349 89788
rect 10285 89728 10349 89732
rect 10365 89788 10429 89792
rect 10365 89732 10369 89788
rect 10369 89732 10425 89788
rect 10425 89732 10429 89788
rect 10365 89728 10429 89732
rect 10445 89788 10509 89792
rect 10445 89732 10449 89788
rect 10449 89732 10505 89788
rect 10505 89732 10509 89788
rect 10445 89728 10509 89732
rect 10525 89788 10589 89792
rect 10525 89732 10529 89788
rect 10529 89732 10585 89788
rect 10585 89732 10589 89788
rect 10525 89728 10589 89732
rect 3285 89244 3349 89248
rect 3285 89188 3289 89244
rect 3289 89188 3345 89244
rect 3345 89188 3349 89244
rect 3285 89184 3349 89188
rect 3365 89244 3429 89248
rect 3365 89188 3369 89244
rect 3369 89188 3425 89244
rect 3425 89188 3429 89244
rect 3365 89184 3429 89188
rect 3445 89244 3509 89248
rect 3445 89188 3449 89244
rect 3449 89188 3505 89244
rect 3505 89188 3509 89244
rect 3445 89184 3509 89188
rect 3525 89244 3589 89248
rect 3525 89188 3529 89244
rect 3529 89188 3585 89244
rect 3585 89188 3589 89244
rect 3525 89184 3589 89188
rect 7952 89244 8016 89248
rect 7952 89188 7956 89244
rect 7956 89188 8012 89244
rect 8012 89188 8016 89244
rect 7952 89184 8016 89188
rect 8032 89244 8096 89248
rect 8032 89188 8036 89244
rect 8036 89188 8092 89244
rect 8092 89188 8096 89244
rect 8032 89184 8096 89188
rect 8112 89244 8176 89248
rect 8112 89188 8116 89244
rect 8116 89188 8172 89244
rect 8172 89188 8176 89244
rect 8112 89184 8176 89188
rect 8192 89244 8256 89248
rect 8192 89188 8196 89244
rect 8196 89188 8252 89244
rect 8252 89188 8256 89244
rect 8192 89184 8256 89188
rect 5618 88700 5682 88704
rect 5618 88644 5622 88700
rect 5622 88644 5678 88700
rect 5678 88644 5682 88700
rect 5618 88640 5682 88644
rect 5698 88700 5762 88704
rect 5698 88644 5702 88700
rect 5702 88644 5758 88700
rect 5758 88644 5762 88700
rect 5698 88640 5762 88644
rect 5778 88700 5842 88704
rect 5778 88644 5782 88700
rect 5782 88644 5838 88700
rect 5838 88644 5842 88700
rect 5778 88640 5842 88644
rect 5858 88700 5922 88704
rect 5858 88644 5862 88700
rect 5862 88644 5918 88700
rect 5918 88644 5922 88700
rect 5858 88640 5922 88644
rect 10285 88700 10349 88704
rect 10285 88644 10289 88700
rect 10289 88644 10345 88700
rect 10345 88644 10349 88700
rect 10285 88640 10349 88644
rect 10365 88700 10429 88704
rect 10365 88644 10369 88700
rect 10369 88644 10425 88700
rect 10425 88644 10429 88700
rect 10365 88640 10429 88644
rect 10445 88700 10509 88704
rect 10445 88644 10449 88700
rect 10449 88644 10505 88700
rect 10505 88644 10509 88700
rect 10445 88640 10509 88644
rect 10525 88700 10589 88704
rect 10525 88644 10529 88700
rect 10529 88644 10585 88700
rect 10585 88644 10589 88700
rect 10525 88640 10589 88644
rect 3285 88156 3349 88160
rect 3285 88100 3289 88156
rect 3289 88100 3345 88156
rect 3345 88100 3349 88156
rect 3285 88096 3349 88100
rect 3365 88156 3429 88160
rect 3365 88100 3369 88156
rect 3369 88100 3425 88156
rect 3425 88100 3429 88156
rect 3365 88096 3429 88100
rect 3445 88156 3509 88160
rect 3445 88100 3449 88156
rect 3449 88100 3505 88156
rect 3505 88100 3509 88156
rect 3445 88096 3509 88100
rect 3525 88156 3589 88160
rect 3525 88100 3529 88156
rect 3529 88100 3585 88156
rect 3585 88100 3589 88156
rect 3525 88096 3589 88100
rect 7952 88156 8016 88160
rect 7952 88100 7956 88156
rect 7956 88100 8012 88156
rect 8012 88100 8016 88156
rect 7952 88096 8016 88100
rect 8032 88156 8096 88160
rect 8032 88100 8036 88156
rect 8036 88100 8092 88156
rect 8092 88100 8096 88156
rect 8032 88096 8096 88100
rect 8112 88156 8176 88160
rect 8112 88100 8116 88156
rect 8116 88100 8172 88156
rect 8172 88100 8176 88156
rect 8112 88096 8176 88100
rect 8192 88156 8256 88160
rect 8192 88100 8196 88156
rect 8196 88100 8252 88156
rect 8252 88100 8256 88156
rect 8192 88096 8256 88100
rect 5618 87612 5682 87616
rect 5618 87556 5622 87612
rect 5622 87556 5678 87612
rect 5678 87556 5682 87612
rect 5618 87552 5682 87556
rect 5698 87612 5762 87616
rect 5698 87556 5702 87612
rect 5702 87556 5758 87612
rect 5758 87556 5762 87612
rect 5698 87552 5762 87556
rect 5778 87612 5842 87616
rect 5778 87556 5782 87612
rect 5782 87556 5838 87612
rect 5838 87556 5842 87612
rect 5778 87552 5842 87556
rect 5858 87612 5922 87616
rect 5858 87556 5862 87612
rect 5862 87556 5918 87612
rect 5918 87556 5922 87612
rect 5858 87552 5922 87556
rect 10285 87612 10349 87616
rect 10285 87556 10289 87612
rect 10289 87556 10345 87612
rect 10345 87556 10349 87612
rect 10285 87552 10349 87556
rect 10365 87612 10429 87616
rect 10365 87556 10369 87612
rect 10369 87556 10425 87612
rect 10425 87556 10429 87612
rect 10365 87552 10429 87556
rect 10445 87612 10509 87616
rect 10445 87556 10449 87612
rect 10449 87556 10505 87612
rect 10505 87556 10509 87612
rect 10445 87552 10509 87556
rect 10525 87612 10589 87616
rect 10525 87556 10529 87612
rect 10529 87556 10585 87612
rect 10585 87556 10589 87612
rect 10525 87552 10589 87556
rect 3285 87068 3349 87072
rect 3285 87012 3289 87068
rect 3289 87012 3345 87068
rect 3345 87012 3349 87068
rect 3285 87008 3349 87012
rect 3365 87068 3429 87072
rect 3365 87012 3369 87068
rect 3369 87012 3425 87068
rect 3425 87012 3429 87068
rect 3365 87008 3429 87012
rect 3445 87068 3509 87072
rect 3445 87012 3449 87068
rect 3449 87012 3505 87068
rect 3505 87012 3509 87068
rect 3445 87008 3509 87012
rect 3525 87068 3589 87072
rect 3525 87012 3529 87068
rect 3529 87012 3585 87068
rect 3585 87012 3589 87068
rect 3525 87008 3589 87012
rect 7952 87068 8016 87072
rect 7952 87012 7956 87068
rect 7956 87012 8012 87068
rect 8012 87012 8016 87068
rect 7952 87008 8016 87012
rect 8032 87068 8096 87072
rect 8032 87012 8036 87068
rect 8036 87012 8092 87068
rect 8092 87012 8096 87068
rect 8032 87008 8096 87012
rect 8112 87068 8176 87072
rect 8112 87012 8116 87068
rect 8116 87012 8172 87068
rect 8172 87012 8176 87068
rect 8112 87008 8176 87012
rect 8192 87068 8256 87072
rect 8192 87012 8196 87068
rect 8196 87012 8252 87068
rect 8252 87012 8256 87068
rect 8192 87008 8256 87012
rect 5618 86524 5682 86528
rect 5618 86468 5622 86524
rect 5622 86468 5678 86524
rect 5678 86468 5682 86524
rect 5618 86464 5682 86468
rect 5698 86524 5762 86528
rect 5698 86468 5702 86524
rect 5702 86468 5758 86524
rect 5758 86468 5762 86524
rect 5698 86464 5762 86468
rect 5778 86524 5842 86528
rect 5778 86468 5782 86524
rect 5782 86468 5838 86524
rect 5838 86468 5842 86524
rect 5778 86464 5842 86468
rect 5858 86524 5922 86528
rect 5858 86468 5862 86524
rect 5862 86468 5918 86524
rect 5918 86468 5922 86524
rect 5858 86464 5922 86468
rect 10285 86524 10349 86528
rect 10285 86468 10289 86524
rect 10289 86468 10345 86524
rect 10345 86468 10349 86524
rect 10285 86464 10349 86468
rect 10365 86524 10429 86528
rect 10365 86468 10369 86524
rect 10369 86468 10425 86524
rect 10425 86468 10429 86524
rect 10365 86464 10429 86468
rect 10445 86524 10509 86528
rect 10445 86468 10449 86524
rect 10449 86468 10505 86524
rect 10505 86468 10509 86524
rect 10445 86464 10509 86468
rect 10525 86524 10589 86528
rect 10525 86468 10529 86524
rect 10529 86468 10585 86524
rect 10585 86468 10589 86524
rect 10525 86464 10589 86468
rect 3285 85980 3349 85984
rect 3285 85924 3289 85980
rect 3289 85924 3345 85980
rect 3345 85924 3349 85980
rect 3285 85920 3349 85924
rect 3365 85980 3429 85984
rect 3365 85924 3369 85980
rect 3369 85924 3425 85980
rect 3425 85924 3429 85980
rect 3365 85920 3429 85924
rect 3445 85980 3509 85984
rect 3445 85924 3449 85980
rect 3449 85924 3505 85980
rect 3505 85924 3509 85980
rect 3445 85920 3509 85924
rect 3525 85980 3589 85984
rect 3525 85924 3529 85980
rect 3529 85924 3585 85980
rect 3585 85924 3589 85980
rect 3525 85920 3589 85924
rect 7952 85980 8016 85984
rect 7952 85924 7956 85980
rect 7956 85924 8012 85980
rect 8012 85924 8016 85980
rect 7952 85920 8016 85924
rect 8032 85980 8096 85984
rect 8032 85924 8036 85980
rect 8036 85924 8092 85980
rect 8092 85924 8096 85980
rect 8032 85920 8096 85924
rect 8112 85980 8176 85984
rect 8112 85924 8116 85980
rect 8116 85924 8172 85980
rect 8172 85924 8176 85980
rect 8112 85920 8176 85924
rect 8192 85980 8256 85984
rect 8192 85924 8196 85980
rect 8196 85924 8252 85980
rect 8252 85924 8256 85980
rect 8192 85920 8256 85924
rect 5618 85436 5682 85440
rect 5618 85380 5622 85436
rect 5622 85380 5678 85436
rect 5678 85380 5682 85436
rect 5618 85376 5682 85380
rect 5698 85436 5762 85440
rect 5698 85380 5702 85436
rect 5702 85380 5758 85436
rect 5758 85380 5762 85436
rect 5698 85376 5762 85380
rect 5778 85436 5842 85440
rect 5778 85380 5782 85436
rect 5782 85380 5838 85436
rect 5838 85380 5842 85436
rect 5778 85376 5842 85380
rect 5858 85436 5922 85440
rect 5858 85380 5862 85436
rect 5862 85380 5918 85436
rect 5918 85380 5922 85436
rect 5858 85376 5922 85380
rect 10285 85436 10349 85440
rect 10285 85380 10289 85436
rect 10289 85380 10345 85436
rect 10345 85380 10349 85436
rect 10285 85376 10349 85380
rect 10365 85436 10429 85440
rect 10365 85380 10369 85436
rect 10369 85380 10425 85436
rect 10425 85380 10429 85436
rect 10365 85376 10429 85380
rect 10445 85436 10509 85440
rect 10445 85380 10449 85436
rect 10449 85380 10505 85436
rect 10505 85380 10509 85436
rect 10445 85376 10509 85380
rect 10525 85436 10589 85440
rect 10525 85380 10529 85436
rect 10529 85380 10585 85436
rect 10585 85380 10589 85436
rect 10525 85376 10589 85380
rect 3285 84892 3349 84896
rect 3285 84836 3289 84892
rect 3289 84836 3345 84892
rect 3345 84836 3349 84892
rect 3285 84832 3349 84836
rect 3365 84892 3429 84896
rect 3365 84836 3369 84892
rect 3369 84836 3425 84892
rect 3425 84836 3429 84892
rect 3365 84832 3429 84836
rect 3445 84892 3509 84896
rect 3445 84836 3449 84892
rect 3449 84836 3505 84892
rect 3505 84836 3509 84892
rect 3445 84832 3509 84836
rect 3525 84892 3589 84896
rect 3525 84836 3529 84892
rect 3529 84836 3585 84892
rect 3585 84836 3589 84892
rect 3525 84832 3589 84836
rect 7952 84892 8016 84896
rect 7952 84836 7956 84892
rect 7956 84836 8012 84892
rect 8012 84836 8016 84892
rect 7952 84832 8016 84836
rect 8032 84892 8096 84896
rect 8032 84836 8036 84892
rect 8036 84836 8092 84892
rect 8092 84836 8096 84892
rect 8032 84832 8096 84836
rect 8112 84892 8176 84896
rect 8112 84836 8116 84892
rect 8116 84836 8172 84892
rect 8172 84836 8176 84892
rect 8112 84832 8176 84836
rect 8192 84892 8256 84896
rect 8192 84836 8196 84892
rect 8196 84836 8252 84892
rect 8252 84836 8256 84892
rect 8192 84832 8256 84836
rect 5618 84348 5682 84352
rect 5618 84292 5622 84348
rect 5622 84292 5678 84348
rect 5678 84292 5682 84348
rect 5618 84288 5682 84292
rect 5698 84348 5762 84352
rect 5698 84292 5702 84348
rect 5702 84292 5758 84348
rect 5758 84292 5762 84348
rect 5698 84288 5762 84292
rect 5778 84348 5842 84352
rect 5778 84292 5782 84348
rect 5782 84292 5838 84348
rect 5838 84292 5842 84348
rect 5778 84288 5842 84292
rect 5858 84348 5922 84352
rect 5858 84292 5862 84348
rect 5862 84292 5918 84348
rect 5918 84292 5922 84348
rect 5858 84288 5922 84292
rect 10285 84348 10349 84352
rect 10285 84292 10289 84348
rect 10289 84292 10345 84348
rect 10345 84292 10349 84348
rect 10285 84288 10349 84292
rect 10365 84348 10429 84352
rect 10365 84292 10369 84348
rect 10369 84292 10425 84348
rect 10425 84292 10429 84348
rect 10365 84288 10429 84292
rect 10445 84348 10509 84352
rect 10445 84292 10449 84348
rect 10449 84292 10505 84348
rect 10505 84292 10509 84348
rect 10445 84288 10509 84292
rect 10525 84348 10589 84352
rect 10525 84292 10529 84348
rect 10529 84292 10585 84348
rect 10585 84292 10589 84348
rect 10525 84288 10589 84292
rect 3285 83804 3349 83808
rect 3285 83748 3289 83804
rect 3289 83748 3345 83804
rect 3345 83748 3349 83804
rect 3285 83744 3349 83748
rect 3365 83804 3429 83808
rect 3365 83748 3369 83804
rect 3369 83748 3425 83804
rect 3425 83748 3429 83804
rect 3365 83744 3429 83748
rect 3445 83804 3509 83808
rect 3445 83748 3449 83804
rect 3449 83748 3505 83804
rect 3505 83748 3509 83804
rect 3445 83744 3509 83748
rect 3525 83804 3589 83808
rect 3525 83748 3529 83804
rect 3529 83748 3585 83804
rect 3585 83748 3589 83804
rect 3525 83744 3589 83748
rect 7952 83804 8016 83808
rect 7952 83748 7956 83804
rect 7956 83748 8012 83804
rect 8012 83748 8016 83804
rect 7952 83744 8016 83748
rect 8032 83804 8096 83808
rect 8032 83748 8036 83804
rect 8036 83748 8092 83804
rect 8092 83748 8096 83804
rect 8032 83744 8096 83748
rect 8112 83804 8176 83808
rect 8112 83748 8116 83804
rect 8116 83748 8172 83804
rect 8172 83748 8176 83804
rect 8112 83744 8176 83748
rect 8192 83804 8256 83808
rect 8192 83748 8196 83804
rect 8196 83748 8252 83804
rect 8252 83748 8256 83804
rect 8192 83744 8256 83748
rect 5618 83260 5682 83264
rect 5618 83204 5622 83260
rect 5622 83204 5678 83260
rect 5678 83204 5682 83260
rect 5618 83200 5682 83204
rect 5698 83260 5762 83264
rect 5698 83204 5702 83260
rect 5702 83204 5758 83260
rect 5758 83204 5762 83260
rect 5698 83200 5762 83204
rect 5778 83260 5842 83264
rect 5778 83204 5782 83260
rect 5782 83204 5838 83260
rect 5838 83204 5842 83260
rect 5778 83200 5842 83204
rect 5858 83260 5922 83264
rect 5858 83204 5862 83260
rect 5862 83204 5918 83260
rect 5918 83204 5922 83260
rect 5858 83200 5922 83204
rect 10285 83260 10349 83264
rect 10285 83204 10289 83260
rect 10289 83204 10345 83260
rect 10345 83204 10349 83260
rect 10285 83200 10349 83204
rect 10365 83260 10429 83264
rect 10365 83204 10369 83260
rect 10369 83204 10425 83260
rect 10425 83204 10429 83260
rect 10365 83200 10429 83204
rect 10445 83260 10509 83264
rect 10445 83204 10449 83260
rect 10449 83204 10505 83260
rect 10505 83204 10509 83260
rect 10445 83200 10509 83204
rect 10525 83260 10589 83264
rect 10525 83204 10529 83260
rect 10529 83204 10585 83260
rect 10585 83204 10589 83260
rect 10525 83200 10589 83204
rect 3285 82716 3349 82720
rect 3285 82660 3289 82716
rect 3289 82660 3345 82716
rect 3345 82660 3349 82716
rect 3285 82656 3349 82660
rect 3365 82716 3429 82720
rect 3365 82660 3369 82716
rect 3369 82660 3425 82716
rect 3425 82660 3429 82716
rect 3365 82656 3429 82660
rect 3445 82716 3509 82720
rect 3445 82660 3449 82716
rect 3449 82660 3505 82716
rect 3505 82660 3509 82716
rect 3445 82656 3509 82660
rect 3525 82716 3589 82720
rect 3525 82660 3529 82716
rect 3529 82660 3585 82716
rect 3585 82660 3589 82716
rect 3525 82656 3589 82660
rect 7952 82716 8016 82720
rect 7952 82660 7956 82716
rect 7956 82660 8012 82716
rect 8012 82660 8016 82716
rect 7952 82656 8016 82660
rect 8032 82716 8096 82720
rect 8032 82660 8036 82716
rect 8036 82660 8092 82716
rect 8092 82660 8096 82716
rect 8032 82656 8096 82660
rect 8112 82716 8176 82720
rect 8112 82660 8116 82716
rect 8116 82660 8172 82716
rect 8172 82660 8176 82716
rect 8112 82656 8176 82660
rect 8192 82716 8256 82720
rect 8192 82660 8196 82716
rect 8196 82660 8252 82716
rect 8252 82660 8256 82716
rect 8192 82656 8256 82660
rect 5618 82172 5682 82176
rect 5618 82116 5622 82172
rect 5622 82116 5678 82172
rect 5678 82116 5682 82172
rect 5618 82112 5682 82116
rect 5698 82172 5762 82176
rect 5698 82116 5702 82172
rect 5702 82116 5758 82172
rect 5758 82116 5762 82172
rect 5698 82112 5762 82116
rect 5778 82172 5842 82176
rect 5778 82116 5782 82172
rect 5782 82116 5838 82172
rect 5838 82116 5842 82172
rect 5778 82112 5842 82116
rect 5858 82172 5922 82176
rect 5858 82116 5862 82172
rect 5862 82116 5918 82172
rect 5918 82116 5922 82172
rect 5858 82112 5922 82116
rect 10285 82172 10349 82176
rect 10285 82116 10289 82172
rect 10289 82116 10345 82172
rect 10345 82116 10349 82172
rect 10285 82112 10349 82116
rect 10365 82172 10429 82176
rect 10365 82116 10369 82172
rect 10369 82116 10425 82172
rect 10425 82116 10429 82172
rect 10365 82112 10429 82116
rect 10445 82172 10509 82176
rect 10445 82116 10449 82172
rect 10449 82116 10505 82172
rect 10505 82116 10509 82172
rect 10445 82112 10509 82116
rect 10525 82172 10589 82176
rect 10525 82116 10529 82172
rect 10529 82116 10585 82172
rect 10585 82116 10589 82172
rect 10525 82112 10589 82116
rect 3285 81628 3349 81632
rect 3285 81572 3289 81628
rect 3289 81572 3345 81628
rect 3345 81572 3349 81628
rect 3285 81568 3349 81572
rect 3365 81628 3429 81632
rect 3365 81572 3369 81628
rect 3369 81572 3425 81628
rect 3425 81572 3429 81628
rect 3365 81568 3429 81572
rect 3445 81628 3509 81632
rect 3445 81572 3449 81628
rect 3449 81572 3505 81628
rect 3505 81572 3509 81628
rect 3445 81568 3509 81572
rect 3525 81628 3589 81632
rect 3525 81572 3529 81628
rect 3529 81572 3585 81628
rect 3585 81572 3589 81628
rect 3525 81568 3589 81572
rect 7952 81628 8016 81632
rect 7952 81572 7956 81628
rect 7956 81572 8012 81628
rect 8012 81572 8016 81628
rect 7952 81568 8016 81572
rect 8032 81628 8096 81632
rect 8032 81572 8036 81628
rect 8036 81572 8092 81628
rect 8092 81572 8096 81628
rect 8032 81568 8096 81572
rect 8112 81628 8176 81632
rect 8112 81572 8116 81628
rect 8116 81572 8172 81628
rect 8172 81572 8176 81628
rect 8112 81568 8176 81572
rect 8192 81628 8256 81632
rect 8192 81572 8196 81628
rect 8196 81572 8252 81628
rect 8252 81572 8256 81628
rect 8192 81568 8256 81572
rect 5618 81084 5682 81088
rect 5618 81028 5622 81084
rect 5622 81028 5678 81084
rect 5678 81028 5682 81084
rect 5618 81024 5682 81028
rect 5698 81084 5762 81088
rect 5698 81028 5702 81084
rect 5702 81028 5758 81084
rect 5758 81028 5762 81084
rect 5698 81024 5762 81028
rect 5778 81084 5842 81088
rect 5778 81028 5782 81084
rect 5782 81028 5838 81084
rect 5838 81028 5842 81084
rect 5778 81024 5842 81028
rect 5858 81084 5922 81088
rect 5858 81028 5862 81084
rect 5862 81028 5918 81084
rect 5918 81028 5922 81084
rect 5858 81024 5922 81028
rect 10285 81084 10349 81088
rect 10285 81028 10289 81084
rect 10289 81028 10345 81084
rect 10345 81028 10349 81084
rect 10285 81024 10349 81028
rect 10365 81084 10429 81088
rect 10365 81028 10369 81084
rect 10369 81028 10425 81084
rect 10425 81028 10429 81084
rect 10365 81024 10429 81028
rect 10445 81084 10509 81088
rect 10445 81028 10449 81084
rect 10449 81028 10505 81084
rect 10505 81028 10509 81084
rect 10445 81024 10509 81028
rect 10525 81084 10589 81088
rect 10525 81028 10529 81084
rect 10529 81028 10585 81084
rect 10585 81028 10589 81084
rect 10525 81024 10589 81028
rect 3285 80540 3349 80544
rect 3285 80484 3289 80540
rect 3289 80484 3345 80540
rect 3345 80484 3349 80540
rect 3285 80480 3349 80484
rect 3365 80540 3429 80544
rect 3365 80484 3369 80540
rect 3369 80484 3425 80540
rect 3425 80484 3429 80540
rect 3365 80480 3429 80484
rect 3445 80540 3509 80544
rect 3445 80484 3449 80540
rect 3449 80484 3505 80540
rect 3505 80484 3509 80540
rect 3445 80480 3509 80484
rect 3525 80540 3589 80544
rect 3525 80484 3529 80540
rect 3529 80484 3585 80540
rect 3585 80484 3589 80540
rect 3525 80480 3589 80484
rect 7952 80540 8016 80544
rect 7952 80484 7956 80540
rect 7956 80484 8012 80540
rect 8012 80484 8016 80540
rect 7952 80480 8016 80484
rect 8032 80540 8096 80544
rect 8032 80484 8036 80540
rect 8036 80484 8092 80540
rect 8092 80484 8096 80540
rect 8032 80480 8096 80484
rect 8112 80540 8176 80544
rect 8112 80484 8116 80540
rect 8116 80484 8172 80540
rect 8172 80484 8176 80540
rect 8112 80480 8176 80484
rect 8192 80540 8256 80544
rect 8192 80484 8196 80540
rect 8196 80484 8252 80540
rect 8252 80484 8256 80540
rect 8192 80480 8256 80484
rect 5618 79996 5682 80000
rect 5618 79940 5622 79996
rect 5622 79940 5678 79996
rect 5678 79940 5682 79996
rect 5618 79936 5682 79940
rect 5698 79996 5762 80000
rect 5698 79940 5702 79996
rect 5702 79940 5758 79996
rect 5758 79940 5762 79996
rect 5698 79936 5762 79940
rect 5778 79996 5842 80000
rect 5778 79940 5782 79996
rect 5782 79940 5838 79996
rect 5838 79940 5842 79996
rect 5778 79936 5842 79940
rect 5858 79996 5922 80000
rect 5858 79940 5862 79996
rect 5862 79940 5918 79996
rect 5918 79940 5922 79996
rect 5858 79936 5922 79940
rect 10285 79996 10349 80000
rect 10285 79940 10289 79996
rect 10289 79940 10345 79996
rect 10345 79940 10349 79996
rect 10285 79936 10349 79940
rect 10365 79996 10429 80000
rect 10365 79940 10369 79996
rect 10369 79940 10425 79996
rect 10425 79940 10429 79996
rect 10365 79936 10429 79940
rect 10445 79996 10509 80000
rect 10445 79940 10449 79996
rect 10449 79940 10505 79996
rect 10505 79940 10509 79996
rect 10445 79936 10509 79940
rect 10525 79996 10589 80000
rect 10525 79940 10529 79996
rect 10529 79940 10585 79996
rect 10585 79940 10589 79996
rect 10525 79936 10589 79940
rect 3285 79452 3349 79456
rect 3285 79396 3289 79452
rect 3289 79396 3345 79452
rect 3345 79396 3349 79452
rect 3285 79392 3349 79396
rect 3365 79452 3429 79456
rect 3365 79396 3369 79452
rect 3369 79396 3425 79452
rect 3425 79396 3429 79452
rect 3365 79392 3429 79396
rect 3445 79452 3509 79456
rect 3445 79396 3449 79452
rect 3449 79396 3505 79452
rect 3505 79396 3509 79452
rect 3445 79392 3509 79396
rect 3525 79452 3589 79456
rect 3525 79396 3529 79452
rect 3529 79396 3585 79452
rect 3585 79396 3589 79452
rect 3525 79392 3589 79396
rect 7952 79452 8016 79456
rect 7952 79396 7956 79452
rect 7956 79396 8012 79452
rect 8012 79396 8016 79452
rect 7952 79392 8016 79396
rect 8032 79452 8096 79456
rect 8032 79396 8036 79452
rect 8036 79396 8092 79452
rect 8092 79396 8096 79452
rect 8032 79392 8096 79396
rect 8112 79452 8176 79456
rect 8112 79396 8116 79452
rect 8116 79396 8172 79452
rect 8172 79396 8176 79452
rect 8112 79392 8176 79396
rect 8192 79452 8256 79456
rect 8192 79396 8196 79452
rect 8196 79396 8252 79452
rect 8252 79396 8256 79452
rect 8192 79392 8256 79396
rect 5618 78908 5682 78912
rect 5618 78852 5622 78908
rect 5622 78852 5678 78908
rect 5678 78852 5682 78908
rect 5618 78848 5682 78852
rect 5698 78908 5762 78912
rect 5698 78852 5702 78908
rect 5702 78852 5758 78908
rect 5758 78852 5762 78908
rect 5698 78848 5762 78852
rect 5778 78908 5842 78912
rect 5778 78852 5782 78908
rect 5782 78852 5838 78908
rect 5838 78852 5842 78908
rect 5778 78848 5842 78852
rect 5858 78908 5922 78912
rect 5858 78852 5862 78908
rect 5862 78852 5918 78908
rect 5918 78852 5922 78908
rect 5858 78848 5922 78852
rect 10285 78908 10349 78912
rect 10285 78852 10289 78908
rect 10289 78852 10345 78908
rect 10345 78852 10349 78908
rect 10285 78848 10349 78852
rect 10365 78908 10429 78912
rect 10365 78852 10369 78908
rect 10369 78852 10425 78908
rect 10425 78852 10429 78908
rect 10365 78848 10429 78852
rect 10445 78908 10509 78912
rect 10445 78852 10449 78908
rect 10449 78852 10505 78908
rect 10505 78852 10509 78908
rect 10445 78848 10509 78852
rect 10525 78908 10589 78912
rect 10525 78852 10529 78908
rect 10529 78852 10585 78908
rect 10585 78852 10589 78908
rect 10525 78848 10589 78852
rect 3285 78364 3349 78368
rect 3285 78308 3289 78364
rect 3289 78308 3345 78364
rect 3345 78308 3349 78364
rect 3285 78304 3349 78308
rect 3365 78364 3429 78368
rect 3365 78308 3369 78364
rect 3369 78308 3425 78364
rect 3425 78308 3429 78364
rect 3365 78304 3429 78308
rect 3445 78364 3509 78368
rect 3445 78308 3449 78364
rect 3449 78308 3505 78364
rect 3505 78308 3509 78364
rect 3445 78304 3509 78308
rect 3525 78364 3589 78368
rect 3525 78308 3529 78364
rect 3529 78308 3585 78364
rect 3585 78308 3589 78364
rect 3525 78304 3589 78308
rect 7952 78364 8016 78368
rect 7952 78308 7956 78364
rect 7956 78308 8012 78364
rect 8012 78308 8016 78364
rect 7952 78304 8016 78308
rect 8032 78364 8096 78368
rect 8032 78308 8036 78364
rect 8036 78308 8092 78364
rect 8092 78308 8096 78364
rect 8032 78304 8096 78308
rect 8112 78364 8176 78368
rect 8112 78308 8116 78364
rect 8116 78308 8172 78364
rect 8172 78308 8176 78364
rect 8112 78304 8176 78308
rect 8192 78364 8256 78368
rect 8192 78308 8196 78364
rect 8196 78308 8252 78364
rect 8252 78308 8256 78364
rect 8192 78304 8256 78308
rect 5618 77820 5682 77824
rect 5618 77764 5622 77820
rect 5622 77764 5678 77820
rect 5678 77764 5682 77820
rect 5618 77760 5682 77764
rect 5698 77820 5762 77824
rect 5698 77764 5702 77820
rect 5702 77764 5758 77820
rect 5758 77764 5762 77820
rect 5698 77760 5762 77764
rect 5778 77820 5842 77824
rect 5778 77764 5782 77820
rect 5782 77764 5838 77820
rect 5838 77764 5842 77820
rect 5778 77760 5842 77764
rect 5858 77820 5922 77824
rect 5858 77764 5862 77820
rect 5862 77764 5918 77820
rect 5918 77764 5922 77820
rect 5858 77760 5922 77764
rect 10285 77820 10349 77824
rect 10285 77764 10289 77820
rect 10289 77764 10345 77820
rect 10345 77764 10349 77820
rect 10285 77760 10349 77764
rect 10365 77820 10429 77824
rect 10365 77764 10369 77820
rect 10369 77764 10425 77820
rect 10425 77764 10429 77820
rect 10365 77760 10429 77764
rect 10445 77820 10509 77824
rect 10445 77764 10449 77820
rect 10449 77764 10505 77820
rect 10505 77764 10509 77820
rect 10445 77760 10509 77764
rect 10525 77820 10589 77824
rect 10525 77764 10529 77820
rect 10529 77764 10585 77820
rect 10585 77764 10589 77820
rect 10525 77760 10589 77764
rect 3285 77276 3349 77280
rect 3285 77220 3289 77276
rect 3289 77220 3345 77276
rect 3345 77220 3349 77276
rect 3285 77216 3349 77220
rect 3365 77276 3429 77280
rect 3365 77220 3369 77276
rect 3369 77220 3425 77276
rect 3425 77220 3429 77276
rect 3365 77216 3429 77220
rect 3445 77276 3509 77280
rect 3445 77220 3449 77276
rect 3449 77220 3505 77276
rect 3505 77220 3509 77276
rect 3445 77216 3509 77220
rect 3525 77276 3589 77280
rect 3525 77220 3529 77276
rect 3529 77220 3585 77276
rect 3585 77220 3589 77276
rect 3525 77216 3589 77220
rect 7952 77276 8016 77280
rect 7952 77220 7956 77276
rect 7956 77220 8012 77276
rect 8012 77220 8016 77276
rect 7952 77216 8016 77220
rect 8032 77276 8096 77280
rect 8032 77220 8036 77276
rect 8036 77220 8092 77276
rect 8092 77220 8096 77276
rect 8032 77216 8096 77220
rect 8112 77276 8176 77280
rect 8112 77220 8116 77276
rect 8116 77220 8172 77276
rect 8172 77220 8176 77276
rect 8112 77216 8176 77220
rect 8192 77276 8256 77280
rect 8192 77220 8196 77276
rect 8196 77220 8252 77276
rect 8252 77220 8256 77276
rect 8192 77216 8256 77220
rect 5618 76732 5682 76736
rect 5618 76676 5622 76732
rect 5622 76676 5678 76732
rect 5678 76676 5682 76732
rect 5618 76672 5682 76676
rect 5698 76732 5762 76736
rect 5698 76676 5702 76732
rect 5702 76676 5758 76732
rect 5758 76676 5762 76732
rect 5698 76672 5762 76676
rect 5778 76732 5842 76736
rect 5778 76676 5782 76732
rect 5782 76676 5838 76732
rect 5838 76676 5842 76732
rect 5778 76672 5842 76676
rect 5858 76732 5922 76736
rect 5858 76676 5862 76732
rect 5862 76676 5918 76732
rect 5918 76676 5922 76732
rect 5858 76672 5922 76676
rect 10285 76732 10349 76736
rect 10285 76676 10289 76732
rect 10289 76676 10345 76732
rect 10345 76676 10349 76732
rect 10285 76672 10349 76676
rect 10365 76732 10429 76736
rect 10365 76676 10369 76732
rect 10369 76676 10425 76732
rect 10425 76676 10429 76732
rect 10365 76672 10429 76676
rect 10445 76732 10509 76736
rect 10445 76676 10449 76732
rect 10449 76676 10505 76732
rect 10505 76676 10509 76732
rect 10445 76672 10509 76676
rect 10525 76732 10589 76736
rect 10525 76676 10529 76732
rect 10529 76676 10585 76732
rect 10585 76676 10589 76732
rect 10525 76672 10589 76676
rect 3285 76188 3349 76192
rect 3285 76132 3289 76188
rect 3289 76132 3345 76188
rect 3345 76132 3349 76188
rect 3285 76128 3349 76132
rect 3365 76188 3429 76192
rect 3365 76132 3369 76188
rect 3369 76132 3425 76188
rect 3425 76132 3429 76188
rect 3365 76128 3429 76132
rect 3445 76188 3509 76192
rect 3445 76132 3449 76188
rect 3449 76132 3505 76188
rect 3505 76132 3509 76188
rect 3445 76128 3509 76132
rect 3525 76188 3589 76192
rect 3525 76132 3529 76188
rect 3529 76132 3585 76188
rect 3585 76132 3589 76188
rect 3525 76128 3589 76132
rect 7952 76188 8016 76192
rect 7952 76132 7956 76188
rect 7956 76132 8012 76188
rect 8012 76132 8016 76188
rect 7952 76128 8016 76132
rect 8032 76188 8096 76192
rect 8032 76132 8036 76188
rect 8036 76132 8092 76188
rect 8092 76132 8096 76188
rect 8032 76128 8096 76132
rect 8112 76188 8176 76192
rect 8112 76132 8116 76188
rect 8116 76132 8172 76188
rect 8172 76132 8176 76188
rect 8112 76128 8176 76132
rect 8192 76188 8256 76192
rect 8192 76132 8196 76188
rect 8196 76132 8252 76188
rect 8252 76132 8256 76188
rect 8192 76128 8256 76132
rect 5618 75644 5682 75648
rect 5618 75588 5622 75644
rect 5622 75588 5678 75644
rect 5678 75588 5682 75644
rect 5618 75584 5682 75588
rect 5698 75644 5762 75648
rect 5698 75588 5702 75644
rect 5702 75588 5758 75644
rect 5758 75588 5762 75644
rect 5698 75584 5762 75588
rect 5778 75644 5842 75648
rect 5778 75588 5782 75644
rect 5782 75588 5838 75644
rect 5838 75588 5842 75644
rect 5778 75584 5842 75588
rect 5858 75644 5922 75648
rect 5858 75588 5862 75644
rect 5862 75588 5918 75644
rect 5918 75588 5922 75644
rect 5858 75584 5922 75588
rect 10285 75644 10349 75648
rect 10285 75588 10289 75644
rect 10289 75588 10345 75644
rect 10345 75588 10349 75644
rect 10285 75584 10349 75588
rect 10365 75644 10429 75648
rect 10365 75588 10369 75644
rect 10369 75588 10425 75644
rect 10425 75588 10429 75644
rect 10365 75584 10429 75588
rect 10445 75644 10509 75648
rect 10445 75588 10449 75644
rect 10449 75588 10505 75644
rect 10505 75588 10509 75644
rect 10445 75584 10509 75588
rect 10525 75644 10589 75648
rect 10525 75588 10529 75644
rect 10529 75588 10585 75644
rect 10585 75588 10589 75644
rect 10525 75584 10589 75588
rect 3285 75100 3349 75104
rect 3285 75044 3289 75100
rect 3289 75044 3345 75100
rect 3345 75044 3349 75100
rect 3285 75040 3349 75044
rect 3365 75100 3429 75104
rect 3365 75044 3369 75100
rect 3369 75044 3425 75100
rect 3425 75044 3429 75100
rect 3365 75040 3429 75044
rect 3445 75100 3509 75104
rect 3445 75044 3449 75100
rect 3449 75044 3505 75100
rect 3505 75044 3509 75100
rect 3445 75040 3509 75044
rect 3525 75100 3589 75104
rect 3525 75044 3529 75100
rect 3529 75044 3585 75100
rect 3585 75044 3589 75100
rect 3525 75040 3589 75044
rect 7952 75100 8016 75104
rect 7952 75044 7956 75100
rect 7956 75044 8012 75100
rect 8012 75044 8016 75100
rect 7952 75040 8016 75044
rect 8032 75100 8096 75104
rect 8032 75044 8036 75100
rect 8036 75044 8092 75100
rect 8092 75044 8096 75100
rect 8032 75040 8096 75044
rect 8112 75100 8176 75104
rect 8112 75044 8116 75100
rect 8116 75044 8172 75100
rect 8172 75044 8176 75100
rect 8112 75040 8176 75044
rect 8192 75100 8256 75104
rect 8192 75044 8196 75100
rect 8196 75044 8252 75100
rect 8252 75044 8256 75100
rect 8192 75040 8256 75044
rect 5618 74556 5682 74560
rect 5618 74500 5622 74556
rect 5622 74500 5678 74556
rect 5678 74500 5682 74556
rect 5618 74496 5682 74500
rect 5698 74556 5762 74560
rect 5698 74500 5702 74556
rect 5702 74500 5758 74556
rect 5758 74500 5762 74556
rect 5698 74496 5762 74500
rect 5778 74556 5842 74560
rect 5778 74500 5782 74556
rect 5782 74500 5838 74556
rect 5838 74500 5842 74556
rect 5778 74496 5842 74500
rect 5858 74556 5922 74560
rect 5858 74500 5862 74556
rect 5862 74500 5918 74556
rect 5918 74500 5922 74556
rect 5858 74496 5922 74500
rect 10285 74556 10349 74560
rect 10285 74500 10289 74556
rect 10289 74500 10345 74556
rect 10345 74500 10349 74556
rect 10285 74496 10349 74500
rect 10365 74556 10429 74560
rect 10365 74500 10369 74556
rect 10369 74500 10425 74556
rect 10425 74500 10429 74556
rect 10365 74496 10429 74500
rect 10445 74556 10509 74560
rect 10445 74500 10449 74556
rect 10449 74500 10505 74556
rect 10505 74500 10509 74556
rect 10445 74496 10509 74500
rect 10525 74556 10589 74560
rect 10525 74500 10529 74556
rect 10529 74500 10585 74556
rect 10585 74500 10589 74556
rect 10525 74496 10589 74500
rect 3285 74012 3349 74016
rect 3285 73956 3289 74012
rect 3289 73956 3345 74012
rect 3345 73956 3349 74012
rect 3285 73952 3349 73956
rect 3365 74012 3429 74016
rect 3365 73956 3369 74012
rect 3369 73956 3425 74012
rect 3425 73956 3429 74012
rect 3365 73952 3429 73956
rect 3445 74012 3509 74016
rect 3445 73956 3449 74012
rect 3449 73956 3505 74012
rect 3505 73956 3509 74012
rect 3445 73952 3509 73956
rect 3525 74012 3589 74016
rect 3525 73956 3529 74012
rect 3529 73956 3585 74012
rect 3585 73956 3589 74012
rect 3525 73952 3589 73956
rect 7952 74012 8016 74016
rect 7952 73956 7956 74012
rect 7956 73956 8012 74012
rect 8012 73956 8016 74012
rect 7952 73952 8016 73956
rect 8032 74012 8096 74016
rect 8032 73956 8036 74012
rect 8036 73956 8092 74012
rect 8092 73956 8096 74012
rect 8032 73952 8096 73956
rect 8112 74012 8176 74016
rect 8112 73956 8116 74012
rect 8116 73956 8172 74012
rect 8172 73956 8176 74012
rect 8112 73952 8176 73956
rect 8192 74012 8256 74016
rect 8192 73956 8196 74012
rect 8196 73956 8252 74012
rect 8252 73956 8256 74012
rect 8192 73952 8256 73956
rect 5618 73468 5682 73472
rect 5618 73412 5622 73468
rect 5622 73412 5678 73468
rect 5678 73412 5682 73468
rect 5618 73408 5682 73412
rect 5698 73468 5762 73472
rect 5698 73412 5702 73468
rect 5702 73412 5758 73468
rect 5758 73412 5762 73468
rect 5698 73408 5762 73412
rect 5778 73468 5842 73472
rect 5778 73412 5782 73468
rect 5782 73412 5838 73468
rect 5838 73412 5842 73468
rect 5778 73408 5842 73412
rect 5858 73468 5922 73472
rect 5858 73412 5862 73468
rect 5862 73412 5918 73468
rect 5918 73412 5922 73468
rect 5858 73408 5922 73412
rect 10285 73468 10349 73472
rect 10285 73412 10289 73468
rect 10289 73412 10345 73468
rect 10345 73412 10349 73468
rect 10285 73408 10349 73412
rect 10365 73468 10429 73472
rect 10365 73412 10369 73468
rect 10369 73412 10425 73468
rect 10425 73412 10429 73468
rect 10365 73408 10429 73412
rect 10445 73468 10509 73472
rect 10445 73412 10449 73468
rect 10449 73412 10505 73468
rect 10505 73412 10509 73468
rect 10445 73408 10509 73412
rect 10525 73468 10589 73472
rect 10525 73412 10529 73468
rect 10529 73412 10585 73468
rect 10585 73412 10589 73468
rect 10525 73408 10589 73412
rect 3285 72924 3349 72928
rect 3285 72868 3289 72924
rect 3289 72868 3345 72924
rect 3345 72868 3349 72924
rect 3285 72864 3349 72868
rect 3365 72924 3429 72928
rect 3365 72868 3369 72924
rect 3369 72868 3425 72924
rect 3425 72868 3429 72924
rect 3365 72864 3429 72868
rect 3445 72924 3509 72928
rect 3445 72868 3449 72924
rect 3449 72868 3505 72924
rect 3505 72868 3509 72924
rect 3445 72864 3509 72868
rect 3525 72924 3589 72928
rect 3525 72868 3529 72924
rect 3529 72868 3585 72924
rect 3585 72868 3589 72924
rect 3525 72864 3589 72868
rect 7952 72924 8016 72928
rect 7952 72868 7956 72924
rect 7956 72868 8012 72924
rect 8012 72868 8016 72924
rect 7952 72864 8016 72868
rect 8032 72924 8096 72928
rect 8032 72868 8036 72924
rect 8036 72868 8092 72924
rect 8092 72868 8096 72924
rect 8032 72864 8096 72868
rect 8112 72924 8176 72928
rect 8112 72868 8116 72924
rect 8116 72868 8172 72924
rect 8172 72868 8176 72924
rect 8112 72864 8176 72868
rect 8192 72924 8256 72928
rect 8192 72868 8196 72924
rect 8196 72868 8252 72924
rect 8252 72868 8256 72924
rect 8192 72864 8256 72868
rect 5618 72380 5682 72384
rect 5618 72324 5622 72380
rect 5622 72324 5678 72380
rect 5678 72324 5682 72380
rect 5618 72320 5682 72324
rect 5698 72380 5762 72384
rect 5698 72324 5702 72380
rect 5702 72324 5758 72380
rect 5758 72324 5762 72380
rect 5698 72320 5762 72324
rect 5778 72380 5842 72384
rect 5778 72324 5782 72380
rect 5782 72324 5838 72380
rect 5838 72324 5842 72380
rect 5778 72320 5842 72324
rect 5858 72380 5922 72384
rect 5858 72324 5862 72380
rect 5862 72324 5918 72380
rect 5918 72324 5922 72380
rect 5858 72320 5922 72324
rect 10285 72380 10349 72384
rect 10285 72324 10289 72380
rect 10289 72324 10345 72380
rect 10345 72324 10349 72380
rect 10285 72320 10349 72324
rect 10365 72380 10429 72384
rect 10365 72324 10369 72380
rect 10369 72324 10425 72380
rect 10425 72324 10429 72380
rect 10365 72320 10429 72324
rect 10445 72380 10509 72384
rect 10445 72324 10449 72380
rect 10449 72324 10505 72380
rect 10505 72324 10509 72380
rect 10445 72320 10509 72324
rect 10525 72380 10589 72384
rect 10525 72324 10529 72380
rect 10529 72324 10585 72380
rect 10585 72324 10589 72380
rect 10525 72320 10589 72324
rect 3285 71836 3349 71840
rect 3285 71780 3289 71836
rect 3289 71780 3345 71836
rect 3345 71780 3349 71836
rect 3285 71776 3349 71780
rect 3365 71836 3429 71840
rect 3365 71780 3369 71836
rect 3369 71780 3425 71836
rect 3425 71780 3429 71836
rect 3365 71776 3429 71780
rect 3445 71836 3509 71840
rect 3445 71780 3449 71836
rect 3449 71780 3505 71836
rect 3505 71780 3509 71836
rect 3445 71776 3509 71780
rect 3525 71836 3589 71840
rect 3525 71780 3529 71836
rect 3529 71780 3585 71836
rect 3585 71780 3589 71836
rect 3525 71776 3589 71780
rect 7952 71836 8016 71840
rect 7952 71780 7956 71836
rect 7956 71780 8012 71836
rect 8012 71780 8016 71836
rect 7952 71776 8016 71780
rect 8032 71836 8096 71840
rect 8032 71780 8036 71836
rect 8036 71780 8092 71836
rect 8092 71780 8096 71836
rect 8032 71776 8096 71780
rect 8112 71836 8176 71840
rect 8112 71780 8116 71836
rect 8116 71780 8172 71836
rect 8172 71780 8176 71836
rect 8112 71776 8176 71780
rect 8192 71836 8256 71840
rect 8192 71780 8196 71836
rect 8196 71780 8252 71836
rect 8252 71780 8256 71836
rect 8192 71776 8256 71780
rect 5618 71292 5682 71296
rect 5618 71236 5622 71292
rect 5622 71236 5678 71292
rect 5678 71236 5682 71292
rect 5618 71232 5682 71236
rect 5698 71292 5762 71296
rect 5698 71236 5702 71292
rect 5702 71236 5758 71292
rect 5758 71236 5762 71292
rect 5698 71232 5762 71236
rect 5778 71292 5842 71296
rect 5778 71236 5782 71292
rect 5782 71236 5838 71292
rect 5838 71236 5842 71292
rect 5778 71232 5842 71236
rect 5858 71292 5922 71296
rect 5858 71236 5862 71292
rect 5862 71236 5918 71292
rect 5918 71236 5922 71292
rect 5858 71232 5922 71236
rect 10285 71292 10349 71296
rect 10285 71236 10289 71292
rect 10289 71236 10345 71292
rect 10345 71236 10349 71292
rect 10285 71232 10349 71236
rect 10365 71292 10429 71296
rect 10365 71236 10369 71292
rect 10369 71236 10425 71292
rect 10425 71236 10429 71292
rect 10365 71232 10429 71236
rect 10445 71292 10509 71296
rect 10445 71236 10449 71292
rect 10449 71236 10505 71292
rect 10505 71236 10509 71292
rect 10445 71232 10509 71236
rect 10525 71292 10589 71296
rect 10525 71236 10529 71292
rect 10529 71236 10585 71292
rect 10585 71236 10589 71292
rect 10525 71232 10589 71236
rect 3285 70748 3349 70752
rect 3285 70692 3289 70748
rect 3289 70692 3345 70748
rect 3345 70692 3349 70748
rect 3285 70688 3349 70692
rect 3365 70748 3429 70752
rect 3365 70692 3369 70748
rect 3369 70692 3425 70748
rect 3425 70692 3429 70748
rect 3365 70688 3429 70692
rect 3445 70748 3509 70752
rect 3445 70692 3449 70748
rect 3449 70692 3505 70748
rect 3505 70692 3509 70748
rect 3445 70688 3509 70692
rect 3525 70748 3589 70752
rect 3525 70692 3529 70748
rect 3529 70692 3585 70748
rect 3585 70692 3589 70748
rect 3525 70688 3589 70692
rect 7952 70748 8016 70752
rect 7952 70692 7956 70748
rect 7956 70692 8012 70748
rect 8012 70692 8016 70748
rect 7952 70688 8016 70692
rect 8032 70748 8096 70752
rect 8032 70692 8036 70748
rect 8036 70692 8092 70748
rect 8092 70692 8096 70748
rect 8032 70688 8096 70692
rect 8112 70748 8176 70752
rect 8112 70692 8116 70748
rect 8116 70692 8172 70748
rect 8172 70692 8176 70748
rect 8112 70688 8176 70692
rect 8192 70748 8256 70752
rect 8192 70692 8196 70748
rect 8196 70692 8252 70748
rect 8252 70692 8256 70748
rect 8192 70688 8256 70692
rect 5618 70204 5682 70208
rect 5618 70148 5622 70204
rect 5622 70148 5678 70204
rect 5678 70148 5682 70204
rect 5618 70144 5682 70148
rect 5698 70204 5762 70208
rect 5698 70148 5702 70204
rect 5702 70148 5758 70204
rect 5758 70148 5762 70204
rect 5698 70144 5762 70148
rect 5778 70204 5842 70208
rect 5778 70148 5782 70204
rect 5782 70148 5838 70204
rect 5838 70148 5842 70204
rect 5778 70144 5842 70148
rect 5858 70204 5922 70208
rect 5858 70148 5862 70204
rect 5862 70148 5918 70204
rect 5918 70148 5922 70204
rect 5858 70144 5922 70148
rect 10285 70204 10349 70208
rect 10285 70148 10289 70204
rect 10289 70148 10345 70204
rect 10345 70148 10349 70204
rect 10285 70144 10349 70148
rect 10365 70204 10429 70208
rect 10365 70148 10369 70204
rect 10369 70148 10425 70204
rect 10425 70148 10429 70204
rect 10365 70144 10429 70148
rect 10445 70204 10509 70208
rect 10445 70148 10449 70204
rect 10449 70148 10505 70204
rect 10505 70148 10509 70204
rect 10445 70144 10509 70148
rect 10525 70204 10589 70208
rect 10525 70148 10529 70204
rect 10529 70148 10585 70204
rect 10585 70148 10589 70204
rect 10525 70144 10589 70148
rect 3285 69660 3349 69664
rect 3285 69604 3289 69660
rect 3289 69604 3345 69660
rect 3345 69604 3349 69660
rect 3285 69600 3349 69604
rect 3365 69660 3429 69664
rect 3365 69604 3369 69660
rect 3369 69604 3425 69660
rect 3425 69604 3429 69660
rect 3365 69600 3429 69604
rect 3445 69660 3509 69664
rect 3445 69604 3449 69660
rect 3449 69604 3505 69660
rect 3505 69604 3509 69660
rect 3445 69600 3509 69604
rect 3525 69660 3589 69664
rect 3525 69604 3529 69660
rect 3529 69604 3585 69660
rect 3585 69604 3589 69660
rect 3525 69600 3589 69604
rect 7952 69660 8016 69664
rect 7952 69604 7956 69660
rect 7956 69604 8012 69660
rect 8012 69604 8016 69660
rect 7952 69600 8016 69604
rect 8032 69660 8096 69664
rect 8032 69604 8036 69660
rect 8036 69604 8092 69660
rect 8092 69604 8096 69660
rect 8032 69600 8096 69604
rect 8112 69660 8176 69664
rect 8112 69604 8116 69660
rect 8116 69604 8172 69660
rect 8172 69604 8176 69660
rect 8112 69600 8176 69604
rect 8192 69660 8256 69664
rect 8192 69604 8196 69660
rect 8196 69604 8252 69660
rect 8252 69604 8256 69660
rect 8192 69600 8256 69604
rect 5618 69116 5682 69120
rect 5618 69060 5622 69116
rect 5622 69060 5678 69116
rect 5678 69060 5682 69116
rect 5618 69056 5682 69060
rect 5698 69116 5762 69120
rect 5698 69060 5702 69116
rect 5702 69060 5758 69116
rect 5758 69060 5762 69116
rect 5698 69056 5762 69060
rect 5778 69116 5842 69120
rect 5778 69060 5782 69116
rect 5782 69060 5838 69116
rect 5838 69060 5842 69116
rect 5778 69056 5842 69060
rect 5858 69116 5922 69120
rect 5858 69060 5862 69116
rect 5862 69060 5918 69116
rect 5918 69060 5922 69116
rect 5858 69056 5922 69060
rect 10285 69116 10349 69120
rect 10285 69060 10289 69116
rect 10289 69060 10345 69116
rect 10345 69060 10349 69116
rect 10285 69056 10349 69060
rect 10365 69116 10429 69120
rect 10365 69060 10369 69116
rect 10369 69060 10425 69116
rect 10425 69060 10429 69116
rect 10365 69056 10429 69060
rect 10445 69116 10509 69120
rect 10445 69060 10449 69116
rect 10449 69060 10505 69116
rect 10505 69060 10509 69116
rect 10445 69056 10509 69060
rect 10525 69116 10589 69120
rect 10525 69060 10529 69116
rect 10529 69060 10585 69116
rect 10585 69060 10589 69116
rect 10525 69056 10589 69060
rect 3285 68572 3349 68576
rect 3285 68516 3289 68572
rect 3289 68516 3345 68572
rect 3345 68516 3349 68572
rect 3285 68512 3349 68516
rect 3365 68572 3429 68576
rect 3365 68516 3369 68572
rect 3369 68516 3425 68572
rect 3425 68516 3429 68572
rect 3365 68512 3429 68516
rect 3445 68572 3509 68576
rect 3445 68516 3449 68572
rect 3449 68516 3505 68572
rect 3505 68516 3509 68572
rect 3445 68512 3509 68516
rect 3525 68572 3589 68576
rect 3525 68516 3529 68572
rect 3529 68516 3585 68572
rect 3585 68516 3589 68572
rect 3525 68512 3589 68516
rect 7952 68572 8016 68576
rect 7952 68516 7956 68572
rect 7956 68516 8012 68572
rect 8012 68516 8016 68572
rect 7952 68512 8016 68516
rect 8032 68572 8096 68576
rect 8032 68516 8036 68572
rect 8036 68516 8092 68572
rect 8092 68516 8096 68572
rect 8032 68512 8096 68516
rect 8112 68572 8176 68576
rect 8112 68516 8116 68572
rect 8116 68516 8172 68572
rect 8172 68516 8176 68572
rect 8112 68512 8176 68516
rect 8192 68572 8256 68576
rect 8192 68516 8196 68572
rect 8196 68516 8252 68572
rect 8252 68516 8256 68572
rect 8192 68512 8256 68516
rect 5618 68028 5682 68032
rect 5618 67972 5622 68028
rect 5622 67972 5678 68028
rect 5678 67972 5682 68028
rect 5618 67968 5682 67972
rect 5698 68028 5762 68032
rect 5698 67972 5702 68028
rect 5702 67972 5758 68028
rect 5758 67972 5762 68028
rect 5698 67968 5762 67972
rect 5778 68028 5842 68032
rect 5778 67972 5782 68028
rect 5782 67972 5838 68028
rect 5838 67972 5842 68028
rect 5778 67968 5842 67972
rect 5858 68028 5922 68032
rect 5858 67972 5862 68028
rect 5862 67972 5918 68028
rect 5918 67972 5922 68028
rect 5858 67968 5922 67972
rect 10285 68028 10349 68032
rect 10285 67972 10289 68028
rect 10289 67972 10345 68028
rect 10345 67972 10349 68028
rect 10285 67968 10349 67972
rect 10365 68028 10429 68032
rect 10365 67972 10369 68028
rect 10369 67972 10425 68028
rect 10425 67972 10429 68028
rect 10365 67968 10429 67972
rect 10445 68028 10509 68032
rect 10445 67972 10449 68028
rect 10449 67972 10505 68028
rect 10505 67972 10509 68028
rect 10445 67968 10509 67972
rect 10525 68028 10589 68032
rect 10525 67972 10529 68028
rect 10529 67972 10585 68028
rect 10585 67972 10589 68028
rect 10525 67968 10589 67972
rect 3285 67484 3349 67488
rect 3285 67428 3289 67484
rect 3289 67428 3345 67484
rect 3345 67428 3349 67484
rect 3285 67424 3349 67428
rect 3365 67484 3429 67488
rect 3365 67428 3369 67484
rect 3369 67428 3425 67484
rect 3425 67428 3429 67484
rect 3365 67424 3429 67428
rect 3445 67484 3509 67488
rect 3445 67428 3449 67484
rect 3449 67428 3505 67484
rect 3505 67428 3509 67484
rect 3445 67424 3509 67428
rect 3525 67484 3589 67488
rect 3525 67428 3529 67484
rect 3529 67428 3585 67484
rect 3585 67428 3589 67484
rect 3525 67424 3589 67428
rect 7952 67484 8016 67488
rect 7952 67428 7956 67484
rect 7956 67428 8012 67484
rect 8012 67428 8016 67484
rect 7952 67424 8016 67428
rect 8032 67484 8096 67488
rect 8032 67428 8036 67484
rect 8036 67428 8092 67484
rect 8092 67428 8096 67484
rect 8032 67424 8096 67428
rect 8112 67484 8176 67488
rect 8112 67428 8116 67484
rect 8116 67428 8172 67484
rect 8172 67428 8176 67484
rect 8112 67424 8176 67428
rect 8192 67484 8256 67488
rect 8192 67428 8196 67484
rect 8196 67428 8252 67484
rect 8252 67428 8256 67484
rect 8192 67424 8256 67428
rect 5618 66940 5682 66944
rect 5618 66884 5622 66940
rect 5622 66884 5678 66940
rect 5678 66884 5682 66940
rect 5618 66880 5682 66884
rect 5698 66940 5762 66944
rect 5698 66884 5702 66940
rect 5702 66884 5758 66940
rect 5758 66884 5762 66940
rect 5698 66880 5762 66884
rect 5778 66940 5842 66944
rect 5778 66884 5782 66940
rect 5782 66884 5838 66940
rect 5838 66884 5842 66940
rect 5778 66880 5842 66884
rect 5858 66940 5922 66944
rect 5858 66884 5862 66940
rect 5862 66884 5918 66940
rect 5918 66884 5922 66940
rect 5858 66880 5922 66884
rect 10285 66940 10349 66944
rect 10285 66884 10289 66940
rect 10289 66884 10345 66940
rect 10345 66884 10349 66940
rect 10285 66880 10349 66884
rect 10365 66940 10429 66944
rect 10365 66884 10369 66940
rect 10369 66884 10425 66940
rect 10425 66884 10429 66940
rect 10365 66880 10429 66884
rect 10445 66940 10509 66944
rect 10445 66884 10449 66940
rect 10449 66884 10505 66940
rect 10505 66884 10509 66940
rect 10445 66880 10509 66884
rect 10525 66940 10589 66944
rect 10525 66884 10529 66940
rect 10529 66884 10585 66940
rect 10585 66884 10589 66940
rect 10525 66880 10589 66884
rect 3285 66396 3349 66400
rect 3285 66340 3289 66396
rect 3289 66340 3345 66396
rect 3345 66340 3349 66396
rect 3285 66336 3349 66340
rect 3365 66396 3429 66400
rect 3365 66340 3369 66396
rect 3369 66340 3425 66396
rect 3425 66340 3429 66396
rect 3365 66336 3429 66340
rect 3445 66396 3509 66400
rect 3445 66340 3449 66396
rect 3449 66340 3505 66396
rect 3505 66340 3509 66396
rect 3445 66336 3509 66340
rect 3525 66396 3589 66400
rect 3525 66340 3529 66396
rect 3529 66340 3585 66396
rect 3585 66340 3589 66396
rect 3525 66336 3589 66340
rect 7952 66396 8016 66400
rect 7952 66340 7956 66396
rect 7956 66340 8012 66396
rect 8012 66340 8016 66396
rect 7952 66336 8016 66340
rect 8032 66396 8096 66400
rect 8032 66340 8036 66396
rect 8036 66340 8092 66396
rect 8092 66340 8096 66396
rect 8032 66336 8096 66340
rect 8112 66396 8176 66400
rect 8112 66340 8116 66396
rect 8116 66340 8172 66396
rect 8172 66340 8176 66396
rect 8112 66336 8176 66340
rect 8192 66396 8256 66400
rect 8192 66340 8196 66396
rect 8196 66340 8252 66396
rect 8252 66340 8256 66396
rect 8192 66336 8256 66340
rect 5618 65852 5682 65856
rect 5618 65796 5622 65852
rect 5622 65796 5678 65852
rect 5678 65796 5682 65852
rect 5618 65792 5682 65796
rect 5698 65852 5762 65856
rect 5698 65796 5702 65852
rect 5702 65796 5758 65852
rect 5758 65796 5762 65852
rect 5698 65792 5762 65796
rect 5778 65852 5842 65856
rect 5778 65796 5782 65852
rect 5782 65796 5838 65852
rect 5838 65796 5842 65852
rect 5778 65792 5842 65796
rect 5858 65852 5922 65856
rect 5858 65796 5862 65852
rect 5862 65796 5918 65852
rect 5918 65796 5922 65852
rect 5858 65792 5922 65796
rect 10285 65852 10349 65856
rect 10285 65796 10289 65852
rect 10289 65796 10345 65852
rect 10345 65796 10349 65852
rect 10285 65792 10349 65796
rect 10365 65852 10429 65856
rect 10365 65796 10369 65852
rect 10369 65796 10425 65852
rect 10425 65796 10429 65852
rect 10365 65792 10429 65796
rect 10445 65852 10509 65856
rect 10445 65796 10449 65852
rect 10449 65796 10505 65852
rect 10505 65796 10509 65852
rect 10445 65792 10509 65796
rect 10525 65852 10589 65856
rect 10525 65796 10529 65852
rect 10529 65796 10585 65852
rect 10585 65796 10589 65852
rect 10525 65792 10589 65796
rect 3285 65308 3349 65312
rect 3285 65252 3289 65308
rect 3289 65252 3345 65308
rect 3345 65252 3349 65308
rect 3285 65248 3349 65252
rect 3365 65308 3429 65312
rect 3365 65252 3369 65308
rect 3369 65252 3425 65308
rect 3425 65252 3429 65308
rect 3365 65248 3429 65252
rect 3445 65308 3509 65312
rect 3445 65252 3449 65308
rect 3449 65252 3505 65308
rect 3505 65252 3509 65308
rect 3445 65248 3509 65252
rect 3525 65308 3589 65312
rect 3525 65252 3529 65308
rect 3529 65252 3585 65308
rect 3585 65252 3589 65308
rect 3525 65248 3589 65252
rect 7952 65308 8016 65312
rect 7952 65252 7956 65308
rect 7956 65252 8012 65308
rect 8012 65252 8016 65308
rect 7952 65248 8016 65252
rect 8032 65308 8096 65312
rect 8032 65252 8036 65308
rect 8036 65252 8092 65308
rect 8092 65252 8096 65308
rect 8032 65248 8096 65252
rect 8112 65308 8176 65312
rect 8112 65252 8116 65308
rect 8116 65252 8172 65308
rect 8172 65252 8176 65308
rect 8112 65248 8176 65252
rect 8192 65308 8256 65312
rect 8192 65252 8196 65308
rect 8196 65252 8252 65308
rect 8252 65252 8256 65308
rect 8192 65248 8256 65252
rect 5618 64764 5682 64768
rect 5618 64708 5622 64764
rect 5622 64708 5678 64764
rect 5678 64708 5682 64764
rect 5618 64704 5682 64708
rect 5698 64764 5762 64768
rect 5698 64708 5702 64764
rect 5702 64708 5758 64764
rect 5758 64708 5762 64764
rect 5698 64704 5762 64708
rect 5778 64764 5842 64768
rect 5778 64708 5782 64764
rect 5782 64708 5838 64764
rect 5838 64708 5842 64764
rect 5778 64704 5842 64708
rect 5858 64764 5922 64768
rect 5858 64708 5862 64764
rect 5862 64708 5918 64764
rect 5918 64708 5922 64764
rect 5858 64704 5922 64708
rect 10285 64764 10349 64768
rect 10285 64708 10289 64764
rect 10289 64708 10345 64764
rect 10345 64708 10349 64764
rect 10285 64704 10349 64708
rect 10365 64764 10429 64768
rect 10365 64708 10369 64764
rect 10369 64708 10425 64764
rect 10425 64708 10429 64764
rect 10365 64704 10429 64708
rect 10445 64764 10509 64768
rect 10445 64708 10449 64764
rect 10449 64708 10505 64764
rect 10505 64708 10509 64764
rect 10445 64704 10509 64708
rect 10525 64764 10589 64768
rect 10525 64708 10529 64764
rect 10529 64708 10585 64764
rect 10585 64708 10589 64764
rect 10525 64704 10589 64708
rect 3285 64220 3349 64224
rect 3285 64164 3289 64220
rect 3289 64164 3345 64220
rect 3345 64164 3349 64220
rect 3285 64160 3349 64164
rect 3365 64220 3429 64224
rect 3365 64164 3369 64220
rect 3369 64164 3425 64220
rect 3425 64164 3429 64220
rect 3365 64160 3429 64164
rect 3445 64220 3509 64224
rect 3445 64164 3449 64220
rect 3449 64164 3505 64220
rect 3505 64164 3509 64220
rect 3445 64160 3509 64164
rect 3525 64220 3589 64224
rect 3525 64164 3529 64220
rect 3529 64164 3585 64220
rect 3585 64164 3589 64220
rect 3525 64160 3589 64164
rect 7952 64220 8016 64224
rect 7952 64164 7956 64220
rect 7956 64164 8012 64220
rect 8012 64164 8016 64220
rect 7952 64160 8016 64164
rect 8032 64220 8096 64224
rect 8032 64164 8036 64220
rect 8036 64164 8092 64220
rect 8092 64164 8096 64220
rect 8032 64160 8096 64164
rect 8112 64220 8176 64224
rect 8112 64164 8116 64220
rect 8116 64164 8172 64220
rect 8172 64164 8176 64220
rect 8112 64160 8176 64164
rect 8192 64220 8256 64224
rect 8192 64164 8196 64220
rect 8196 64164 8252 64220
rect 8252 64164 8256 64220
rect 8192 64160 8256 64164
rect 5618 63676 5682 63680
rect 5618 63620 5622 63676
rect 5622 63620 5678 63676
rect 5678 63620 5682 63676
rect 5618 63616 5682 63620
rect 5698 63676 5762 63680
rect 5698 63620 5702 63676
rect 5702 63620 5758 63676
rect 5758 63620 5762 63676
rect 5698 63616 5762 63620
rect 5778 63676 5842 63680
rect 5778 63620 5782 63676
rect 5782 63620 5838 63676
rect 5838 63620 5842 63676
rect 5778 63616 5842 63620
rect 5858 63676 5922 63680
rect 5858 63620 5862 63676
rect 5862 63620 5918 63676
rect 5918 63620 5922 63676
rect 5858 63616 5922 63620
rect 10285 63676 10349 63680
rect 10285 63620 10289 63676
rect 10289 63620 10345 63676
rect 10345 63620 10349 63676
rect 10285 63616 10349 63620
rect 10365 63676 10429 63680
rect 10365 63620 10369 63676
rect 10369 63620 10425 63676
rect 10425 63620 10429 63676
rect 10365 63616 10429 63620
rect 10445 63676 10509 63680
rect 10445 63620 10449 63676
rect 10449 63620 10505 63676
rect 10505 63620 10509 63676
rect 10445 63616 10509 63620
rect 10525 63676 10589 63680
rect 10525 63620 10529 63676
rect 10529 63620 10585 63676
rect 10585 63620 10589 63676
rect 10525 63616 10589 63620
rect 3285 63132 3349 63136
rect 3285 63076 3289 63132
rect 3289 63076 3345 63132
rect 3345 63076 3349 63132
rect 3285 63072 3349 63076
rect 3365 63132 3429 63136
rect 3365 63076 3369 63132
rect 3369 63076 3425 63132
rect 3425 63076 3429 63132
rect 3365 63072 3429 63076
rect 3445 63132 3509 63136
rect 3445 63076 3449 63132
rect 3449 63076 3505 63132
rect 3505 63076 3509 63132
rect 3445 63072 3509 63076
rect 3525 63132 3589 63136
rect 3525 63076 3529 63132
rect 3529 63076 3585 63132
rect 3585 63076 3589 63132
rect 3525 63072 3589 63076
rect 7952 63132 8016 63136
rect 7952 63076 7956 63132
rect 7956 63076 8012 63132
rect 8012 63076 8016 63132
rect 7952 63072 8016 63076
rect 8032 63132 8096 63136
rect 8032 63076 8036 63132
rect 8036 63076 8092 63132
rect 8092 63076 8096 63132
rect 8032 63072 8096 63076
rect 8112 63132 8176 63136
rect 8112 63076 8116 63132
rect 8116 63076 8172 63132
rect 8172 63076 8176 63132
rect 8112 63072 8176 63076
rect 8192 63132 8256 63136
rect 8192 63076 8196 63132
rect 8196 63076 8252 63132
rect 8252 63076 8256 63132
rect 8192 63072 8256 63076
rect 5618 62588 5682 62592
rect 5618 62532 5622 62588
rect 5622 62532 5678 62588
rect 5678 62532 5682 62588
rect 5618 62528 5682 62532
rect 5698 62588 5762 62592
rect 5698 62532 5702 62588
rect 5702 62532 5758 62588
rect 5758 62532 5762 62588
rect 5698 62528 5762 62532
rect 5778 62588 5842 62592
rect 5778 62532 5782 62588
rect 5782 62532 5838 62588
rect 5838 62532 5842 62588
rect 5778 62528 5842 62532
rect 5858 62588 5922 62592
rect 5858 62532 5862 62588
rect 5862 62532 5918 62588
rect 5918 62532 5922 62588
rect 5858 62528 5922 62532
rect 10285 62588 10349 62592
rect 10285 62532 10289 62588
rect 10289 62532 10345 62588
rect 10345 62532 10349 62588
rect 10285 62528 10349 62532
rect 10365 62588 10429 62592
rect 10365 62532 10369 62588
rect 10369 62532 10425 62588
rect 10425 62532 10429 62588
rect 10365 62528 10429 62532
rect 10445 62588 10509 62592
rect 10445 62532 10449 62588
rect 10449 62532 10505 62588
rect 10505 62532 10509 62588
rect 10445 62528 10509 62532
rect 10525 62588 10589 62592
rect 10525 62532 10529 62588
rect 10529 62532 10585 62588
rect 10585 62532 10589 62588
rect 10525 62528 10589 62532
rect 3285 62044 3349 62048
rect 3285 61988 3289 62044
rect 3289 61988 3345 62044
rect 3345 61988 3349 62044
rect 3285 61984 3349 61988
rect 3365 62044 3429 62048
rect 3365 61988 3369 62044
rect 3369 61988 3425 62044
rect 3425 61988 3429 62044
rect 3365 61984 3429 61988
rect 3445 62044 3509 62048
rect 3445 61988 3449 62044
rect 3449 61988 3505 62044
rect 3505 61988 3509 62044
rect 3445 61984 3509 61988
rect 3525 62044 3589 62048
rect 3525 61988 3529 62044
rect 3529 61988 3585 62044
rect 3585 61988 3589 62044
rect 3525 61984 3589 61988
rect 7952 62044 8016 62048
rect 7952 61988 7956 62044
rect 7956 61988 8012 62044
rect 8012 61988 8016 62044
rect 7952 61984 8016 61988
rect 8032 62044 8096 62048
rect 8032 61988 8036 62044
rect 8036 61988 8092 62044
rect 8092 61988 8096 62044
rect 8032 61984 8096 61988
rect 8112 62044 8176 62048
rect 8112 61988 8116 62044
rect 8116 61988 8172 62044
rect 8172 61988 8176 62044
rect 8112 61984 8176 61988
rect 8192 62044 8256 62048
rect 8192 61988 8196 62044
rect 8196 61988 8252 62044
rect 8252 61988 8256 62044
rect 8192 61984 8256 61988
rect 5618 61500 5682 61504
rect 5618 61444 5622 61500
rect 5622 61444 5678 61500
rect 5678 61444 5682 61500
rect 5618 61440 5682 61444
rect 5698 61500 5762 61504
rect 5698 61444 5702 61500
rect 5702 61444 5758 61500
rect 5758 61444 5762 61500
rect 5698 61440 5762 61444
rect 5778 61500 5842 61504
rect 5778 61444 5782 61500
rect 5782 61444 5838 61500
rect 5838 61444 5842 61500
rect 5778 61440 5842 61444
rect 5858 61500 5922 61504
rect 5858 61444 5862 61500
rect 5862 61444 5918 61500
rect 5918 61444 5922 61500
rect 5858 61440 5922 61444
rect 10285 61500 10349 61504
rect 10285 61444 10289 61500
rect 10289 61444 10345 61500
rect 10345 61444 10349 61500
rect 10285 61440 10349 61444
rect 10365 61500 10429 61504
rect 10365 61444 10369 61500
rect 10369 61444 10425 61500
rect 10425 61444 10429 61500
rect 10365 61440 10429 61444
rect 10445 61500 10509 61504
rect 10445 61444 10449 61500
rect 10449 61444 10505 61500
rect 10505 61444 10509 61500
rect 10445 61440 10509 61444
rect 10525 61500 10589 61504
rect 10525 61444 10529 61500
rect 10529 61444 10585 61500
rect 10585 61444 10589 61500
rect 10525 61440 10589 61444
rect 3285 60956 3349 60960
rect 3285 60900 3289 60956
rect 3289 60900 3345 60956
rect 3345 60900 3349 60956
rect 3285 60896 3349 60900
rect 3365 60956 3429 60960
rect 3365 60900 3369 60956
rect 3369 60900 3425 60956
rect 3425 60900 3429 60956
rect 3365 60896 3429 60900
rect 3445 60956 3509 60960
rect 3445 60900 3449 60956
rect 3449 60900 3505 60956
rect 3505 60900 3509 60956
rect 3445 60896 3509 60900
rect 3525 60956 3589 60960
rect 3525 60900 3529 60956
rect 3529 60900 3585 60956
rect 3585 60900 3589 60956
rect 3525 60896 3589 60900
rect 7952 60956 8016 60960
rect 7952 60900 7956 60956
rect 7956 60900 8012 60956
rect 8012 60900 8016 60956
rect 7952 60896 8016 60900
rect 8032 60956 8096 60960
rect 8032 60900 8036 60956
rect 8036 60900 8092 60956
rect 8092 60900 8096 60956
rect 8032 60896 8096 60900
rect 8112 60956 8176 60960
rect 8112 60900 8116 60956
rect 8116 60900 8172 60956
rect 8172 60900 8176 60956
rect 8112 60896 8176 60900
rect 8192 60956 8256 60960
rect 8192 60900 8196 60956
rect 8196 60900 8252 60956
rect 8252 60900 8256 60956
rect 8192 60896 8256 60900
rect 5618 60412 5682 60416
rect 5618 60356 5622 60412
rect 5622 60356 5678 60412
rect 5678 60356 5682 60412
rect 5618 60352 5682 60356
rect 5698 60412 5762 60416
rect 5698 60356 5702 60412
rect 5702 60356 5758 60412
rect 5758 60356 5762 60412
rect 5698 60352 5762 60356
rect 5778 60412 5842 60416
rect 5778 60356 5782 60412
rect 5782 60356 5838 60412
rect 5838 60356 5842 60412
rect 5778 60352 5842 60356
rect 5858 60412 5922 60416
rect 5858 60356 5862 60412
rect 5862 60356 5918 60412
rect 5918 60356 5922 60412
rect 5858 60352 5922 60356
rect 10285 60412 10349 60416
rect 10285 60356 10289 60412
rect 10289 60356 10345 60412
rect 10345 60356 10349 60412
rect 10285 60352 10349 60356
rect 10365 60412 10429 60416
rect 10365 60356 10369 60412
rect 10369 60356 10425 60412
rect 10425 60356 10429 60412
rect 10365 60352 10429 60356
rect 10445 60412 10509 60416
rect 10445 60356 10449 60412
rect 10449 60356 10505 60412
rect 10505 60356 10509 60412
rect 10445 60352 10509 60356
rect 10525 60412 10589 60416
rect 10525 60356 10529 60412
rect 10529 60356 10585 60412
rect 10585 60356 10589 60412
rect 10525 60352 10589 60356
rect 3285 59868 3349 59872
rect 3285 59812 3289 59868
rect 3289 59812 3345 59868
rect 3345 59812 3349 59868
rect 3285 59808 3349 59812
rect 3365 59868 3429 59872
rect 3365 59812 3369 59868
rect 3369 59812 3425 59868
rect 3425 59812 3429 59868
rect 3365 59808 3429 59812
rect 3445 59868 3509 59872
rect 3445 59812 3449 59868
rect 3449 59812 3505 59868
rect 3505 59812 3509 59868
rect 3445 59808 3509 59812
rect 3525 59868 3589 59872
rect 3525 59812 3529 59868
rect 3529 59812 3585 59868
rect 3585 59812 3589 59868
rect 3525 59808 3589 59812
rect 7952 59868 8016 59872
rect 7952 59812 7956 59868
rect 7956 59812 8012 59868
rect 8012 59812 8016 59868
rect 7952 59808 8016 59812
rect 8032 59868 8096 59872
rect 8032 59812 8036 59868
rect 8036 59812 8092 59868
rect 8092 59812 8096 59868
rect 8032 59808 8096 59812
rect 8112 59868 8176 59872
rect 8112 59812 8116 59868
rect 8116 59812 8172 59868
rect 8172 59812 8176 59868
rect 8112 59808 8176 59812
rect 8192 59868 8256 59872
rect 8192 59812 8196 59868
rect 8196 59812 8252 59868
rect 8252 59812 8256 59868
rect 8192 59808 8256 59812
rect 5618 59324 5682 59328
rect 5618 59268 5622 59324
rect 5622 59268 5678 59324
rect 5678 59268 5682 59324
rect 5618 59264 5682 59268
rect 5698 59324 5762 59328
rect 5698 59268 5702 59324
rect 5702 59268 5758 59324
rect 5758 59268 5762 59324
rect 5698 59264 5762 59268
rect 5778 59324 5842 59328
rect 5778 59268 5782 59324
rect 5782 59268 5838 59324
rect 5838 59268 5842 59324
rect 5778 59264 5842 59268
rect 5858 59324 5922 59328
rect 5858 59268 5862 59324
rect 5862 59268 5918 59324
rect 5918 59268 5922 59324
rect 5858 59264 5922 59268
rect 10285 59324 10349 59328
rect 10285 59268 10289 59324
rect 10289 59268 10345 59324
rect 10345 59268 10349 59324
rect 10285 59264 10349 59268
rect 10365 59324 10429 59328
rect 10365 59268 10369 59324
rect 10369 59268 10425 59324
rect 10425 59268 10429 59324
rect 10365 59264 10429 59268
rect 10445 59324 10509 59328
rect 10445 59268 10449 59324
rect 10449 59268 10505 59324
rect 10505 59268 10509 59324
rect 10445 59264 10509 59268
rect 10525 59324 10589 59328
rect 10525 59268 10529 59324
rect 10529 59268 10585 59324
rect 10585 59268 10589 59324
rect 10525 59264 10589 59268
rect 3285 58780 3349 58784
rect 3285 58724 3289 58780
rect 3289 58724 3345 58780
rect 3345 58724 3349 58780
rect 3285 58720 3349 58724
rect 3365 58780 3429 58784
rect 3365 58724 3369 58780
rect 3369 58724 3425 58780
rect 3425 58724 3429 58780
rect 3365 58720 3429 58724
rect 3445 58780 3509 58784
rect 3445 58724 3449 58780
rect 3449 58724 3505 58780
rect 3505 58724 3509 58780
rect 3445 58720 3509 58724
rect 3525 58780 3589 58784
rect 3525 58724 3529 58780
rect 3529 58724 3585 58780
rect 3585 58724 3589 58780
rect 3525 58720 3589 58724
rect 7952 58780 8016 58784
rect 7952 58724 7956 58780
rect 7956 58724 8012 58780
rect 8012 58724 8016 58780
rect 7952 58720 8016 58724
rect 8032 58780 8096 58784
rect 8032 58724 8036 58780
rect 8036 58724 8092 58780
rect 8092 58724 8096 58780
rect 8032 58720 8096 58724
rect 8112 58780 8176 58784
rect 8112 58724 8116 58780
rect 8116 58724 8172 58780
rect 8172 58724 8176 58780
rect 8112 58720 8176 58724
rect 8192 58780 8256 58784
rect 8192 58724 8196 58780
rect 8196 58724 8252 58780
rect 8252 58724 8256 58780
rect 8192 58720 8256 58724
rect 5618 58236 5682 58240
rect 5618 58180 5622 58236
rect 5622 58180 5678 58236
rect 5678 58180 5682 58236
rect 5618 58176 5682 58180
rect 5698 58236 5762 58240
rect 5698 58180 5702 58236
rect 5702 58180 5758 58236
rect 5758 58180 5762 58236
rect 5698 58176 5762 58180
rect 5778 58236 5842 58240
rect 5778 58180 5782 58236
rect 5782 58180 5838 58236
rect 5838 58180 5842 58236
rect 5778 58176 5842 58180
rect 5858 58236 5922 58240
rect 5858 58180 5862 58236
rect 5862 58180 5918 58236
rect 5918 58180 5922 58236
rect 5858 58176 5922 58180
rect 10285 58236 10349 58240
rect 10285 58180 10289 58236
rect 10289 58180 10345 58236
rect 10345 58180 10349 58236
rect 10285 58176 10349 58180
rect 10365 58236 10429 58240
rect 10365 58180 10369 58236
rect 10369 58180 10425 58236
rect 10425 58180 10429 58236
rect 10365 58176 10429 58180
rect 10445 58236 10509 58240
rect 10445 58180 10449 58236
rect 10449 58180 10505 58236
rect 10505 58180 10509 58236
rect 10445 58176 10509 58180
rect 10525 58236 10589 58240
rect 10525 58180 10529 58236
rect 10529 58180 10585 58236
rect 10585 58180 10589 58236
rect 10525 58176 10589 58180
rect 3285 57692 3349 57696
rect 3285 57636 3289 57692
rect 3289 57636 3345 57692
rect 3345 57636 3349 57692
rect 3285 57632 3349 57636
rect 3365 57692 3429 57696
rect 3365 57636 3369 57692
rect 3369 57636 3425 57692
rect 3425 57636 3429 57692
rect 3365 57632 3429 57636
rect 3445 57692 3509 57696
rect 3445 57636 3449 57692
rect 3449 57636 3505 57692
rect 3505 57636 3509 57692
rect 3445 57632 3509 57636
rect 3525 57692 3589 57696
rect 3525 57636 3529 57692
rect 3529 57636 3585 57692
rect 3585 57636 3589 57692
rect 3525 57632 3589 57636
rect 7952 57692 8016 57696
rect 7952 57636 7956 57692
rect 7956 57636 8012 57692
rect 8012 57636 8016 57692
rect 7952 57632 8016 57636
rect 8032 57692 8096 57696
rect 8032 57636 8036 57692
rect 8036 57636 8092 57692
rect 8092 57636 8096 57692
rect 8032 57632 8096 57636
rect 8112 57692 8176 57696
rect 8112 57636 8116 57692
rect 8116 57636 8172 57692
rect 8172 57636 8176 57692
rect 8112 57632 8176 57636
rect 8192 57692 8256 57696
rect 8192 57636 8196 57692
rect 8196 57636 8252 57692
rect 8252 57636 8256 57692
rect 8192 57632 8256 57636
rect 5618 57148 5682 57152
rect 5618 57092 5622 57148
rect 5622 57092 5678 57148
rect 5678 57092 5682 57148
rect 5618 57088 5682 57092
rect 5698 57148 5762 57152
rect 5698 57092 5702 57148
rect 5702 57092 5758 57148
rect 5758 57092 5762 57148
rect 5698 57088 5762 57092
rect 5778 57148 5842 57152
rect 5778 57092 5782 57148
rect 5782 57092 5838 57148
rect 5838 57092 5842 57148
rect 5778 57088 5842 57092
rect 5858 57148 5922 57152
rect 5858 57092 5862 57148
rect 5862 57092 5918 57148
rect 5918 57092 5922 57148
rect 5858 57088 5922 57092
rect 10285 57148 10349 57152
rect 10285 57092 10289 57148
rect 10289 57092 10345 57148
rect 10345 57092 10349 57148
rect 10285 57088 10349 57092
rect 10365 57148 10429 57152
rect 10365 57092 10369 57148
rect 10369 57092 10425 57148
rect 10425 57092 10429 57148
rect 10365 57088 10429 57092
rect 10445 57148 10509 57152
rect 10445 57092 10449 57148
rect 10449 57092 10505 57148
rect 10505 57092 10509 57148
rect 10445 57088 10509 57092
rect 10525 57148 10589 57152
rect 10525 57092 10529 57148
rect 10529 57092 10585 57148
rect 10585 57092 10589 57148
rect 10525 57088 10589 57092
rect 3285 56604 3349 56608
rect 3285 56548 3289 56604
rect 3289 56548 3345 56604
rect 3345 56548 3349 56604
rect 3285 56544 3349 56548
rect 3365 56604 3429 56608
rect 3365 56548 3369 56604
rect 3369 56548 3425 56604
rect 3425 56548 3429 56604
rect 3365 56544 3429 56548
rect 3445 56604 3509 56608
rect 3445 56548 3449 56604
rect 3449 56548 3505 56604
rect 3505 56548 3509 56604
rect 3445 56544 3509 56548
rect 3525 56604 3589 56608
rect 3525 56548 3529 56604
rect 3529 56548 3585 56604
rect 3585 56548 3589 56604
rect 3525 56544 3589 56548
rect 7952 56604 8016 56608
rect 7952 56548 7956 56604
rect 7956 56548 8012 56604
rect 8012 56548 8016 56604
rect 7952 56544 8016 56548
rect 8032 56604 8096 56608
rect 8032 56548 8036 56604
rect 8036 56548 8092 56604
rect 8092 56548 8096 56604
rect 8032 56544 8096 56548
rect 8112 56604 8176 56608
rect 8112 56548 8116 56604
rect 8116 56548 8172 56604
rect 8172 56548 8176 56604
rect 8112 56544 8176 56548
rect 8192 56604 8256 56608
rect 8192 56548 8196 56604
rect 8196 56548 8252 56604
rect 8252 56548 8256 56604
rect 8192 56544 8256 56548
rect 5618 56060 5682 56064
rect 5618 56004 5622 56060
rect 5622 56004 5678 56060
rect 5678 56004 5682 56060
rect 5618 56000 5682 56004
rect 5698 56060 5762 56064
rect 5698 56004 5702 56060
rect 5702 56004 5758 56060
rect 5758 56004 5762 56060
rect 5698 56000 5762 56004
rect 5778 56060 5842 56064
rect 5778 56004 5782 56060
rect 5782 56004 5838 56060
rect 5838 56004 5842 56060
rect 5778 56000 5842 56004
rect 5858 56060 5922 56064
rect 5858 56004 5862 56060
rect 5862 56004 5918 56060
rect 5918 56004 5922 56060
rect 5858 56000 5922 56004
rect 10285 56060 10349 56064
rect 10285 56004 10289 56060
rect 10289 56004 10345 56060
rect 10345 56004 10349 56060
rect 10285 56000 10349 56004
rect 10365 56060 10429 56064
rect 10365 56004 10369 56060
rect 10369 56004 10425 56060
rect 10425 56004 10429 56060
rect 10365 56000 10429 56004
rect 10445 56060 10509 56064
rect 10445 56004 10449 56060
rect 10449 56004 10505 56060
rect 10505 56004 10509 56060
rect 10445 56000 10509 56004
rect 10525 56060 10589 56064
rect 10525 56004 10529 56060
rect 10529 56004 10585 56060
rect 10585 56004 10589 56060
rect 10525 56000 10589 56004
rect 3285 55516 3349 55520
rect 3285 55460 3289 55516
rect 3289 55460 3345 55516
rect 3345 55460 3349 55516
rect 3285 55456 3349 55460
rect 3365 55516 3429 55520
rect 3365 55460 3369 55516
rect 3369 55460 3425 55516
rect 3425 55460 3429 55516
rect 3365 55456 3429 55460
rect 3445 55516 3509 55520
rect 3445 55460 3449 55516
rect 3449 55460 3505 55516
rect 3505 55460 3509 55516
rect 3445 55456 3509 55460
rect 3525 55516 3589 55520
rect 3525 55460 3529 55516
rect 3529 55460 3585 55516
rect 3585 55460 3589 55516
rect 3525 55456 3589 55460
rect 7952 55516 8016 55520
rect 7952 55460 7956 55516
rect 7956 55460 8012 55516
rect 8012 55460 8016 55516
rect 7952 55456 8016 55460
rect 8032 55516 8096 55520
rect 8032 55460 8036 55516
rect 8036 55460 8092 55516
rect 8092 55460 8096 55516
rect 8032 55456 8096 55460
rect 8112 55516 8176 55520
rect 8112 55460 8116 55516
rect 8116 55460 8172 55516
rect 8172 55460 8176 55516
rect 8112 55456 8176 55460
rect 8192 55516 8256 55520
rect 8192 55460 8196 55516
rect 8196 55460 8252 55516
rect 8252 55460 8256 55516
rect 8192 55456 8256 55460
rect 5618 54972 5682 54976
rect 5618 54916 5622 54972
rect 5622 54916 5678 54972
rect 5678 54916 5682 54972
rect 5618 54912 5682 54916
rect 5698 54972 5762 54976
rect 5698 54916 5702 54972
rect 5702 54916 5758 54972
rect 5758 54916 5762 54972
rect 5698 54912 5762 54916
rect 5778 54972 5842 54976
rect 5778 54916 5782 54972
rect 5782 54916 5838 54972
rect 5838 54916 5842 54972
rect 5778 54912 5842 54916
rect 5858 54972 5922 54976
rect 5858 54916 5862 54972
rect 5862 54916 5918 54972
rect 5918 54916 5922 54972
rect 5858 54912 5922 54916
rect 10285 54972 10349 54976
rect 10285 54916 10289 54972
rect 10289 54916 10345 54972
rect 10345 54916 10349 54972
rect 10285 54912 10349 54916
rect 10365 54972 10429 54976
rect 10365 54916 10369 54972
rect 10369 54916 10425 54972
rect 10425 54916 10429 54972
rect 10365 54912 10429 54916
rect 10445 54972 10509 54976
rect 10445 54916 10449 54972
rect 10449 54916 10505 54972
rect 10505 54916 10509 54972
rect 10445 54912 10509 54916
rect 10525 54972 10589 54976
rect 10525 54916 10529 54972
rect 10529 54916 10585 54972
rect 10585 54916 10589 54972
rect 10525 54912 10589 54916
rect 3285 54428 3349 54432
rect 3285 54372 3289 54428
rect 3289 54372 3345 54428
rect 3345 54372 3349 54428
rect 3285 54368 3349 54372
rect 3365 54428 3429 54432
rect 3365 54372 3369 54428
rect 3369 54372 3425 54428
rect 3425 54372 3429 54428
rect 3365 54368 3429 54372
rect 3445 54428 3509 54432
rect 3445 54372 3449 54428
rect 3449 54372 3505 54428
rect 3505 54372 3509 54428
rect 3445 54368 3509 54372
rect 3525 54428 3589 54432
rect 3525 54372 3529 54428
rect 3529 54372 3585 54428
rect 3585 54372 3589 54428
rect 3525 54368 3589 54372
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 5618 53884 5682 53888
rect 5618 53828 5622 53884
rect 5622 53828 5678 53884
rect 5678 53828 5682 53884
rect 5618 53824 5682 53828
rect 5698 53884 5762 53888
rect 5698 53828 5702 53884
rect 5702 53828 5758 53884
rect 5758 53828 5762 53884
rect 5698 53824 5762 53828
rect 5778 53884 5842 53888
rect 5778 53828 5782 53884
rect 5782 53828 5838 53884
rect 5838 53828 5842 53884
rect 5778 53824 5842 53828
rect 5858 53884 5922 53888
rect 5858 53828 5862 53884
rect 5862 53828 5918 53884
rect 5918 53828 5922 53884
rect 5858 53824 5922 53828
rect 10285 53884 10349 53888
rect 10285 53828 10289 53884
rect 10289 53828 10345 53884
rect 10345 53828 10349 53884
rect 10285 53824 10349 53828
rect 10365 53884 10429 53888
rect 10365 53828 10369 53884
rect 10369 53828 10425 53884
rect 10425 53828 10429 53884
rect 10365 53824 10429 53828
rect 10445 53884 10509 53888
rect 10445 53828 10449 53884
rect 10449 53828 10505 53884
rect 10505 53828 10509 53884
rect 10445 53824 10509 53828
rect 10525 53884 10589 53888
rect 10525 53828 10529 53884
rect 10529 53828 10585 53884
rect 10585 53828 10589 53884
rect 10525 53824 10589 53828
rect 3285 53340 3349 53344
rect 3285 53284 3289 53340
rect 3289 53284 3345 53340
rect 3345 53284 3349 53340
rect 3285 53280 3349 53284
rect 3365 53340 3429 53344
rect 3365 53284 3369 53340
rect 3369 53284 3425 53340
rect 3425 53284 3429 53340
rect 3365 53280 3429 53284
rect 3445 53340 3509 53344
rect 3445 53284 3449 53340
rect 3449 53284 3505 53340
rect 3505 53284 3509 53340
rect 3445 53280 3509 53284
rect 3525 53340 3589 53344
rect 3525 53284 3529 53340
rect 3529 53284 3585 53340
rect 3585 53284 3589 53340
rect 3525 53280 3589 53284
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 5618 52796 5682 52800
rect 5618 52740 5622 52796
rect 5622 52740 5678 52796
rect 5678 52740 5682 52796
rect 5618 52736 5682 52740
rect 5698 52796 5762 52800
rect 5698 52740 5702 52796
rect 5702 52740 5758 52796
rect 5758 52740 5762 52796
rect 5698 52736 5762 52740
rect 5778 52796 5842 52800
rect 5778 52740 5782 52796
rect 5782 52740 5838 52796
rect 5838 52740 5842 52796
rect 5778 52736 5842 52740
rect 5858 52796 5922 52800
rect 5858 52740 5862 52796
rect 5862 52740 5918 52796
rect 5918 52740 5922 52796
rect 5858 52736 5922 52740
rect 10285 52796 10349 52800
rect 10285 52740 10289 52796
rect 10289 52740 10345 52796
rect 10345 52740 10349 52796
rect 10285 52736 10349 52740
rect 10365 52796 10429 52800
rect 10365 52740 10369 52796
rect 10369 52740 10425 52796
rect 10425 52740 10429 52796
rect 10365 52736 10429 52740
rect 10445 52796 10509 52800
rect 10445 52740 10449 52796
rect 10449 52740 10505 52796
rect 10505 52740 10509 52796
rect 10445 52736 10509 52740
rect 10525 52796 10589 52800
rect 10525 52740 10529 52796
rect 10529 52740 10585 52796
rect 10585 52740 10589 52796
rect 10525 52736 10589 52740
rect 3285 52252 3349 52256
rect 3285 52196 3289 52252
rect 3289 52196 3345 52252
rect 3345 52196 3349 52252
rect 3285 52192 3349 52196
rect 3365 52252 3429 52256
rect 3365 52196 3369 52252
rect 3369 52196 3425 52252
rect 3425 52196 3429 52252
rect 3365 52192 3429 52196
rect 3445 52252 3509 52256
rect 3445 52196 3449 52252
rect 3449 52196 3505 52252
rect 3505 52196 3509 52252
rect 3445 52192 3509 52196
rect 3525 52252 3589 52256
rect 3525 52196 3529 52252
rect 3529 52196 3585 52252
rect 3585 52196 3589 52252
rect 3525 52192 3589 52196
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 5618 51708 5682 51712
rect 5618 51652 5622 51708
rect 5622 51652 5678 51708
rect 5678 51652 5682 51708
rect 5618 51648 5682 51652
rect 5698 51708 5762 51712
rect 5698 51652 5702 51708
rect 5702 51652 5758 51708
rect 5758 51652 5762 51708
rect 5698 51648 5762 51652
rect 5778 51708 5842 51712
rect 5778 51652 5782 51708
rect 5782 51652 5838 51708
rect 5838 51652 5842 51708
rect 5778 51648 5842 51652
rect 5858 51708 5922 51712
rect 5858 51652 5862 51708
rect 5862 51652 5918 51708
rect 5918 51652 5922 51708
rect 5858 51648 5922 51652
rect 10285 51708 10349 51712
rect 10285 51652 10289 51708
rect 10289 51652 10345 51708
rect 10345 51652 10349 51708
rect 10285 51648 10349 51652
rect 10365 51708 10429 51712
rect 10365 51652 10369 51708
rect 10369 51652 10425 51708
rect 10425 51652 10429 51708
rect 10365 51648 10429 51652
rect 10445 51708 10509 51712
rect 10445 51652 10449 51708
rect 10449 51652 10505 51708
rect 10505 51652 10509 51708
rect 10445 51648 10509 51652
rect 10525 51708 10589 51712
rect 10525 51652 10529 51708
rect 10529 51652 10585 51708
rect 10585 51652 10589 51708
rect 10525 51648 10589 51652
rect 3285 51164 3349 51168
rect 3285 51108 3289 51164
rect 3289 51108 3345 51164
rect 3345 51108 3349 51164
rect 3285 51104 3349 51108
rect 3365 51164 3429 51168
rect 3365 51108 3369 51164
rect 3369 51108 3425 51164
rect 3425 51108 3429 51164
rect 3365 51104 3429 51108
rect 3445 51164 3509 51168
rect 3445 51108 3449 51164
rect 3449 51108 3505 51164
rect 3505 51108 3509 51164
rect 3445 51104 3509 51108
rect 3525 51164 3589 51168
rect 3525 51108 3529 51164
rect 3529 51108 3585 51164
rect 3585 51108 3589 51164
rect 3525 51104 3589 51108
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 5618 50620 5682 50624
rect 5618 50564 5622 50620
rect 5622 50564 5678 50620
rect 5678 50564 5682 50620
rect 5618 50560 5682 50564
rect 5698 50620 5762 50624
rect 5698 50564 5702 50620
rect 5702 50564 5758 50620
rect 5758 50564 5762 50620
rect 5698 50560 5762 50564
rect 5778 50620 5842 50624
rect 5778 50564 5782 50620
rect 5782 50564 5838 50620
rect 5838 50564 5842 50620
rect 5778 50560 5842 50564
rect 5858 50620 5922 50624
rect 5858 50564 5862 50620
rect 5862 50564 5918 50620
rect 5918 50564 5922 50620
rect 5858 50560 5922 50564
rect 10285 50620 10349 50624
rect 10285 50564 10289 50620
rect 10289 50564 10345 50620
rect 10345 50564 10349 50620
rect 10285 50560 10349 50564
rect 10365 50620 10429 50624
rect 10365 50564 10369 50620
rect 10369 50564 10425 50620
rect 10425 50564 10429 50620
rect 10365 50560 10429 50564
rect 10445 50620 10509 50624
rect 10445 50564 10449 50620
rect 10449 50564 10505 50620
rect 10505 50564 10509 50620
rect 10445 50560 10509 50564
rect 10525 50620 10589 50624
rect 10525 50564 10529 50620
rect 10529 50564 10585 50620
rect 10585 50564 10589 50620
rect 10525 50560 10589 50564
rect 3285 50076 3349 50080
rect 3285 50020 3289 50076
rect 3289 50020 3345 50076
rect 3345 50020 3349 50076
rect 3285 50016 3349 50020
rect 3365 50076 3429 50080
rect 3365 50020 3369 50076
rect 3369 50020 3425 50076
rect 3425 50020 3429 50076
rect 3365 50016 3429 50020
rect 3445 50076 3509 50080
rect 3445 50020 3449 50076
rect 3449 50020 3505 50076
rect 3505 50020 3509 50076
rect 3445 50016 3509 50020
rect 3525 50076 3589 50080
rect 3525 50020 3529 50076
rect 3529 50020 3585 50076
rect 3585 50020 3589 50076
rect 3525 50016 3589 50020
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 5618 49532 5682 49536
rect 5618 49476 5622 49532
rect 5622 49476 5678 49532
rect 5678 49476 5682 49532
rect 5618 49472 5682 49476
rect 5698 49532 5762 49536
rect 5698 49476 5702 49532
rect 5702 49476 5758 49532
rect 5758 49476 5762 49532
rect 5698 49472 5762 49476
rect 5778 49532 5842 49536
rect 5778 49476 5782 49532
rect 5782 49476 5838 49532
rect 5838 49476 5842 49532
rect 5778 49472 5842 49476
rect 5858 49532 5922 49536
rect 5858 49476 5862 49532
rect 5862 49476 5918 49532
rect 5918 49476 5922 49532
rect 5858 49472 5922 49476
rect 10285 49532 10349 49536
rect 10285 49476 10289 49532
rect 10289 49476 10345 49532
rect 10345 49476 10349 49532
rect 10285 49472 10349 49476
rect 10365 49532 10429 49536
rect 10365 49476 10369 49532
rect 10369 49476 10425 49532
rect 10425 49476 10429 49532
rect 10365 49472 10429 49476
rect 10445 49532 10509 49536
rect 10445 49476 10449 49532
rect 10449 49476 10505 49532
rect 10505 49476 10509 49532
rect 10445 49472 10509 49476
rect 10525 49532 10589 49536
rect 10525 49476 10529 49532
rect 10529 49476 10585 49532
rect 10585 49476 10589 49532
rect 10525 49472 10589 49476
rect 3285 48988 3349 48992
rect 3285 48932 3289 48988
rect 3289 48932 3345 48988
rect 3345 48932 3349 48988
rect 3285 48928 3349 48932
rect 3365 48988 3429 48992
rect 3365 48932 3369 48988
rect 3369 48932 3425 48988
rect 3425 48932 3429 48988
rect 3365 48928 3429 48932
rect 3445 48988 3509 48992
rect 3445 48932 3449 48988
rect 3449 48932 3505 48988
rect 3505 48932 3509 48988
rect 3445 48928 3509 48932
rect 3525 48988 3589 48992
rect 3525 48932 3529 48988
rect 3529 48932 3585 48988
rect 3585 48932 3589 48988
rect 3525 48928 3589 48932
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 5618 48444 5682 48448
rect 5618 48388 5622 48444
rect 5622 48388 5678 48444
rect 5678 48388 5682 48444
rect 5618 48384 5682 48388
rect 5698 48444 5762 48448
rect 5698 48388 5702 48444
rect 5702 48388 5758 48444
rect 5758 48388 5762 48444
rect 5698 48384 5762 48388
rect 5778 48444 5842 48448
rect 5778 48388 5782 48444
rect 5782 48388 5838 48444
rect 5838 48388 5842 48444
rect 5778 48384 5842 48388
rect 5858 48444 5922 48448
rect 5858 48388 5862 48444
rect 5862 48388 5918 48444
rect 5918 48388 5922 48444
rect 5858 48384 5922 48388
rect 10285 48444 10349 48448
rect 10285 48388 10289 48444
rect 10289 48388 10345 48444
rect 10345 48388 10349 48444
rect 10285 48384 10349 48388
rect 10365 48444 10429 48448
rect 10365 48388 10369 48444
rect 10369 48388 10425 48444
rect 10425 48388 10429 48444
rect 10365 48384 10429 48388
rect 10445 48444 10509 48448
rect 10445 48388 10449 48444
rect 10449 48388 10505 48444
rect 10505 48388 10509 48444
rect 10445 48384 10509 48388
rect 10525 48444 10589 48448
rect 10525 48388 10529 48444
rect 10529 48388 10585 48444
rect 10585 48388 10589 48444
rect 10525 48384 10589 48388
rect 3285 47900 3349 47904
rect 3285 47844 3289 47900
rect 3289 47844 3345 47900
rect 3345 47844 3349 47900
rect 3285 47840 3349 47844
rect 3365 47900 3429 47904
rect 3365 47844 3369 47900
rect 3369 47844 3425 47900
rect 3425 47844 3429 47900
rect 3365 47840 3429 47844
rect 3445 47900 3509 47904
rect 3445 47844 3449 47900
rect 3449 47844 3505 47900
rect 3505 47844 3509 47900
rect 3445 47840 3509 47844
rect 3525 47900 3589 47904
rect 3525 47844 3529 47900
rect 3529 47844 3585 47900
rect 3585 47844 3589 47900
rect 3525 47840 3589 47844
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 5618 47356 5682 47360
rect 5618 47300 5622 47356
rect 5622 47300 5678 47356
rect 5678 47300 5682 47356
rect 5618 47296 5682 47300
rect 5698 47356 5762 47360
rect 5698 47300 5702 47356
rect 5702 47300 5758 47356
rect 5758 47300 5762 47356
rect 5698 47296 5762 47300
rect 5778 47356 5842 47360
rect 5778 47300 5782 47356
rect 5782 47300 5838 47356
rect 5838 47300 5842 47356
rect 5778 47296 5842 47300
rect 5858 47356 5922 47360
rect 5858 47300 5862 47356
rect 5862 47300 5918 47356
rect 5918 47300 5922 47356
rect 5858 47296 5922 47300
rect 10285 47356 10349 47360
rect 10285 47300 10289 47356
rect 10289 47300 10345 47356
rect 10345 47300 10349 47356
rect 10285 47296 10349 47300
rect 10365 47356 10429 47360
rect 10365 47300 10369 47356
rect 10369 47300 10425 47356
rect 10425 47300 10429 47356
rect 10365 47296 10429 47300
rect 10445 47356 10509 47360
rect 10445 47300 10449 47356
rect 10449 47300 10505 47356
rect 10505 47300 10509 47356
rect 10445 47296 10509 47300
rect 10525 47356 10589 47360
rect 10525 47300 10529 47356
rect 10529 47300 10585 47356
rect 10585 47300 10589 47356
rect 10525 47296 10589 47300
rect 3285 46812 3349 46816
rect 3285 46756 3289 46812
rect 3289 46756 3345 46812
rect 3345 46756 3349 46812
rect 3285 46752 3349 46756
rect 3365 46812 3429 46816
rect 3365 46756 3369 46812
rect 3369 46756 3425 46812
rect 3425 46756 3429 46812
rect 3365 46752 3429 46756
rect 3445 46812 3509 46816
rect 3445 46756 3449 46812
rect 3449 46756 3505 46812
rect 3505 46756 3509 46812
rect 3445 46752 3509 46756
rect 3525 46812 3589 46816
rect 3525 46756 3529 46812
rect 3529 46756 3585 46812
rect 3585 46756 3589 46812
rect 3525 46752 3589 46756
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 5618 46268 5682 46272
rect 5618 46212 5622 46268
rect 5622 46212 5678 46268
rect 5678 46212 5682 46268
rect 5618 46208 5682 46212
rect 5698 46268 5762 46272
rect 5698 46212 5702 46268
rect 5702 46212 5758 46268
rect 5758 46212 5762 46268
rect 5698 46208 5762 46212
rect 5778 46268 5842 46272
rect 5778 46212 5782 46268
rect 5782 46212 5838 46268
rect 5838 46212 5842 46268
rect 5778 46208 5842 46212
rect 5858 46268 5922 46272
rect 5858 46212 5862 46268
rect 5862 46212 5918 46268
rect 5918 46212 5922 46268
rect 5858 46208 5922 46212
rect 10285 46268 10349 46272
rect 10285 46212 10289 46268
rect 10289 46212 10345 46268
rect 10345 46212 10349 46268
rect 10285 46208 10349 46212
rect 10365 46268 10429 46272
rect 10365 46212 10369 46268
rect 10369 46212 10425 46268
rect 10425 46212 10429 46268
rect 10365 46208 10429 46212
rect 10445 46268 10509 46272
rect 10445 46212 10449 46268
rect 10449 46212 10505 46268
rect 10505 46212 10509 46268
rect 10445 46208 10509 46212
rect 10525 46268 10589 46272
rect 10525 46212 10529 46268
rect 10529 46212 10585 46268
rect 10585 46212 10589 46268
rect 10525 46208 10589 46212
rect 3285 45724 3349 45728
rect 3285 45668 3289 45724
rect 3289 45668 3345 45724
rect 3345 45668 3349 45724
rect 3285 45664 3349 45668
rect 3365 45724 3429 45728
rect 3365 45668 3369 45724
rect 3369 45668 3425 45724
rect 3425 45668 3429 45724
rect 3365 45664 3429 45668
rect 3445 45724 3509 45728
rect 3445 45668 3449 45724
rect 3449 45668 3505 45724
rect 3505 45668 3509 45724
rect 3445 45664 3509 45668
rect 3525 45724 3589 45728
rect 3525 45668 3529 45724
rect 3529 45668 3585 45724
rect 3585 45668 3589 45724
rect 3525 45664 3589 45668
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 5618 45180 5682 45184
rect 5618 45124 5622 45180
rect 5622 45124 5678 45180
rect 5678 45124 5682 45180
rect 5618 45120 5682 45124
rect 5698 45180 5762 45184
rect 5698 45124 5702 45180
rect 5702 45124 5758 45180
rect 5758 45124 5762 45180
rect 5698 45120 5762 45124
rect 5778 45180 5842 45184
rect 5778 45124 5782 45180
rect 5782 45124 5838 45180
rect 5838 45124 5842 45180
rect 5778 45120 5842 45124
rect 5858 45180 5922 45184
rect 5858 45124 5862 45180
rect 5862 45124 5918 45180
rect 5918 45124 5922 45180
rect 5858 45120 5922 45124
rect 10285 45180 10349 45184
rect 10285 45124 10289 45180
rect 10289 45124 10345 45180
rect 10345 45124 10349 45180
rect 10285 45120 10349 45124
rect 10365 45180 10429 45184
rect 10365 45124 10369 45180
rect 10369 45124 10425 45180
rect 10425 45124 10429 45180
rect 10365 45120 10429 45124
rect 10445 45180 10509 45184
rect 10445 45124 10449 45180
rect 10449 45124 10505 45180
rect 10505 45124 10509 45180
rect 10445 45120 10509 45124
rect 10525 45180 10589 45184
rect 10525 45124 10529 45180
rect 10529 45124 10585 45180
rect 10585 45124 10589 45180
rect 10525 45120 10589 45124
rect 3285 44636 3349 44640
rect 3285 44580 3289 44636
rect 3289 44580 3345 44636
rect 3345 44580 3349 44636
rect 3285 44576 3349 44580
rect 3365 44636 3429 44640
rect 3365 44580 3369 44636
rect 3369 44580 3425 44636
rect 3425 44580 3429 44636
rect 3365 44576 3429 44580
rect 3445 44636 3509 44640
rect 3445 44580 3449 44636
rect 3449 44580 3505 44636
rect 3505 44580 3509 44636
rect 3445 44576 3509 44580
rect 3525 44636 3589 44640
rect 3525 44580 3529 44636
rect 3529 44580 3585 44636
rect 3585 44580 3589 44636
rect 3525 44576 3589 44580
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 5618 44092 5682 44096
rect 5618 44036 5622 44092
rect 5622 44036 5678 44092
rect 5678 44036 5682 44092
rect 5618 44032 5682 44036
rect 5698 44092 5762 44096
rect 5698 44036 5702 44092
rect 5702 44036 5758 44092
rect 5758 44036 5762 44092
rect 5698 44032 5762 44036
rect 5778 44092 5842 44096
rect 5778 44036 5782 44092
rect 5782 44036 5838 44092
rect 5838 44036 5842 44092
rect 5778 44032 5842 44036
rect 5858 44092 5922 44096
rect 5858 44036 5862 44092
rect 5862 44036 5918 44092
rect 5918 44036 5922 44092
rect 5858 44032 5922 44036
rect 10285 44092 10349 44096
rect 10285 44036 10289 44092
rect 10289 44036 10345 44092
rect 10345 44036 10349 44092
rect 10285 44032 10349 44036
rect 10365 44092 10429 44096
rect 10365 44036 10369 44092
rect 10369 44036 10425 44092
rect 10425 44036 10429 44092
rect 10365 44032 10429 44036
rect 10445 44092 10509 44096
rect 10445 44036 10449 44092
rect 10449 44036 10505 44092
rect 10505 44036 10509 44092
rect 10445 44032 10509 44036
rect 10525 44092 10589 44096
rect 10525 44036 10529 44092
rect 10529 44036 10585 44092
rect 10585 44036 10589 44092
rect 10525 44032 10589 44036
rect 3285 43548 3349 43552
rect 3285 43492 3289 43548
rect 3289 43492 3345 43548
rect 3345 43492 3349 43548
rect 3285 43488 3349 43492
rect 3365 43548 3429 43552
rect 3365 43492 3369 43548
rect 3369 43492 3425 43548
rect 3425 43492 3429 43548
rect 3365 43488 3429 43492
rect 3445 43548 3509 43552
rect 3445 43492 3449 43548
rect 3449 43492 3505 43548
rect 3505 43492 3509 43548
rect 3445 43488 3509 43492
rect 3525 43548 3589 43552
rect 3525 43492 3529 43548
rect 3529 43492 3585 43548
rect 3585 43492 3589 43548
rect 3525 43488 3589 43492
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 5618 43004 5682 43008
rect 5618 42948 5622 43004
rect 5622 42948 5678 43004
rect 5678 42948 5682 43004
rect 5618 42944 5682 42948
rect 5698 43004 5762 43008
rect 5698 42948 5702 43004
rect 5702 42948 5758 43004
rect 5758 42948 5762 43004
rect 5698 42944 5762 42948
rect 5778 43004 5842 43008
rect 5778 42948 5782 43004
rect 5782 42948 5838 43004
rect 5838 42948 5842 43004
rect 5778 42944 5842 42948
rect 5858 43004 5922 43008
rect 5858 42948 5862 43004
rect 5862 42948 5918 43004
rect 5918 42948 5922 43004
rect 5858 42944 5922 42948
rect 10285 43004 10349 43008
rect 10285 42948 10289 43004
rect 10289 42948 10345 43004
rect 10345 42948 10349 43004
rect 10285 42944 10349 42948
rect 10365 43004 10429 43008
rect 10365 42948 10369 43004
rect 10369 42948 10425 43004
rect 10425 42948 10429 43004
rect 10365 42944 10429 42948
rect 10445 43004 10509 43008
rect 10445 42948 10449 43004
rect 10449 42948 10505 43004
rect 10505 42948 10509 43004
rect 10445 42944 10509 42948
rect 10525 43004 10589 43008
rect 10525 42948 10529 43004
rect 10529 42948 10585 43004
rect 10585 42948 10589 43004
rect 10525 42944 10589 42948
rect 3285 42460 3349 42464
rect 3285 42404 3289 42460
rect 3289 42404 3345 42460
rect 3345 42404 3349 42460
rect 3285 42400 3349 42404
rect 3365 42460 3429 42464
rect 3365 42404 3369 42460
rect 3369 42404 3425 42460
rect 3425 42404 3429 42460
rect 3365 42400 3429 42404
rect 3445 42460 3509 42464
rect 3445 42404 3449 42460
rect 3449 42404 3505 42460
rect 3505 42404 3509 42460
rect 3445 42400 3509 42404
rect 3525 42460 3589 42464
rect 3525 42404 3529 42460
rect 3529 42404 3585 42460
rect 3585 42404 3589 42460
rect 3525 42400 3589 42404
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 5618 41916 5682 41920
rect 5618 41860 5622 41916
rect 5622 41860 5678 41916
rect 5678 41860 5682 41916
rect 5618 41856 5682 41860
rect 5698 41916 5762 41920
rect 5698 41860 5702 41916
rect 5702 41860 5758 41916
rect 5758 41860 5762 41916
rect 5698 41856 5762 41860
rect 5778 41916 5842 41920
rect 5778 41860 5782 41916
rect 5782 41860 5838 41916
rect 5838 41860 5842 41916
rect 5778 41856 5842 41860
rect 5858 41916 5922 41920
rect 5858 41860 5862 41916
rect 5862 41860 5918 41916
rect 5918 41860 5922 41916
rect 5858 41856 5922 41860
rect 10285 41916 10349 41920
rect 10285 41860 10289 41916
rect 10289 41860 10345 41916
rect 10345 41860 10349 41916
rect 10285 41856 10349 41860
rect 10365 41916 10429 41920
rect 10365 41860 10369 41916
rect 10369 41860 10425 41916
rect 10425 41860 10429 41916
rect 10365 41856 10429 41860
rect 10445 41916 10509 41920
rect 10445 41860 10449 41916
rect 10449 41860 10505 41916
rect 10505 41860 10509 41916
rect 10445 41856 10509 41860
rect 10525 41916 10589 41920
rect 10525 41860 10529 41916
rect 10529 41860 10585 41916
rect 10585 41860 10589 41916
rect 10525 41856 10589 41860
rect 3285 41372 3349 41376
rect 3285 41316 3289 41372
rect 3289 41316 3345 41372
rect 3345 41316 3349 41372
rect 3285 41312 3349 41316
rect 3365 41372 3429 41376
rect 3365 41316 3369 41372
rect 3369 41316 3425 41372
rect 3425 41316 3429 41372
rect 3365 41312 3429 41316
rect 3445 41372 3509 41376
rect 3445 41316 3449 41372
rect 3449 41316 3505 41372
rect 3505 41316 3509 41372
rect 3445 41312 3509 41316
rect 3525 41372 3589 41376
rect 3525 41316 3529 41372
rect 3529 41316 3585 41372
rect 3585 41316 3589 41372
rect 3525 41312 3589 41316
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 5618 40828 5682 40832
rect 5618 40772 5622 40828
rect 5622 40772 5678 40828
rect 5678 40772 5682 40828
rect 5618 40768 5682 40772
rect 5698 40828 5762 40832
rect 5698 40772 5702 40828
rect 5702 40772 5758 40828
rect 5758 40772 5762 40828
rect 5698 40768 5762 40772
rect 5778 40828 5842 40832
rect 5778 40772 5782 40828
rect 5782 40772 5838 40828
rect 5838 40772 5842 40828
rect 5778 40768 5842 40772
rect 5858 40828 5922 40832
rect 5858 40772 5862 40828
rect 5862 40772 5918 40828
rect 5918 40772 5922 40828
rect 5858 40768 5922 40772
rect 10285 40828 10349 40832
rect 10285 40772 10289 40828
rect 10289 40772 10345 40828
rect 10345 40772 10349 40828
rect 10285 40768 10349 40772
rect 10365 40828 10429 40832
rect 10365 40772 10369 40828
rect 10369 40772 10425 40828
rect 10425 40772 10429 40828
rect 10365 40768 10429 40772
rect 10445 40828 10509 40832
rect 10445 40772 10449 40828
rect 10449 40772 10505 40828
rect 10505 40772 10509 40828
rect 10445 40768 10509 40772
rect 10525 40828 10589 40832
rect 10525 40772 10529 40828
rect 10529 40772 10585 40828
rect 10585 40772 10589 40828
rect 10525 40768 10589 40772
rect 3285 40284 3349 40288
rect 3285 40228 3289 40284
rect 3289 40228 3345 40284
rect 3345 40228 3349 40284
rect 3285 40224 3349 40228
rect 3365 40284 3429 40288
rect 3365 40228 3369 40284
rect 3369 40228 3425 40284
rect 3425 40228 3429 40284
rect 3365 40224 3429 40228
rect 3445 40284 3509 40288
rect 3445 40228 3449 40284
rect 3449 40228 3505 40284
rect 3505 40228 3509 40284
rect 3445 40224 3509 40228
rect 3525 40284 3589 40288
rect 3525 40228 3529 40284
rect 3529 40228 3585 40284
rect 3585 40228 3589 40284
rect 3525 40224 3589 40228
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 5618 39740 5682 39744
rect 5618 39684 5622 39740
rect 5622 39684 5678 39740
rect 5678 39684 5682 39740
rect 5618 39680 5682 39684
rect 5698 39740 5762 39744
rect 5698 39684 5702 39740
rect 5702 39684 5758 39740
rect 5758 39684 5762 39740
rect 5698 39680 5762 39684
rect 5778 39740 5842 39744
rect 5778 39684 5782 39740
rect 5782 39684 5838 39740
rect 5838 39684 5842 39740
rect 5778 39680 5842 39684
rect 5858 39740 5922 39744
rect 5858 39684 5862 39740
rect 5862 39684 5918 39740
rect 5918 39684 5922 39740
rect 5858 39680 5922 39684
rect 10285 39740 10349 39744
rect 10285 39684 10289 39740
rect 10289 39684 10345 39740
rect 10345 39684 10349 39740
rect 10285 39680 10349 39684
rect 10365 39740 10429 39744
rect 10365 39684 10369 39740
rect 10369 39684 10425 39740
rect 10425 39684 10429 39740
rect 10365 39680 10429 39684
rect 10445 39740 10509 39744
rect 10445 39684 10449 39740
rect 10449 39684 10505 39740
rect 10505 39684 10509 39740
rect 10445 39680 10509 39684
rect 10525 39740 10589 39744
rect 10525 39684 10529 39740
rect 10529 39684 10585 39740
rect 10585 39684 10589 39740
rect 10525 39680 10589 39684
rect 3285 39196 3349 39200
rect 3285 39140 3289 39196
rect 3289 39140 3345 39196
rect 3345 39140 3349 39196
rect 3285 39136 3349 39140
rect 3365 39196 3429 39200
rect 3365 39140 3369 39196
rect 3369 39140 3425 39196
rect 3425 39140 3429 39196
rect 3365 39136 3429 39140
rect 3445 39196 3509 39200
rect 3445 39140 3449 39196
rect 3449 39140 3505 39196
rect 3505 39140 3509 39196
rect 3445 39136 3509 39140
rect 3525 39196 3589 39200
rect 3525 39140 3529 39196
rect 3529 39140 3585 39196
rect 3585 39140 3589 39196
rect 3525 39136 3589 39140
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 5618 38652 5682 38656
rect 5618 38596 5622 38652
rect 5622 38596 5678 38652
rect 5678 38596 5682 38652
rect 5618 38592 5682 38596
rect 5698 38652 5762 38656
rect 5698 38596 5702 38652
rect 5702 38596 5758 38652
rect 5758 38596 5762 38652
rect 5698 38592 5762 38596
rect 5778 38652 5842 38656
rect 5778 38596 5782 38652
rect 5782 38596 5838 38652
rect 5838 38596 5842 38652
rect 5778 38592 5842 38596
rect 5858 38652 5922 38656
rect 5858 38596 5862 38652
rect 5862 38596 5918 38652
rect 5918 38596 5922 38652
rect 5858 38592 5922 38596
rect 10285 38652 10349 38656
rect 10285 38596 10289 38652
rect 10289 38596 10345 38652
rect 10345 38596 10349 38652
rect 10285 38592 10349 38596
rect 10365 38652 10429 38656
rect 10365 38596 10369 38652
rect 10369 38596 10425 38652
rect 10425 38596 10429 38652
rect 10365 38592 10429 38596
rect 10445 38652 10509 38656
rect 10445 38596 10449 38652
rect 10449 38596 10505 38652
rect 10505 38596 10509 38652
rect 10445 38592 10509 38596
rect 10525 38652 10589 38656
rect 10525 38596 10529 38652
rect 10529 38596 10585 38652
rect 10585 38596 10589 38652
rect 10525 38592 10589 38596
rect 3285 38108 3349 38112
rect 3285 38052 3289 38108
rect 3289 38052 3345 38108
rect 3345 38052 3349 38108
rect 3285 38048 3349 38052
rect 3365 38108 3429 38112
rect 3365 38052 3369 38108
rect 3369 38052 3425 38108
rect 3425 38052 3429 38108
rect 3365 38048 3429 38052
rect 3445 38108 3509 38112
rect 3445 38052 3449 38108
rect 3449 38052 3505 38108
rect 3505 38052 3509 38108
rect 3445 38048 3509 38052
rect 3525 38108 3589 38112
rect 3525 38052 3529 38108
rect 3529 38052 3585 38108
rect 3585 38052 3589 38108
rect 3525 38048 3589 38052
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 5618 37564 5682 37568
rect 5618 37508 5622 37564
rect 5622 37508 5678 37564
rect 5678 37508 5682 37564
rect 5618 37504 5682 37508
rect 5698 37564 5762 37568
rect 5698 37508 5702 37564
rect 5702 37508 5758 37564
rect 5758 37508 5762 37564
rect 5698 37504 5762 37508
rect 5778 37564 5842 37568
rect 5778 37508 5782 37564
rect 5782 37508 5838 37564
rect 5838 37508 5842 37564
rect 5778 37504 5842 37508
rect 5858 37564 5922 37568
rect 5858 37508 5862 37564
rect 5862 37508 5918 37564
rect 5918 37508 5922 37564
rect 5858 37504 5922 37508
rect 10285 37564 10349 37568
rect 10285 37508 10289 37564
rect 10289 37508 10345 37564
rect 10345 37508 10349 37564
rect 10285 37504 10349 37508
rect 10365 37564 10429 37568
rect 10365 37508 10369 37564
rect 10369 37508 10425 37564
rect 10425 37508 10429 37564
rect 10365 37504 10429 37508
rect 10445 37564 10509 37568
rect 10445 37508 10449 37564
rect 10449 37508 10505 37564
rect 10505 37508 10509 37564
rect 10445 37504 10509 37508
rect 10525 37564 10589 37568
rect 10525 37508 10529 37564
rect 10529 37508 10585 37564
rect 10585 37508 10589 37564
rect 10525 37504 10589 37508
rect 3285 37020 3349 37024
rect 3285 36964 3289 37020
rect 3289 36964 3345 37020
rect 3345 36964 3349 37020
rect 3285 36960 3349 36964
rect 3365 37020 3429 37024
rect 3365 36964 3369 37020
rect 3369 36964 3425 37020
rect 3425 36964 3429 37020
rect 3365 36960 3429 36964
rect 3445 37020 3509 37024
rect 3445 36964 3449 37020
rect 3449 36964 3505 37020
rect 3505 36964 3509 37020
rect 3445 36960 3509 36964
rect 3525 37020 3589 37024
rect 3525 36964 3529 37020
rect 3529 36964 3585 37020
rect 3585 36964 3589 37020
rect 3525 36960 3589 36964
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 5618 36476 5682 36480
rect 5618 36420 5622 36476
rect 5622 36420 5678 36476
rect 5678 36420 5682 36476
rect 5618 36416 5682 36420
rect 5698 36476 5762 36480
rect 5698 36420 5702 36476
rect 5702 36420 5758 36476
rect 5758 36420 5762 36476
rect 5698 36416 5762 36420
rect 5778 36476 5842 36480
rect 5778 36420 5782 36476
rect 5782 36420 5838 36476
rect 5838 36420 5842 36476
rect 5778 36416 5842 36420
rect 5858 36476 5922 36480
rect 5858 36420 5862 36476
rect 5862 36420 5918 36476
rect 5918 36420 5922 36476
rect 5858 36416 5922 36420
rect 10285 36476 10349 36480
rect 10285 36420 10289 36476
rect 10289 36420 10345 36476
rect 10345 36420 10349 36476
rect 10285 36416 10349 36420
rect 10365 36476 10429 36480
rect 10365 36420 10369 36476
rect 10369 36420 10425 36476
rect 10425 36420 10429 36476
rect 10365 36416 10429 36420
rect 10445 36476 10509 36480
rect 10445 36420 10449 36476
rect 10449 36420 10505 36476
rect 10505 36420 10509 36476
rect 10445 36416 10509 36420
rect 10525 36476 10589 36480
rect 10525 36420 10529 36476
rect 10529 36420 10585 36476
rect 10585 36420 10589 36476
rect 10525 36416 10589 36420
rect 3285 35932 3349 35936
rect 3285 35876 3289 35932
rect 3289 35876 3345 35932
rect 3345 35876 3349 35932
rect 3285 35872 3349 35876
rect 3365 35932 3429 35936
rect 3365 35876 3369 35932
rect 3369 35876 3425 35932
rect 3425 35876 3429 35932
rect 3365 35872 3429 35876
rect 3445 35932 3509 35936
rect 3445 35876 3449 35932
rect 3449 35876 3505 35932
rect 3505 35876 3509 35932
rect 3445 35872 3509 35876
rect 3525 35932 3589 35936
rect 3525 35876 3529 35932
rect 3529 35876 3585 35932
rect 3585 35876 3589 35932
rect 3525 35872 3589 35876
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 5618 35388 5682 35392
rect 5618 35332 5622 35388
rect 5622 35332 5678 35388
rect 5678 35332 5682 35388
rect 5618 35328 5682 35332
rect 5698 35388 5762 35392
rect 5698 35332 5702 35388
rect 5702 35332 5758 35388
rect 5758 35332 5762 35388
rect 5698 35328 5762 35332
rect 5778 35388 5842 35392
rect 5778 35332 5782 35388
rect 5782 35332 5838 35388
rect 5838 35332 5842 35388
rect 5778 35328 5842 35332
rect 5858 35388 5922 35392
rect 5858 35332 5862 35388
rect 5862 35332 5918 35388
rect 5918 35332 5922 35388
rect 5858 35328 5922 35332
rect 10285 35388 10349 35392
rect 10285 35332 10289 35388
rect 10289 35332 10345 35388
rect 10345 35332 10349 35388
rect 10285 35328 10349 35332
rect 10365 35388 10429 35392
rect 10365 35332 10369 35388
rect 10369 35332 10425 35388
rect 10425 35332 10429 35388
rect 10365 35328 10429 35332
rect 10445 35388 10509 35392
rect 10445 35332 10449 35388
rect 10449 35332 10505 35388
rect 10505 35332 10509 35388
rect 10445 35328 10509 35332
rect 10525 35388 10589 35392
rect 10525 35332 10529 35388
rect 10529 35332 10585 35388
rect 10585 35332 10589 35388
rect 10525 35328 10589 35332
rect 3285 34844 3349 34848
rect 3285 34788 3289 34844
rect 3289 34788 3345 34844
rect 3345 34788 3349 34844
rect 3285 34784 3349 34788
rect 3365 34844 3429 34848
rect 3365 34788 3369 34844
rect 3369 34788 3425 34844
rect 3425 34788 3429 34844
rect 3365 34784 3429 34788
rect 3445 34844 3509 34848
rect 3445 34788 3449 34844
rect 3449 34788 3505 34844
rect 3505 34788 3509 34844
rect 3445 34784 3509 34788
rect 3525 34844 3589 34848
rect 3525 34788 3529 34844
rect 3529 34788 3585 34844
rect 3585 34788 3589 34844
rect 3525 34784 3589 34788
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 5618 34300 5682 34304
rect 5618 34244 5622 34300
rect 5622 34244 5678 34300
rect 5678 34244 5682 34300
rect 5618 34240 5682 34244
rect 5698 34300 5762 34304
rect 5698 34244 5702 34300
rect 5702 34244 5758 34300
rect 5758 34244 5762 34300
rect 5698 34240 5762 34244
rect 5778 34300 5842 34304
rect 5778 34244 5782 34300
rect 5782 34244 5838 34300
rect 5838 34244 5842 34300
rect 5778 34240 5842 34244
rect 5858 34300 5922 34304
rect 5858 34244 5862 34300
rect 5862 34244 5918 34300
rect 5918 34244 5922 34300
rect 5858 34240 5922 34244
rect 10285 34300 10349 34304
rect 10285 34244 10289 34300
rect 10289 34244 10345 34300
rect 10345 34244 10349 34300
rect 10285 34240 10349 34244
rect 10365 34300 10429 34304
rect 10365 34244 10369 34300
rect 10369 34244 10425 34300
rect 10425 34244 10429 34300
rect 10365 34240 10429 34244
rect 10445 34300 10509 34304
rect 10445 34244 10449 34300
rect 10449 34244 10505 34300
rect 10505 34244 10509 34300
rect 10445 34240 10509 34244
rect 10525 34300 10589 34304
rect 10525 34244 10529 34300
rect 10529 34244 10585 34300
rect 10585 34244 10589 34300
rect 10525 34240 10589 34244
rect 3285 33756 3349 33760
rect 3285 33700 3289 33756
rect 3289 33700 3345 33756
rect 3345 33700 3349 33756
rect 3285 33696 3349 33700
rect 3365 33756 3429 33760
rect 3365 33700 3369 33756
rect 3369 33700 3425 33756
rect 3425 33700 3429 33756
rect 3365 33696 3429 33700
rect 3445 33756 3509 33760
rect 3445 33700 3449 33756
rect 3449 33700 3505 33756
rect 3505 33700 3509 33756
rect 3445 33696 3509 33700
rect 3525 33756 3589 33760
rect 3525 33700 3529 33756
rect 3529 33700 3585 33756
rect 3585 33700 3589 33756
rect 3525 33696 3589 33700
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 5618 33212 5682 33216
rect 5618 33156 5622 33212
rect 5622 33156 5678 33212
rect 5678 33156 5682 33212
rect 5618 33152 5682 33156
rect 5698 33212 5762 33216
rect 5698 33156 5702 33212
rect 5702 33156 5758 33212
rect 5758 33156 5762 33212
rect 5698 33152 5762 33156
rect 5778 33212 5842 33216
rect 5778 33156 5782 33212
rect 5782 33156 5838 33212
rect 5838 33156 5842 33212
rect 5778 33152 5842 33156
rect 5858 33212 5922 33216
rect 5858 33156 5862 33212
rect 5862 33156 5918 33212
rect 5918 33156 5922 33212
rect 5858 33152 5922 33156
rect 10285 33212 10349 33216
rect 10285 33156 10289 33212
rect 10289 33156 10345 33212
rect 10345 33156 10349 33212
rect 10285 33152 10349 33156
rect 10365 33212 10429 33216
rect 10365 33156 10369 33212
rect 10369 33156 10425 33212
rect 10425 33156 10429 33212
rect 10365 33152 10429 33156
rect 10445 33212 10509 33216
rect 10445 33156 10449 33212
rect 10449 33156 10505 33212
rect 10505 33156 10509 33212
rect 10445 33152 10509 33156
rect 10525 33212 10589 33216
rect 10525 33156 10529 33212
rect 10529 33156 10585 33212
rect 10585 33156 10589 33212
rect 10525 33152 10589 33156
rect 3285 32668 3349 32672
rect 3285 32612 3289 32668
rect 3289 32612 3345 32668
rect 3345 32612 3349 32668
rect 3285 32608 3349 32612
rect 3365 32668 3429 32672
rect 3365 32612 3369 32668
rect 3369 32612 3425 32668
rect 3425 32612 3429 32668
rect 3365 32608 3429 32612
rect 3445 32668 3509 32672
rect 3445 32612 3449 32668
rect 3449 32612 3505 32668
rect 3505 32612 3509 32668
rect 3445 32608 3509 32612
rect 3525 32668 3589 32672
rect 3525 32612 3529 32668
rect 3529 32612 3585 32668
rect 3585 32612 3589 32668
rect 3525 32608 3589 32612
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 5618 32124 5682 32128
rect 5618 32068 5622 32124
rect 5622 32068 5678 32124
rect 5678 32068 5682 32124
rect 5618 32064 5682 32068
rect 5698 32124 5762 32128
rect 5698 32068 5702 32124
rect 5702 32068 5758 32124
rect 5758 32068 5762 32124
rect 5698 32064 5762 32068
rect 5778 32124 5842 32128
rect 5778 32068 5782 32124
rect 5782 32068 5838 32124
rect 5838 32068 5842 32124
rect 5778 32064 5842 32068
rect 5858 32124 5922 32128
rect 5858 32068 5862 32124
rect 5862 32068 5918 32124
rect 5918 32068 5922 32124
rect 5858 32064 5922 32068
rect 10285 32124 10349 32128
rect 10285 32068 10289 32124
rect 10289 32068 10345 32124
rect 10345 32068 10349 32124
rect 10285 32064 10349 32068
rect 10365 32124 10429 32128
rect 10365 32068 10369 32124
rect 10369 32068 10425 32124
rect 10425 32068 10429 32124
rect 10365 32064 10429 32068
rect 10445 32124 10509 32128
rect 10445 32068 10449 32124
rect 10449 32068 10505 32124
rect 10505 32068 10509 32124
rect 10445 32064 10509 32068
rect 10525 32124 10589 32128
rect 10525 32068 10529 32124
rect 10529 32068 10585 32124
rect 10585 32068 10589 32124
rect 10525 32064 10589 32068
rect 3285 31580 3349 31584
rect 3285 31524 3289 31580
rect 3289 31524 3345 31580
rect 3345 31524 3349 31580
rect 3285 31520 3349 31524
rect 3365 31580 3429 31584
rect 3365 31524 3369 31580
rect 3369 31524 3425 31580
rect 3425 31524 3429 31580
rect 3365 31520 3429 31524
rect 3445 31580 3509 31584
rect 3445 31524 3449 31580
rect 3449 31524 3505 31580
rect 3505 31524 3509 31580
rect 3445 31520 3509 31524
rect 3525 31580 3589 31584
rect 3525 31524 3529 31580
rect 3529 31524 3585 31580
rect 3585 31524 3589 31580
rect 3525 31520 3589 31524
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 5618 31036 5682 31040
rect 5618 30980 5622 31036
rect 5622 30980 5678 31036
rect 5678 30980 5682 31036
rect 5618 30976 5682 30980
rect 5698 31036 5762 31040
rect 5698 30980 5702 31036
rect 5702 30980 5758 31036
rect 5758 30980 5762 31036
rect 5698 30976 5762 30980
rect 5778 31036 5842 31040
rect 5778 30980 5782 31036
rect 5782 30980 5838 31036
rect 5838 30980 5842 31036
rect 5778 30976 5842 30980
rect 5858 31036 5922 31040
rect 5858 30980 5862 31036
rect 5862 30980 5918 31036
rect 5918 30980 5922 31036
rect 5858 30976 5922 30980
rect 10285 31036 10349 31040
rect 10285 30980 10289 31036
rect 10289 30980 10345 31036
rect 10345 30980 10349 31036
rect 10285 30976 10349 30980
rect 10365 31036 10429 31040
rect 10365 30980 10369 31036
rect 10369 30980 10425 31036
rect 10425 30980 10429 31036
rect 10365 30976 10429 30980
rect 10445 31036 10509 31040
rect 10445 30980 10449 31036
rect 10449 30980 10505 31036
rect 10505 30980 10509 31036
rect 10445 30976 10509 30980
rect 10525 31036 10589 31040
rect 10525 30980 10529 31036
rect 10529 30980 10585 31036
rect 10585 30980 10589 31036
rect 10525 30976 10589 30980
rect 3285 30492 3349 30496
rect 3285 30436 3289 30492
rect 3289 30436 3345 30492
rect 3345 30436 3349 30492
rect 3285 30432 3349 30436
rect 3365 30492 3429 30496
rect 3365 30436 3369 30492
rect 3369 30436 3425 30492
rect 3425 30436 3429 30492
rect 3365 30432 3429 30436
rect 3445 30492 3509 30496
rect 3445 30436 3449 30492
rect 3449 30436 3505 30492
rect 3505 30436 3509 30492
rect 3445 30432 3509 30436
rect 3525 30492 3589 30496
rect 3525 30436 3529 30492
rect 3529 30436 3585 30492
rect 3585 30436 3589 30492
rect 3525 30432 3589 30436
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 5618 29948 5682 29952
rect 5618 29892 5622 29948
rect 5622 29892 5678 29948
rect 5678 29892 5682 29948
rect 5618 29888 5682 29892
rect 5698 29948 5762 29952
rect 5698 29892 5702 29948
rect 5702 29892 5758 29948
rect 5758 29892 5762 29948
rect 5698 29888 5762 29892
rect 5778 29948 5842 29952
rect 5778 29892 5782 29948
rect 5782 29892 5838 29948
rect 5838 29892 5842 29948
rect 5778 29888 5842 29892
rect 5858 29948 5922 29952
rect 5858 29892 5862 29948
rect 5862 29892 5918 29948
rect 5918 29892 5922 29948
rect 5858 29888 5922 29892
rect 10285 29948 10349 29952
rect 10285 29892 10289 29948
rect 10289 29892 10345 29948
rect 10345 29892 10349 29948
rect 10285 29888 10349 29892
rect 10365 29948 10429 29952
rect 10365 29892 10369 29948
rect 10369 29892 10425 29948
rect 10425 29892 10429 29948
rect 10365 29888 10429 29892
rect 10445 29948 10509 29952
rect 10445 29892 10449 29948
rect 10449 29892 10505 29948
rect 10505 29892 10509 29948
rect 10445 29888 10509 29892
rect 10525 29948 10589 29952
rect 10525 29892 10529 29948
rect 10529 29892 10585 29948
rect 10585 29892 10589 29948
rect 10525 29888 10589 29892
rect 3285 29404 3349 29408
rect 3285 29348 3289 29404
rect 3289 29348 3345 29404
rect 3345 29348 3349 29404
rect 3285 29344 3349 29348
rect 3365 29404 3429 29408
rect 3365 29348 3369 29404
rect 3369 29348 3425 29404
rect 3425 29348 3429 29404
rect 3365 29344 3429 29348
rect 3445 29404 3509 29408
rect 3445 29348 3449 29404
rect 3449 29348 3505 29404
rect 3505 29348 3509 29404
rect 3445 29344 3509 29348
rect 3525 29404 3589 29408
rect 3525 29348 3529 29404
rect 3529 29348 3585 29404
rect 3585 29348 3589 29404
rect 3525 29344 3589 29348
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 5618 28860 5682 28864
rect 5618 28804 5622 28860
rect 5622 28804 5678 28860
rect 5678 28804 5682 28860
rect 5618 28800 5682 28804
rect 5698 28860 5762 28864
rect 5698 28804 5702 28860
rect 5702 28804 5758 28860
rect 5758 28804 5762 28860
rect 5698 28800 5762 28804
rect 5778 28860 5842 28864
rect 5778 28804 5782 28860
rect 5782 28804 5838 28860
rect 5838 28804 5842 28860
rect 5778 28800 5842 28804
rect 5858 28860 5922 28864
rect 5858 28804 5862 28860
rect 5862 28804 5918 28860
rect 5918 28804 5922 28860
rect 5858 28800 5922 28804
rect 10285 28860 10349 28864
rect 10285 28804 10289 28860
rect 10289 28804 10345 28860
rect 10345 28804 10349 28860
rect 10285 28800 10349 28804
rect 10365 28860 10429 28864
rect 10365 28804 10369 28860
rect 10369 28804 10425 28860
rect 10425 28804 10429 28860
rect 10365 28800 10429 28804
rect 10445 28860 10509 28864
rect 10445 28804 10449 28860
rect 10449 28804 10505 28860
rect 10505 28804 10509 28860
rect 10445 28800 10509 28804
rect 10525 28860 10589 28864
rect 10525 28804 10529 28860
rect 10529 28804 10585 28860
rect 10585 28804 10589 28860
rect 10525 28800 10589 28804
rect 3285 28316 3349 28320
rect 3285 28260 3289 28316
rect 3289 28260 3345 28316
rect 3345 28260 3349 28316
rect 3285 28256 3349 28260
rect 3365 28316 3429 28320
rect 3365 28260 3369 28316
rect 3369 28260 3425 28316
rect 3425 28260 3429 28316
rect 3365 28256 3429 28260
rect 3445 28316 3509 28320
rect 3445 28260 3449 28316
rect 3449 28260 3505 28316
rect 3505 28260 3509 28316
rect 3445 28256 3509 28260
rect 3525 28316 3589 28320
rect 3525 28260 3529 28316
rect 3529 28260 3585 28316
rect 3585 28260 3589 28316
rect 3525 28256 3589 28260
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 5618 27772 5682 27776
rect 5618 27716 5622 27772
rect 5622 27716 5678 27772
rect 5678 27716 5682 27772
rect 5618 27712 5682 27716
rect 5698 27772 5762 27776
rect 5698 27716 5702 27772
rect 5702 27716 5758 27772
rect 5758 27716 5762 27772
rect 5698 27712 5762 27716
rect 5778 27772 5842 27776
rect 5778 27716 5782 27772
rect 5782 27716 5838 27772
rect 5838 27716 5842 27772
rect 5778 27712 5842 27716
rect 5858 27772 5922 27776
rect 5858 27716 5862 27772
rect 5862 27716 5918 27772
rect 5918 27716 5922 27772
rect 5858 27712 5922 27716
rect 10285 27772 10349 27776
rect 10285 27716 10289 27772
rect 10289 27716 10345 27772
rect 10345 27716 10349 27772
rect 10285 27712 10349 27716
rect 10365 27772 10429 27776
rect 10365 27716 10369 27772
rect 10369 27716 10425 27772
rect 10425 27716 10429 27772
rect 10365 27712 10429 27716
rect 10445 27772 10509 27776
rect 10445 27716 10449 27772
rect 10449 27716 10505 27772
rect 10505 27716 10509 27772
rect 10445 27712 10509 27716
rect 10525 27772 10589 27776
rect 10525 27716 10529 27772
rect 10529 27716 10585 27772
rect 10585 27716 10589 27772
rect 10525 27712 10589 27716
rect 3285 27228 3349 27232
rect 3285 27172 3289 27228
rect 3289 27172 3345 27228
rect 3345 27172 3349 27228
rect 3285 27168 3349 27172
rect 3365 27228 3429 27232
rect 3365 27172 3369 27228
rect 3369 27172 3425 27228
rect 3425 27172 3429 27228
rect 3365 27168 3429 27172
rect 3445 27228 3509 27232
rect 3445 27172 3449 27228
rect 3449 27172 3505 27228
rect 3505 27172 3509 27228
rect 3445 27168 3509 27172
rect 3525 27228 3589 27232
rect 3525 27172 3529 27228
rect 3529 27172 3585 27228
rect 3585 27172 3589 27228
rect 3525 27168 3589 27172
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 5618 26684 5682 26688
rect 5618 26628 5622 26684
rect 5622 26628 5678 26684
rect 5678 26628 5682 26684
rect 5618 26624 5682 26628
rect 5698 26684 5762 26688
rect 5698 26628 5702 26684
rect 5702 26628 5758 26684
rect 5758 26628 5762 26684
rect 5698 26624 5762 26628
rect 5778 26684 5842 26688
rect 5778 26628 5782 26684
rect 5782 26628 5838 26684
rect 5838 26628 5842 26684
rect 5778 26624 5842 26628
rect 5858 26684 5922 26688
rect 5858 26628 5862 26684
rect 5862 26628 5918 26684
rect 5918 26628 5922 26684
rect 5858 26624 5922 26628
rect 10285 26684 10349 26688
rect 10285 26628 10289 26684
rect 10289 26628 10345 26684
rect 10345 26628 10349 26684
rect 10285 26624 10349 26628
rect 10365 26684 10429 26688
rect 10365 26628 10369 26684
rect 10369 26628 10425 26684
rect 10425 26628 10429 26684
rect 10365 26624 10429 26628
rect 10445 26684 10509 26688
rect 10445 26628 10449 26684
rect 10449 26628 10505 26684
rect 10505 26628 10509 26684
rect 10445 26624 10509 26628
rect 10525 26684 10589 26688
rect 10525 26628 10529 26684
rect 10529 26628 10585 26684
rect 10585 26628 10589 26684
rect 10525 26624 10589 26628
rect 3285 26140 3349 26144
rect 3285 26084 3289 26140
rect 3289 26084 3345 26140
rect 3345 26084 3349 26140
rect 3285 26080 3349 26084
rect 3365 26140 3429 26144
rect 3365 26084 3369 26140
rect 3369 26084 3425 26140
rect 3425 26084 3429 26140
rect 3365 26080 3429 26084
rect 3445 26140 3509 26144
rect 3445 26084 3449 26140
rect 3449 26084 3505 26140
rect 3505 26084 3509 26140
rect 3445 26080 3509 26084
rect 3525 26140 3589 26144
rect 3525 26084 3529 26140
rect 3529 26084 3585 26140
rect 3585 26084 3589 26140
rect 3525 26080 3589 26084
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 5618 25596 5682 25600
rect 5618 25540 5622 25596
rect 5622 25540 5678 25596
rect 5678 25540 5682 25596
rect 5618 25536 5682 25540
rect 5698 25596 5762 25600
rect 5698 25540 5702 25596
rect 5702 25540 5758 25596
rect 5758 25540 5762 25596
rect 5698 25536 5762 25540
rect 5778 25596 5842 25600
rect 5778 25540 5782 25596
rect 5782 25540 5838 25596
rect 5838 25540 5842 25596
rect 5778 25536 5842 25540
rect 5858 25596 5922 25600
rect 5858 25540 5862 25596
rect 5862 25540 5918 25596
rect 5918 25540 5922 25596
rect 5858 25536 5922 25540
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 3285 25052 3349 25056
rect 3285 24996 3289 25052
rect 3289 24996 3345 25052
rect 3345 24996 3349 25052
rect 3285 24992 3349 24996
rect 3365 25052 3429 25056
rect 3365 24996 3369 25052
rect 3369 24996 3425 25052
rect 3425 24996 3429 25052
rect 3365 24992 3429 24996
rect 3445 25052 3509 25056
rect 3445 24996 3449 25052
rect 3449 24996 3505 25052
rect 3505 24996 3509 25052
rect 3445 24992 3509 24996
rect 3525 25052 3589 25056
rect 3525 24996 3529 25052
rect 3529 24996 3585 25052
rect 3585 24996 3589 25052
rect 3525 24992 3589 24996
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 5618 24508 5682 24512
rect 5618 24452 5622 24508
rect 5622 24452 5678 24508
rect 5678 24452 5682 24508
rect 5618 24448 5682 24452
rect 5698 24508 5762 24512
rect 5698 24452 5702 24508
rect 5702 24452 5758 24508
rect 5758 24452 5762 24508
rect 5698 24448 5762 24452
rect 5778 24508 5842 24512
rect 5778 24452 5782 24508
rect 5782 24452 5838 24508
rect 5838 24452 5842 24508
rect 5778 24448 5842 24452
rect 5858 24508 5922 24512
rect 5858 24452 5862 24508
rect 5862 24452 5918 24508
rect 5918 24452 5922 24508
rect 5858 24448 5922 24452
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 3285 23964 3349 23968
rect 3285 23908 3289 23964
rect 3289 23908 3345 23964
rect 3345 23908 3349 23964
rect 3285 23904 3349 23908
rect 3365 23964 3429 23968
rect 3365 23908 3369 23964
rect 3369 23908 3425 23964
rect 3425 23908 3429 23964
rect 3365 23904 3429 23908
rect 3445 23964 3509 23968
rect 3445 23908 3449 23964
rect 3449 23908 3505 23964
rect 3505 23908 3509 23964
rect 3445 23904 3509 23908
rect 3525 23964 3589 23968
rect 3525 23908 3529 23964
rect 3529 23908 3585 23964
rect 3585 23908 3589 23964
rect 3525 23904 3589 23908
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 5618 23420 5682 23424
rect 5618 23364 5622 23420
rect 5622 23364 5678 23420
rect 5678 23364 5682 23420
rect 5618 23360 5682 23364
rect 5698 23420 5762 23424
rect 5698 23364 5702 23420
rect 5702 23364 5758 23420
rect 5758 23364 5762 23420
rect 5698 23360 5762 23364
rect 5778 23420 5842 23424
rect 5778 23364 5782 23420
rect 5782 23364 5838 23420
rect 5838 23364 5842 23420
rect 5778 23360 5842 23364
rect 5858 23420 5922 23424
rect 5858 23364 5862 23420
rect 5862 23364 5918 23420
rect 5918 23364 5922 23420
rect 5858 23360 5922 23364
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 3285 22876 3349 22880
rect 3285 22820 3289 22876
rect 3289 22820 3345 22876
rect 3345 22820 3349 22876
rect 3285 22816 3349 22820
rect 3365 22876 3429 22880
rect 3365 22820 3369 22876
rect 3369 22820 3425 22876
rect 3425 22820 3429 22876
rect 3365 22816 3429 22820
rect 3445 22876 3509 22880
rect 3445 22820 3449 22876
rect 3449 22820 3505 22876
rect 3505 22820 3509 22876
rect 3445 22816 3509 22820
rect 3525 22876 3589 22880
rect 3525 22820 3529 22876
rect 3529 22820 3585 22876
rect 3585 22820 3589 22876
rect 3525 22816 3589 22820
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 5618 22332 5682 22336
rect 5618 22276 5622 22332
rect 5622 22276 5678 22332
rect 5678 22276 5682 22332
rect 5618 22272 5682 22276
rect 5698 22332 5762 22336
rect 5698 22276 5702 22332
rect 5702 22276 5758 22332
rect 5758 22276 5762 22332
rect 5698 22272 5762 22276
rect 5778 22332 5842 22336
rect 5778 22276 5782 22332
rect 5782 22276 5838 22332
rect 5838 22276 5842 22332
rect 5778 22272 5842 22276
rect 5858 22332 5922 22336
rect 5858 22276 5862 22332
rect 5862 22276 5918 22332
rect 5918 22276 5922 22332
rect 5858 22272 5922 22276
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 3285 21788 3349 21792
rect 3285 21732 3289 21788
rect 3289 21732 3345 21788
rect 3345 21732 3349 21788
rect 3285 21728 3349 21732
rect 3365 21788 3429 21792
rect 3365 21732 3369 21788
rect 3369 21732 3425 21788
rect 3425 21732 3429 21788
rect 3365 21728 3429 21732
rect 3445 21788 3509 21792
rect 3445 21732 3449 21788
rect 3449 21732 3505 21788
rect 3505 21732 3509 21788
rect 3445 21728 3509 21732
rect 3525 21788 3589 21792
rect 3525 21732 3529 21788
rect 3529 21732 3585 21788
rect 3585 21732 3589 21788
rect 3525 21728 3589 21732
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 5618 21244 5682 21248
rect 5618 21188 5622 21244
rect 5622 21188 5678 21244
rect 5678 21188 5682 21244
rect 5618 21184 5682 21188
rect 5698 21244 5762 21248
rect 5698 21188 5702 21244
rect 5702 21188 5758 21244
rect 5758 21188 5762 21244
rect 5698 21184 5762 21188
rect 5778 21244 5842 21248
rect 5778 21188 5782 21244
rect 5782 21188 5838 21244
rect 5838 21188 5842 21244
rect 5778 21184 5842 21188
rect 5858 21244 5922 21248
rect 5858 21188 5862 21244
rect 5862 21188 5918 21244
rect 5918 21188 5922 21244
rect 5858 21184 5922 21188
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 3285 20700 3349 20704
rect 3285 20644 3289 20700
rect 3289 20644 3345 20700
rect 3345 20644 3349 20700
rect 3285 20640 3349 20644
rect 3365 20700 3429 20704
rect 3365 20644 3369 20700
rect 3369 20644 3425 20700
rect 3425 20644 3429 20700
rect 3365 20640 3429 20644
rect 3445 20700 3509 20704
rect 3445 20644 3449 20700
rect 3449 20644 3505 20700
rect 3505 20644 3509 20700
rect 3445 20640 3509 20644
rect 3525 20700 3589 20704
rect 3525 20644 3529 20700
rect 3529 20644 3585 20700
rect 3585 20644 3589 20700
rect 3525 20640 3589 20644
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 5618 20156 5682 20160
rect 5618 20100 5622 20156
rect 5622 20100 5678 20156
rect 5678 20100 5682 20156
rect 5618 20096 5682 20100
rect 5698 20156 5762 20160
rect 5698 20100 5702 20156
rect 5702 20100 5758 20156
rect 5758 20100 5762 20156
rect 5698 20096 5762 20100
rect 5778 20156 5842 20160
rect 5778 20100 5782 20156
rect 5782 20100 5838 20156
rect 5838 20100 5842 20156
rect 5778 20096 5842 20100
rect 5858 20156 5922 20160
rect 5858 20100 5862 20156
rect 5862 20100 5918 20156
rect 5918 20100 5922 20156
rect 5858 20096 5922 20100
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 3285 19612 3349 19616
rect 3285 19556 3289 19612
rect 3289 19556 3345 19612
rect 3345 19556 3349 19612
rect 3285 19552 3349 19556
rect 3365 19612 3429 19616
rect 3365 19556 3369 19612
rect 3369 19556 3425 19612
rect 3425 19556 3429 19612
rect 3365 19552 3429 19556
rect 3445 19612 3509 19616
rect 3445 19556 3449 19612
rect 3449 19556 3505 19612
rect 3505 19556 3509 19612
rect 3445 19552 3509 19556
rect 3525 19612 3589 19616
rect 3525 19556 3529 19612
rect 3529 19556 3585 19612
rect 3585 19556 3589 19612
rect 3525 19552 3589 19556
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 5618 19068 5682 19072
rect 5618 19012 5622 19068
rect 5622 19012 5678 19068
rect 5678 19012 5682 19068
rect 5618 19008 5682 19012
rect 5698 19068 5762 19072
rect 5698 19012 5702 19068
rect 5702 19012 5758 19068
rect 5758 19012 5762 19068
rect 5698 19008 5762 19012
rect 5778 19068 5842 19072
rect 5778 19012 5782 19068
rect 5782 19012 5838 19068
rect 5838 19012 5842 19068
rect 5778 19008 5842 19012
rect 5858 19068 5922 19072
rect 5858 19012 5862 19068
rect 5862 19012 5918 19068
rect 5918 19012 5922 19068
rect 5858 19008 5922 19012
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 3285 18524 3349 18528
rect 3285 18468 3289 18524
rect 3289 18468 3345 18524
rect 3345 18468 3349 18524
rect 3285 18464 3349 18468
rect 3365 18524 3429 18528
rect 3365 18468 3369 18524
rect 3369 18468 3425 18524
rect 3425 18468 3429 18524
rect 3365 18464 3429 18468
rect 3445 18524 3509 18528
rect 3445 18468 3449 18524
rect 3449 18468 3505 18524
rect 3505 18468 3509 18524
rect 3445 18464 3509 18468
rect 3525 18524 3589 18528
rect 3525 18468 3529 18524
rect 3529 18468 3585 18524
rect 3585 18468 3589 18524
rect 3525 18464 3589 18468
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 5618 17980 5682 17984
rect 5618 17924 5622 17980
rect 5622 17924 5678 17980
rect 5678 17924 5682 17980
rect 5618 17920 5682 17924
rect 5698 17980 5762 17984
rect 5698 17924 5702 17980
rect 5702 17924 5758 17980
rect 5758 17924 5762 17980
rect 5698 17920 5762 17924
rect 5778 17980 5842 17984
rect 5778 17924 5782 17980
rect 5782 17924 5838 17980
rect 5838 17924 5842 17980
rect 5778 17920 5842 17924
rect 5858 17980 5922 17984
rect 5858 17924 5862 17980
rect 5862 17924 5918 17980
rect 5918 17924 5922 17980
rect 5858 17920 5922 17924
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 3285 17436 3349 17440
rect 3285 17380 3289 17436
rect 3289 17380 3345 17436
rect 3345 17380 3349 17436
rect 3285 17376 3349 17380
rect 3365 17436 3429 17440
rect 3365 17380 3369 17436
rect 3369 17380 3425 17436
rect 3425 17380 3429 17436
rect 3365 17376 3429 17380
rect 3445 17436 3509 17440
rect 3445 17380 3449 17436
rect 3449 17380 3505 17436
rect 3505 17380 3509 17436
rect 3445 17376 3509 17380
rect 3525 17436 3589 17440
rect 3525 17380 3529 17436
rect 3529 17380 3585 17436
rect 3585 17380 3589 17436
rect 3525 17376 3589 17380
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 5618 16892 5682 16896
rect 5618 16836 5622 16892
rect 5622 16836 5678 16892
rect 5678 16836 5682 16892
rect 5618 16832 5682 16836
rect 5698 16892 5762 16896
rect 5698 16836 5702 16892
rect 5702 16836 5758 16892
rect 5758 16836 5762 16892
rect 5698 16832 5762 16836
rect 5778 16892 5842 16896
rect 5778 16836 5782 16892
rect 5782 16836 5838 16892
rect 5838 16836 5842 16892
rect 5778 16832 5842 16836
rect 5858 16892 5922 16896
rect 5858 16836 5862 16892
rect 5862 16836 5918 16892
rect 5918 16836 5922 16892
rect 5858 16832 5922 16836
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 3285 16348 3349 16352
rect 3285 16292 3289 16348
rect 3289 16292 3345 16348
rect 3345 16292 3349 16348
rect 3285 16288 3349 16292
rect 3365 16348 3429 16352
rect 3365 16292 3369 16348
rect 3369 16292 3425 16348
rect 3425 16292 3429 16348
rect 3365 16288 3429 16292
rect 3445 16348 3509 16352
rect 3445 16292 3449 16348
rect 3449 16292 3505 16348
rect 3505 16292 3509 16348
rect 3445 16288 3509 16292
rect 3525 16348 3589 16352
rect 3525 16292 3529 16348
rect 3529 16292 3585 16348
rect 3585 16292 3589 16348
rect 3525 16288 3589 16292
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 5618 15804 5682 15808
rect 5618 15748 5622 15804
rect 5622 15748 5678 15804
rect 5678 15748 5682 15804
rect 5618 15744 5682 15748
rect 5698 15804 5762 15808
rect 5698 15748 5702 15804
rect 5702 15748 5758 15804
rect 5758 15748 5762 15804
rect 5698 15744 5762 15748
rect 5778 15804 5842 15808
rect 5778 15748 5782 15804
rect 5782 15748 5838 15804
rect 5838 15748 5842 15804
rect 5778 15744 5842 15748
rect 5858 15804 5922 15808
rect 5858 15748 5862 15804
rect 5862 15748 5918 15804
rect 5918 15748 5922 15804
rect 5858 15744 5922 15748
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 3285 15260 3349 15264
rect 3285 15204 3289 15260
rect 3289 15204 3345 15260
rect 3345 15204 3349 15260
rect 3285 15200 3349 15204
rect 3365 15260 3429 15264
rect 3365 15204 3369 15260
rect 3369 15204 3425 15260
rect 3425 15204 3429 15260
rect 3365 15200 3429 15204
rect 3445 15260 3509 15264
rect 3445 15204 3449 15260
rect 3449 15204 3505 15260
rect 3505 15204 3509 15260
rect 3445 15200 3509 15204
rect 3525 15260 3589 15264
rect 3525 15204 3529 15260
rect 3529 15204 3585 15260
rect 3585 15204 3589 15260
rect 3525 15200 3589 15204
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 5618 14716 5682 14720
rect 5618 14660 5622 14716
rect 5622 14660 5678 14716
rect 5678 14660 5682 14716
rect 5618 14656 5682 14660
rect 5698 14716 5762 14720
rect 5698 14660 5702 14716
rect 5702 14660 5758 14716
rect 5758 14660 5762 14716
rect 5698 14656 5762 14660
rect 5778 14716 5842 14720
rect 5778 14660 5782 14716
rect 5782 14660 5838 14716
rect 5838 14660 5842 14716
rect 5778 14656 5842 14660
rect 5858 14716 5922 14720
rect 5858 14660 5862 14716
rect 5862 14660 5918 14716
rect 5918 14660 5922 14716
rect 5858 14656 5922 14660
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 3285 14172 3349 14176
rect 3285 14116 3289 14172
rect 3289 14116 3345 14172
rect 3345 14116 3349 14172
rect 3285 14112 3349 14116
rect 3365 14172 3429 14176
rect 3365 14116 3369 14172
rect 3369 14116 3425 14172
rect 3425 14116 3429 14172
rect 3365 14112 3429 14116
rect 3445 14172 3509 14176
rect 3445 14116 3449 14172
rect 3449 14116 3505 14172
rect 3505 14116 3509 14172
rect 3445 14112 3509 14116
rect 3525 14172 3589 14176
rect 3525 14116 3529 14172
rect 3529 14116 3585 14172
rect 3585 14116 3589 14172
rect 3525 14112 3589 14116
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 5618 13628 5682 13632
rect 5618 13572 5622 13628
rect 5622 13572 5678 13628
rect 5678 13572 5682 13628
rect 5618 13568 5682 13572
rect 5698 13628 5762 13632
rect 5698 13572 5702 13628
rect 5702 13572 5758 13628
rect 5758 13572 5762 13628
rect 5698 13568 5762 13572
rect 5778 13628 5842 13632
rect 5778 13572 5782 13628
rect 5782 13572 5838 13628
rect 5838 13572 5842 13628
rect 5778 13568 5842 13572
rect 5858 13628 5922 13632
rect 5858 13572 5862 13628
rect 5862 13572 5918 13628
rect 5918 13572 5922 13628
rect 5858 13568 5922 13572
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 3285 13084 3349 13088
rect 3285 13028 3289 13084
rect 3289 13028 3345 13084
rect 3345 13028 3349 13084
rect 3285 13024 3349 13028
rect 3365 13084 3429 13088
rect 3365 13028 3369 13084
rect 3369 13028 3425 13084
rect 3425 13028 3429 13084
rect 3365 13024 3429 13028
rect 3445 13084 3509 13088
rect 3445 13028 3449 13084
rect 3449 13028 3505 13084
rect 3505 13028 3509 13084
rect 3445 13024 3509 13028
rect 3525 13084 3589 13088
rect 3525 13028 3529 13084
rect 3529 13028 3585 13084
rect 3585 13028 3589 13084
rect 3525 13024 3589 13028
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 5618 12540 5682 12544
rect 5618 12484 5622 12540
rect 5622 12484 5678 12540
rect 5678 12484 5682 12540
rect 5618 12480 5682 12484
rect 5698 12540 5762 12544
rect 5698 12484 5702 12540
rect 5702 12484 5758 12540
rect 5758 12484 5762 12540
rect 5698 12480 5762 12484
rect 5778 12540 5842 12544
rect 5778 12484 5782 12540
rect 5782 12484 5838 12540
rect 5838 12484 5842 12540
rect 5778 12480 5842 12484
rect 5858 12540 5922 12544
rect 5858 12484 5862 12540
rect 5862 12484 5918 12540
rect 5918 12484 5922 12540
rect 5858 12480 5922 12484
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 3285 11996 3349 12000
rect 3285 11940 3289 11996
rect 3289 11940 3345 11996
rect 3345 11940 3349 11996
rect 3285 11936 3349 11940
rect 3365 11996 3429 12000
rect 3365 11940 3369 11996
rect 3369 11940 3425 11996
rect 3425 11940 3429 11996
rect 3365 11936 3429 11940
rect 3445 11996 3509 12000
rect 3445 11940 3449 11996
rect 3449 11940 3505 11996
rect 3505 11940 3509 11996
rect 3445 11936 3509 11940
rect 3525 11996 3589 12000
rect 3525 11940 3529 11996
rect 3529 11940 3585 11996
rect 3585 11940 3589 11996
rect 3525 11936 3589 11940
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 5618 11452 5682 11456
rect 5618 11396 5622 11452
rect 5622 11396 5678 11452
rect 5678 11396 5682 11452
rect 5618 11392 5682 11396
rect 5698 11452 5762 11456
rect 5698 11396 5702 11452
rect 5702 11396 5758 11452
rect 5758 11396 5762 11452
rect 5698 11392 5762 11396
rect 5778 11452 5842 11456
rect 5778 11396 5782 11452
rect 5782 11396 5838 11452
rect 5838 11396 5842 11452
rect 5778 11392 5842 11396
rect 5858 11452 5922 11456
rect 5858 11396 5862 11452
rect 5862 11396 5918 11452
rect 5918 11396 5922 11452
rect 5858 11392 5922 11396
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 3285 10908 3349 10912
rect 3285 10852 3289 10908
rect 3289 10852 3345 10908
rect 3345 10852 3349 10908
rect 3285 10848 3349 10852
rect 3365 10908 3429 10912
rect 3365 10852 3369 10908
rect 3369 10852 3425 10908
rect 3425 10852 3429 10908
rect 3365 10848 3429 10852
rect 3445 10908 3509 10912
rect 3445 10852 3449 10908
rect 3449 10852 3505 10908
rect 3505 10852 3509 10908
rect 3445 10848 3509 10852
rect 3525 10908 3589 10912
rect 3525 10852 3529 10908
rect 3529 10852 3585 10908
rect 3585 10852 3589 10908
rect 3525 10848 3589 10852
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 5618 10364 5682 10368
rect 5618 10308 5622 10364
rect 5622 10308 5678 10364
rect 5678 10308 5682 10364
rect 5618 10304 5682 10308
rect 5698 10364 5762 10368
rect 5698 10308 5702 10364
rect 5702 10308 5758 10364
rect 5758 10308 5762 10364
rect 5698 10304 5762 10308
rect 5778 10364 5842 10368
rect 5778 10308 5782 10364
rect 5782 10308 5838 10364
rect 5838 10308 5842 10364
rect 5778 10304 5842 10308
rect 5858 10364 5922 10368
rect 5858 10308 5862 10364
rect 5862 10308 5918 10364
rect 5918 10308 5922 10364
rect 5858 10304 5922 10308
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 3285 9820 3349 9824
rect 3285 9764 3289 9820
rect 3289 9764 3345 9820
rect 3345 9764 3349 9820
rect 3285 9760 3349 9764
rect 3365 9820 3429 9824
rect 3365 9764 3369 9820
rect 3369 9764 3425 9820
rect 3425 9764 3429 9820
rect 3365 9760 3429 9764
rect 3445 9820 3509 9824
rect 3445 9764 3449 9820
rect 3449 9764 3505 9820
rect 3505 9764 3509 9820
rect 3445 9760 3509 9764
rect 3525 9820 3589 9824
rect 3525 9764 3529 9820
rect 3529 9764 3585 9820
rect 3585 9764 3589 9820
rect 3525 9760 3589 9764
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 5618 9276 5682 9280
rect 5618 9220 5622 9276
rect 5622 9220 5678 9276
rect 5678 9220 5682 9276
rect 5618 9216 5682 9220
rect 5698 9276 5762 9280
rect 5698 9220 5702 9276
rect 5702 9220 5758 9276
rect 5758 9220 5762 9276
rect 5698 9216 5762 9220
rect 5778 9276 5842 9280
rect 5778 9220 5782 9276
rect 5782 9220 5838 9276
rect 5838 9220 5842 9276
rect 5778 9216 5842 9220
rect 5858 9276 5922 9280
rect 5858 9220 5862 9276
rect 5862 9220 5918 9276
rect 5918 9220 5922 9276
rect 5858 9216 5922 9220
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 3285 8732 3349 8736
rect 3285 8676 3289 8732
rect 3289 8676 3345 8732
rect 3345 8676 3349 8732
rect 3285 8672 3349 8676
rect 3365 8732 3429 8736
rect 3365 8676 3369 8732
rect 3369 8676 3425 8732
rect 3425 8676 3429 8732
rect 3365 8672 3429 8676
rect 3445 8732 3509 8736
rect 3445 8676 3449 8732
rect 3449 8676 3505 8732
rect 3505 8676 3509 8732
rect 3445 8672 3509 8676
rect 3525 8732 3589 8736
rect 3525 8676 3529 8732
rect 3529 8676 3585 8732
rect 3585 8676 3589 8732
rect 3525 8672 3589 8676
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 5618 8188 5682 8192
rect 5618 8132 5622 8188
rect 5622 8132 5678 8188
rect 5678 8132 5682 8188
rect 5618 8128 5682 8132
rect 5698 8188 5762 8192
rect 5698 8132 5702 8188
rect 5702 8132 5758 8188
rect 5758 8132 5762 8188
rect 5698 8128 5762 8132
rect 5778 8188 5842 8192
rect 5778 8132 5782 8188
rect 5782 8132 5838 8188
rect 5838 8132 5842 8188
rect 5778 8128 5842 8132
rect 5858 8188 5922 8192
rect 5858 8132 5862 8188
rect 5862 8132 5918 8188
rect 5918 8132 5922 8188
rect 5858 8128 5922 8132
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 3285 7644 3349 7648
rect 3285 7588 3289 7644
rect 3289 7588 3345 7644
rect 3345 7588 3349 7644
rect 3285 7584 3349 7588
rect 3365 7644 3429 7648
rect 3365 7588 3369 7644
rect 3369 7588 3425 7644
rect 3425 7588 3429 7644
rect 3365 7584 3429 7588
rect 3445 7644 3509 7648
rect 3445 7588 3449 7644
rect 3449 7588 3505 7644
rect 3505 7588 3509 7644
rect 3445 7584 3509 7588
rect 3525 7644 3589 7648
rect 3525 7588 3529 7644
rect 3529 7588 3585 7644
rect 3585 7588 3589 7644
rect 3525 7584 3589 7588
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 5618 7100 5682 7104
rect 5618 7044 5622 7100
rect 5622 7044 5678 7100
rect 5678 7044 5682 7100
rect 5618 7040 5682 7044
rect 5698 7100 5762 7104
rect 5698 7044 5702 7100
rect 5702 7044 5758 7100
rect 5758 7044 5762 7100
rect 5698 7040 5762 7044
rect 5778 7100 5842 7104
rect 5778 7044 5782 7100
rect 5782 7044 5838 7100
rect 5838 7044 5842 7100
rect 5778 7040 5842 7044
rect 5858 7100 5922 7104
rect 5858 7044 5862 7100
rect 5862 7044 5918 7100
rect 5918 7044 5922 7100
rect 5858 7040 5922 7044
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 3285 6556 3349 6560
rect 3285 6500 3289 6556
rect 3289 6500 3345 6556
rect 3345 6500 3349 6556
rect 3285 6496 3349 6500
rect 3365 6556 3429 6560
rect 3365 6500 3369 6556
rect 3369 6500 3425 6556
rect 3425 6500 3429 6556
rect 3365 6496 3429 6500
rect 3445 6556 3509 6560
rect 3445 6500 3449 6556
rect 3449 6500 3505 6556
rect 3505 6500 3509 6556
rect 3445 6496 3509 6500
rect 3525 6556 3589 6560
rect 3525 6500 3529 6556
rect 3529 6500 3585 6556
rect 3585 6500 3589 6556
rect 3525 6496 3589 6500
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 5618 6012 5682 6016
rect 5618 5956 5622 6012
rect 5622 5956 5678 6012
rect 5678 5956 5682 6012
rect 5618 5952 5682 5956
rect 5698 6012 5762 6016
rect 5698 5956 5702 6012
rect 5702 5956 5758 6012
rect 5758 5956 5762 6012
rect 5698 5952 5762 5956
rect 5778 6012 5842 6016
rect 5778 5956 5782 6012
rect 5782 5956 5838 6012
rect 5838 5956 5842 6012
rect 5778 5952 5842 5956
rect 5858 6012 5922 6016
rect 5858 5956 5862 6012
rect 5862 5956 5918 6012
rect 5918 5956 5922 6012
rect 5858 5952 5922 5956
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 3285 5468 3349 5472
rect 3285 5412 3289 5468
rect 3289 5412 3345 5468
rect 3345 5412 3349 5468
rect 3285 5408 3349 5412
rect 3365 5468 3429 5472
rect 3365 5412 3369 5468
rect 3369 5412 3425 5468
rect 3425 5412 3429 5468
rect 3365 5408 3429 5412
rect 3445 5468 3509 5472
rect 3445 5412 3449 5468
rect 3449 5412 3505 5468
rect 3505 5412 3509 5468
rect 3445 5408 3509 5412
rect 3525 5468 3589 5472
rect 3525 5412 3529 5468
rect 3529 5412 3585 5468
rect 3585 5412 3589 5468
rect 3525 5408 3589 5412
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 5618 4924 5682 4928
rect 5618 4868 5622 4924
rect 5622 4868 5678 4924
rect 5678 4868 5682 4924
rect 5618 4864 5682 4868
rect 5698 4924 5762 4928
rect 5698 4868 5702 4924
rect 5702 4868 5758 4924
rect 5758 4868 5762 4924
rect 5698 4864 5762 4868
rect 5778 4924 5842 4928
rect 5778 4868 5782 4924
rect 5782 4868 5838 4924
rect 5838 4868 5842 4924
rect 5778 4864 5842 4868
rect 5858 4924 5922 4928
rect 5858 4868 5862 4924
rect 5862 4868 5918 4924
rect 5918 4868 5922 4924
rect 5858 4864 5922 4868
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 3285 4380 3349 4384
rect 3285 4324 3289 4380
rect 3289 4324 3345 4380
rect 3345 4324 3349 4380
rect 3285 4320 3349 4324
rect 3365 4380 3429 4384
rect 3365 4324 3369 4380
rect 3369 4324 3425 4380
rect 3425 4324 3429 4380
rect 3365 4320 3429 4324
rect 3445 4380 3509 4384
rect 3445 4324 3449 4380
rect 3449 4324 3505 4380
rect 3505 4324 3509 4380
rect 3445 4320 3509 4324
rect 3525 4380 3589 4384
rect 3525 4324 3529 4380
rect 3529 4324 3585 4380
rect 3585 4324 3589 4380
rect 3525 4320 3589 4324
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 5618 3836 5682 3840
rect 5618 3780 5622 3836
rect 5622 3780 5678 3836
rect 5678 3780 5682 3836
rect 5618 3776 5682 3780
rect 5698 3836 5762 3840
rect 5698 3780 5702 3836
rect 5702 3780 5758 3836
rect 5758 3780 5762 3836
rect 5698 3776 5762 3780
rect 5778 3836 5842 3840
rect 5778 3780 5782 3836
rect 5782 3780 5838 3836
rect 5838 3780 5842 3836
rect 5778 3776 5842 3780
rect 5858 3836 5922 3840
rect 5858 3780 5862 3836
rect 5862 3780 5918 3836
rect 5918 3780 5922 3836
rect 5858 3776 5922 3780
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 3285 3292 3349 3296
rect 3285 3236 3289 3292
rect 3289 3236 3345 3292
rect 3345 3236 3349 3292
rect 3285 3232 3349 3236
rect 3365 3292 3429 3296
rect 3365 3236 3369 3292
rect 3369 3236 3425 3292
rect 3425 3236 3429 3292
rect 3365 3232 3429 3236
rect 3445 3292 3509 3296
rect 3445 3236 3449 3292
rect 3449 3236 3505 3292
rect 3505 3236 3509 3292
rect 3445 3232 3509 3236
rect 3525 3292 3589 3296
rect 3525 3236 3529 3292
rect 3529 3236 3585 3292
rect 3585 3236 3589 3292
rect 3525 3232 3589 3236
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 5618 2748 5682 2752
rect 5618 2692 5622 2748
rect 5622 2692 5678 2748
rect 5678 2692 5682 2748
rect 5618 2688 5682 2692
rect 5698 2748 5762 2752
rect 5698 2692 5702 2748
rect 5702 2692 5758 2748
rect 5758 2692 5762 2748
rect 5698 2688 5762 2692
rect 5778 2748 5842 2752
rect 5778 2692 5782 2748
rect 5782 2692 5838 2748
rect 5838 2692 5842 2748
rect 5778 2688 5842 2692
rect 5858 2748 5922 2752
rect 5858 2692 5862 2748
rect 5862 2692 5918 2748
rect 5918 2692 5922 2748
rect 5858 2688 5922 2692
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 3285 2204 3349 2208
rect 3285 2148 3289 2204
rect 3289 2148 3345 2204
rect 3345 2148 3349 2204
rect 3285 2144 3349 2148
rect 3365 2204 3429 2208
rect 3365 2148 3369 2204
rect 3369 2148 3425 2204
rect 3425 2148 3429 2204
rect 3365 2144 3429 2148
rect 3445 2204 3509 2208
rect 3445 2148 3449 2204
rect 3449 2148 3505 2204
rect 3505 2148 3509 2204
rect 3445 2144 3509 2148
rect 3525 2204 3589 2208
rect 3525 2148 3529 2204
rect 3529 2148 3585 2204
rect 3585 2148 3589 2204
rect 3525 2144 3589 2148
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
<< metal4 >>
rect 3277 106656 3597 106672
rect 3277 106592 3285 106656
rect 3349 106592 3365 106656
rect 3429 106592 3445 106656
rect 3509 106592 3525 106656
rect 3589 106592 3597 106656
rect 3277 105568 3597 106592
rect 3277 105504 3285 105568
rect 3349 105504 3365 105568
rect 3429 105504 3445 105568
rect 3509 105504 3525 105568
rect 3589 105504 3597 105568
rect 3277 104480 3597 105504
rect 3277 104416 3285 104480
rect 3349 104416 3365 104480
rect 3429 104416 3445 104480
rect 3509 104416 3525 104480
rect 3589 104416 3597 104480
rect 3277 103392 3597 104416
rect 3277 103328 3285 103392
rect 3349 103328 3365 103392
rect 3429 103328 3445 103392
rect 3509 103328 3525 103392
rect 3589 103328 3597 103392
rect 3277 102304 3597 103328
rect 3277 102240 3285 102304
rect 3349 102240 3365 102304
rect 3429 102240 3445 102304
rect 3509 102240 3525 102304
rect 3589 102240 3597 102304
rect 3277 101216 3597 102240
rect 3277 101152 3285 101216
rect 3349 101152 3365 101216
rect 3429 101152 3445 101216
rect 3509 101152 3525 101216
rect 3589 101152 3597 101216
rect 3277 100128 3597 101152
rect 3277 100064 3285 100128
rect 3349 100064 3365 100128
rect 3429 100064 3445 100128
rect 3509 100064 3525 100128
rect 3589 100064 3597 100128
rect 3277 99040 3597 100064
rect 3277 98976 3285 99040
rect 3349 98976 3365 99040
rect 3429 98976 3445 99040
rect 3509 98976 3525 99040
rect 3589 98976 3597 99040
rect 3277 97952 3597 98976
rect 3277 97888 3285 97952
rect 3349 97888 3365 97952
rect 3429 97888 3445 97952
rect 3509 97888 3525 97952
rect 3589 97888 3597 97952
rect 3277 96864 3597 97888
rect 3277 96800 3285 96864
rect 3349 96800 3365 96864
rect 3429 96800 3445 96864
rect 3509 96800 3525 96864
rect 3589 96800 3597 96864
rect 3277 95776 3597 96800
rect 3277 95712 3285 95776
rect 3349 95712 3365 95776
rect 3429 95712 3445 95776
rect 3509 95712 3525 95776
rect 3589 95712 3597 95776
rect 3277 94688 3597 95712
rect 3277 94624 3285 94688
rect 3349 94624 3365 94688
rect 3429 94624 3445 94688
rect 3509 94624 3525 94688
rect 3589 94624 3597 94688
rect 3277 93600 3597 94624
rect 3277 93536 3285 93600
rect 3349 93536 3365 93600
rect 3429 93536 3445 93600
rect 3509 93536 3525 93600
rect 3589 93536 3597 93600
rect 3277 92512 3597 93536
rect 3277 92448 3285 92512
rect 3349 92448 3365 92512
rect 3429 92448 3445 92512
rect 3509 92448 3525 92512
rect 3589 92448 3597 92512
rect 3277 91424 3597 92448
rect 3277 91360 3285 91424
rect 3349 91360 3365 91424
rect 3429 91360 3445 91424
rect 3509 91360 3525 91424
rect 3589 91360 3597 91424
rect 3277 90336 3597 91360
rect 3277 90272 3285 90336
rect 3349 90272 3365 90336
rect 3429 90272 3445 90336
rect 3509 90272 3525 90336
rect 3589 90272 3597 90336
rect 3277 89248 3597 90272
rect 3277 89184 3285 89248
rect 3349 89184 3365 89248
rect 3429 89184 3445 89248
rect 3509 89184 3525 89248
rect 3589 89184 3597 89248
rect 3277 88160 3597 89184
rect 3277 88096 3285 88160
rect 3349 88096 3365 88160
rect 3429 88096 3445 88160
rect 3509 88096 3525 88160
rect 3589 88096 3597 88160
rect 3277 87072 3597 88096
rect 3277 87008 3285 87072
rect 3349 87008 3365 87072
rect 3429 87008 3445 87072
rect 3509 87008 3525 87072
rect 3589 87008 3597 87072
rect 3277 85984 3597 87008
rect 3277 85920 3285 85984
rect 3349 85920 3365 85984
rect 3429 85920 3445 85984
rect 3509 85920 3525 85984
rect 3589 85920 3597 85984
rect 3277 84896 3597 85920
rect 3277 84832 3285 84896
rect 3349 84832 3365 84896
rect 3429 84832 3445 84896
rect 3509 84832 3525 84896
rect 3589 84832 3597 84896
rect 3277 83808 3597 84832
rect 3277 83744 3285 83808
rect 3349 83744 3365 83808
rect 3429 83744 3445 83808
rect 3509 83744 3525 83808
rect 3589 83744 3597 83808
rect 3277 82720 3597 83744
rect 3277 82656 3285 82720
rect 3349 82656 3365 82720
rect 3429 82656 3445 82720
rect 3509 82656 3525 82720
rect 3589 82656 3597 82720
rect 3277 81632 3597 82656
rect 3277 81568 3285 81632
rect 3349 81568 3365 81632
rect 3429 81568 3445 81632
rect 3509 81568 3525 81632
rect 3589 81568 3597 81632
rect 3277 80544 3597 81568
rect 3277 80480 3285 80544
rect 3349 80480 3365 80544
rect 3429 80480 3445 80544
rect 3509 80480 3525 80544
rect 3589 80480 3597 80544
rect 3277 79456 3597 80480
rect 3277 79392 3285 79456
rect 3349 79392 3365 79456
rect 3429 79392 3445 79456
rect 3509 79392 3525 79456
rect 3589 79392 3597 79456
rect 3277 78368 3597 79392
rect 3277 78304 3285 78368
rect 3349 78304 3365 78368
rect 3429 78304 3445 78368
rect 3509 78304 3525 78368
rect 3589 78304 3597 78368
rect 3277 77280 3597 78304
rect 3277 77216 3285 77280
rect 3349 77216 3365 77280
rect 3429 77216 3445 77280
rect 3509 77216 3525 77280
rect 3589 77216 3597 77280
rect 3277 76192 3597 77216
rect 3277 76128 3285 76192
rect 3349 76128 3365 76192
rect 3429 76128 3445 76192
rect 3509 76128 3525 76192
rect 3589 76128 3597 76192
rect 3277 75104 3597 76128
rect 3277 75040 3285 75104
rect 3349 75040 3365 75104
rect 3429 75040 3445 75104
rect 3509 75040 3525 75104
rect 3589 75040 3597 75104
rect 3277 74016 3597 75040
rect 3277 73952 3285 74016
rect 3349 73952 3365 74016
rect 3429 73952 3445 74016
rect 3509 73952 3525 74016
rect 3589 73952 3597 74016
rect 3277 72928 3597 73952
rect 3277 72864 3285 72928
rect 3349 72864 3365 72928
rect 3429 72864 3445 72928
rect 3509 72864 3525 72928
rect 3589 72864 3597 72928
rect 3277 71840 3597 72864
rect 3277 71776 3285 71840
rect 3349 71776 3365 71840
rect 3429 71776 3445 71840
rect 3509 71776 3525 71840
rect 3589 71776 3597 71840
rect 3277 70752 3597 71776
rect 3277 70688 3285 70752
rect 3349 70688 3365 70752
rect 3429 70688 3445 70752
rect 3509 70688 3525 70752
rect 3589 70688 3597 70752
rect 3277 69664 3597 70688
rect 3277 69600 3285 69664
rect 3349 69600 3365 69664
rect 3429 69600 3445 69664
rect 3509 69600 3525 69664
rect 3589 69600 3597 69664
rect 3277 68576 3597 69600
rect 3277 68512 3285 68576
rect 3349 68512 3365 68576
rect 3429 68512 3445 68576
rect 3509 68512 3525 68576
rect 3589 68512 3597 68576
rect 3277 67488 3597 68512
rect 3277 67424 3285 67488
rect 3349 67424 3365 67488
rect 3429 67424 3445 67488
rect 3509 67424 3525 67488
rect 3589 67424 3597 67488
rect 3277 66400 3597 67424
rect 3277 66336 3285 66400
rect 3349 66336 3365 66400
rect 3429 66336 3445 66400
rect 3509 66336 3525 66400
rect 3589 66336 3597 66400
rect 3277 65312 3597 66336
rect 3277 65248 3285 65312
rect 3349 65248 3365 65312
rect 3429 65248 3445 65312
rect 3509 65248 3525 65312
rect 3589 65248 3597 65312
rect 3277 64224 3597 65248
rect 3277 64160 3285 64224
rect 3349 64160 3365 64224
rect 3429 64160 3445 64224
rect 3509 64160 3525 64224
rect 3589 64160 3597 64224
rect 3277 63136 3597 64160
rect 3277 63072 3285 63136
rect 3349 63072 3365 63136
rect 3429 63072 3445 63136
rect 3509 63072 3525 63136
rect 3589 63072 3597 63136
rect 3277 62048 3597 63072
rect 3277 61984 3285 62048
rect 3349 61984 3365 62048
rect 3429 61984 3445 62048
rect 3509 61984 3525 62048
rect 3589 61984 3597 62048
rect 3277 60960 3597 61984
rect 3277 60896 3285 60960
rect 3349 60896 3365 60960
rect 3429 60896 3445 60960
rect 3509 60896 3525 60960
rect 3589 60896 3597 60960
rect 3277 59872 3597 60896
rect 3277 59808 3285 59872
rect 3349 59808 3365 59872
rect 3429 59808 3445 59872
rect 3509 59808 3525 59872
rect 3589 59808 3597 59872
rect 3277 58784 3597 59808
rect 3277 58720 3285 58784
rect 3349 58720 3365 58784
rect 3429 58720 3445 58784
rect 3509 58720 3525 58784
rect 3589 58720 3597 58784
rect 3277 57696 3597 58720
rect 3277 57632 3285 57696
rect 3349 57632 3365 57696
rect 3429 57632 3445 57696
rect 3509 57632 3525 57696
rect 3589 57632 3597 57696
rect 3277 56608 3597 57632
rect 3277 56544 3285 56608
rect 3349 56544 3365 56608
rect 3429 56544 3445 56608
rect 3509 56544 3525 56608
rect 3589 56544 3597 56608
rect 3277 55520 3597 56544
rect 3277 55456 3285 55520
rect 3349 55456 3365 55520
rect 3429 55456 3445 55520
rect 3509 55456 3525 55520
rect 3589 55456 3597 55520
rect 3277 54432 3597 55456
rect 3277 54368 3285 54432
rect 3349 54368 3365 54432
rect 3429 54368 3445 54432
rect 3509 54368 3525 54432
rect 3589 54368 3597 54432
rect 3277 53344 3597 54368
rect 3277 53280 3285 53344
rect 3349 53280 3365 53344
rect 3429 53280 3445 53344
rect 3509 53280 3525 53344
rect 3589 53280 3597 53344
rect 3277 52256 3597 53280
rect 3277 52192 3285 52256
rect 3349 52192 3365 52256
rect 3429 52192 3445 52256
rect 3509 52192 3525 52256
rect 3589 52192 3597 52256
rect 3277 51168 3597 52192
rect 3277 51104 3285 51168
rect 3349 51104 3365 51168
rect 3429 51104 3445 51168
rect 3509 51104 3525 51168
rect 3589 51104 3597 51168
rect 3277 50080 3597 51104
rect 3277 50016 3285 50080
rect 3349 50016 3365 50080
rect 3429 50016 3445 50080
rect 3509 50016 3525 50080
rect 3589 50016 3597 50080
rect 3277 48992 3597 50016
rect 3277 48928 3285 48992
rect 3349 48928 3365 48992
rect 3429 48928 3445 48992
rect 3509 48928 3525 48992
rect 3589 48928 3597 48992
rect 3277 47904 3597 48928
rect 3277 47840 3285 47904
rect 3349 47840 3365 47904
rect 3429 47840 3445 47904
rect 3509 47840 3525 47904
rect 3589 47840 3597 47904
rect 3277 46816 3597 47840
rect 3277 46752 3285 46816
rect 3349 46752 3365 46816
rect 3429 46752 3445 46816
rect 3509 46752 3525 46816
rect 3589 46752 3597 46816
rect 3277 45728 3597 46752
rect 3277 45664 3285 45728
rect 3349 45664 3365 45728
rect 3429 45664 3445 45728
rect 3509 45664 3525 45728
rect 3589 45664 3597 45728
rect 3277 44640 3597 45664
rect 3277 44576 3285 44640
rect 3349 44576 3365 44640
rect 3429 44576 3445 44640
rect 3509 44576 3525 44640
rect 3589 44576 3597 44640
rect 3277 43552 3597 44576
rect 3277 43488 3285 43552
rect 3349 43488 3365 43552
rect 3429 43488 3445 43552
rect 3509 43488 3525 43552
rect 3589 43488 3597 43552
rect 3277 42464 3597 43488
rect 3277 42400 3285 42464
rect 3349 42400 3365 42464
rect 3429 42400 3445 42464
rect 3509 42400 3525 42464
rect 3589 42400 3597 42464
rect 3277 41376 3597 42400
rect 3277 41312 3285 41376
rect 3349 41312 3365 41376
rect 3429 41312 3445 41376
rect 3509 41312 3525 41376
rect 3589 41312 3597 41376
rect 3277 40288 3597 41312
rect 3277 40224 3285 40288
rect 3349 40224 3365 40288
rect 3429 40224 3445 40288
rect 3509 40224 3525 40288
rect 3589 40224 3597 40288
rect 3277 39200 3597 40224
rect 3277 39136 3285 39200
rect 3349 39136 3365 39200
rect 3429 39136 3445 39200
rect 3509 39136 3525 39200
rect 3589 39136 3597 39200
rect 3277 38112 3597 39136
rect 3277 38048 3285 38112
rect 3349 38048 3365 38112
rect 3429 38048 3445 38112
rect 3509 38048 3525 38112
rect 3589 38048 3597 38112
rect 3277 37024 3597 38048
rect 3277 36960 3285 37024
rect 3349 36960 3365 37024
rect 3429 36960 3445 37024
rect 3509 36960 3525 37024
rect 3589 36960 3597 37024
rect 3277 35936 3597 36960
rect 3277 35872 3285 35936
rect 3349 35872 3365 35936
rect 3429 35872 3445 35936
rect 3509 35872 3525 35936
rect 3589 35872 3597 35936
rect 3277 34848 3597 35872
rect 3277 34784 3285 34848
rect 3349 34784 3365 34848
rect 3429 34784 3445 34848
rect 3509 34784 3525 34848
rect 3589 34784 3597 34848
rect 3277 33760 3597 34784
rect 3277 33696 3285 33760
rect 3349 33696 3365 33760
rect 3429 33696 3445 33760
rect 3509 33696 3525 33760
rect 3589 33696 3597 33760
rect 3277 32672 3597 33696
rect 3277 32608 3285 32672
rect 3349 32608 3365 32672
rect 3429 32608 3445 32672
rect 3509 32608 3525 32672
rect 3589 32608 3597 32672
rect 3277 31584 3597 32608
rect 3277 31520 3285 31584
rect 3349 31520 3365 31584
rect 3429 31520 3445 31584
rect 3509 31520 3525 31584
rect 3589 31520 3597 31584
rect 3277 30496 3597 31520
rect 3277 30432 3285 30496
rect 3349 30432 3365 30496
rect 3429 30432 3445 30496
rect 3509 30432 3525 30496
rect 3589 30432 3597 30496
rect 3277 29408 3597 30432
rect 3277 29344 3285 29408
rect 3349 29344 3365 29408
rect 3429 29344 3445 29408
rect 3509 29344 3525 29408
rect 3589 29344 3597 29408
rect 3277 28320 3597 29344
rect 3277 28256 3285 28320
rect 3349 28256 3365 28320
rect 3429 28256 3445 28320
rect 3509 28256 3525 28320
rect 3589 28256 3597 28320
rect 3277 27232 3597 28256
rect 3277 27168 3285 27232
rect 3349 27168 3365 27232
rect 3429 27168 3445 27232
rect 3509 27168 3525 27232
rect 3589 27168 3597 27232
rect 3277 26144 3597 27168
rect 3277 26080 3285 26144
rect 3349 26080 3365 26144
rect 3429 26080 3445 26144
rect 3509 26080 3525 26144
rect 3589 26080 3597 26144
rect 3277 25056 3597 26080
rect 3277 24992 3285 25056
rect 3349 24992 3365 25056
rect 3429 24992 3445 25056
rect 3509 24992 3525 25056
rect 3589 24992 3597 25056
rect 3277 23968 3597 24992
rect 3277 23904 3285 23968
rect 3349 23904 3365 23968
rect 3429 23904 3445 23968
rect 3509 23904 3525 23968
rect 3589 23904 3597 23968
rect 3277 22880 3597 23904
rect 3277 22816 3285 22880
rect 3349 22816 3365 22880
rect 3429 22816 3445 22880
rect 3509 22816 3525 22880
rect 3589 22816 3597 22880
rect 3277 21792 3597 22816
rect 3277 21728 3285 21792
rect 3349 21728 3365 21792
rect 3429 21728 3445 21792
rect 3509 21728 3525 21792
rect 3589 21728 3597 21792
rect 3277 20704 3597 21728
rect 3277 20640 3285 20704
rect 3349 20640 3365 20704
rect 3429 20640 3445 20704
rect 3509 20640 3525 20704
rect 3589 20640 3597 20704
rect 3277 19616 3597 20640
rect 3277 19552 3285 19616
rect 3349 19552 3365 19616
rect 3429 19552 3445 19616
rect 3509 19552 3525 19616
rect 3589 19552 3597 19616
rect 3277 18528 3597 19552
rect 3277 18464 3285 18528
rect 3349 18464 3365 18528
rect 3429 18464 3445 18528
rect 3509 18464 3525 18528
rect 3589 18464 3597 18528
rect 3277 17440 3597 18464
rect 3277 17376 3285 17440
rect 3349 17376 3365 17440
rect 3429 17376 3445 17440
rect 3509 17376 3525 17440
rect 3589 17376 3597 17440
rect 3277 16352 3597 17376
rect 3277 16288 3285 16352
rect 3349 16288 3365 16352
rect 3429 16288 3445 16352
rect 3509 16288 3525 16352
rect 3589 16288 3597 16352
rect 3277 15264 3597 16288
rect 3277 15200 3285 15264
rect 3349 15200 3365 15264
rect 3429 15200 3445 15264
rect 3509 15200 3525 15264
rect 3589 15200 3597 15264
rect 3277 14176 3597 15200
rect 3277 14112 3285 14176
rect 3349 14112 3365 14176
rect 3429 14112 3445 14176
rect 3509 14112 3525 14176
rect 3589 14112 3597 14176
rect 3277 13088 3597 14112
rect 3277 13024 3285 13088
rect 3349 13024 3365 13088
rect 3429 13024 3445 13088
rect 3509 13024 3525 13088
rect 3589 13024 3597 13088
rect 3277 12000 3597 13024
rect 3277 11936 3285 12000
rect 3349 11936 3365 12000
rect 3429 11936 3445 12000
rect 3509 11936 3525 12000
rect 3589 11936 3597 12000
rect 3277 10912 3597 11936
rect 3277 10848 3285 10912
rect 3349 10848 3365 10912
rect 3429 10848 3445 10912
rect 3509 10848 3525 10912
rect 3589 10848 3597 10912
rect 3277 9824 3597 10848
rect 3277 9760 3285 9824
rect 3349 9760 3365 9824
rect 3429 9760 3445 9824
rect 3509 9760 3525 9824
rect 3589 9760 3597 9824
rect 3277 8736 3597 9760
rect 3277 8672 3285 8736
rect 3349 8672 3365 8736
rect 3429 8672 3445 8736
rect 3509 8672 3525 8736
rect 3589 8672 3597 8736
rect 3277 7648 3597 8672
rect 3277 7584 3285 7648
rect 3349 7584 3365 7648
rect 3429 7584 3445 7648
rect 3509 7584 3525 7648
rect 3589 7584 3597 7648
rect 3277 6560 3597 7584
rect 3277 6496 3285 6560
rect 3349 6496 3365 6560
rect 3429 6496 3445 6560
rect 3509 6496 3525 6560
rect 3589 6496 3597 6560
rect 3277 5472 3597 6496
rect 3277 5408 3285 5472
rect 3349 5408 3365 5472
rect 3429 5408 3445 5472
rect 3509 5408 3525 5472
rect 3589 5408 3597 5472
rect 3277 4384 3597 5408
rect 3277 4320 3285 4384
rect 3349 4320 3365 4384
rect 3429 4320 3445 4384
rect 3509 4320 3525 4384
rect 3589 4320 3597 4384
rect 3277 3296 3597 4320
rect 3277 3232 3285 3296
rect 3349 3232 3365 3296
rect 3429 3232 3445 3296
rect 3509 3232 3525 3296
rect 3589 3232 3597 3296
rect 3277 2208 3597 3232
rect 3277 2144 3285 2208
rect 3349 2144 3365 2208
rect 3429 2144 3445 2208
rect 3509 2144 3525 2208
rect 3589 2144 3597 2208
rect 3277 2128 3597 2144
rect 5610 106112 5931 106672
rect 5610 106048 5618 106112
rect 5682 106048 5698 106112
rect 5762 106048 5778 106112
rect 5842 106048 5858 106112
rect 5922 106048 5931 106112
rect 5610 105024 5931 106048
rect 5610 104960 5618 105024
rect 5682 104960 5698 105024
rect 5762 104960 5778 105024
rect 5842 104960 5858 105024
rect 5922 104960 5931 105024
rect 5610 103936 5931 104960
rect 5610 103872 5618 103936
rect 5682 103872 5698 103936
rect 5762 103872 5778 103936
rect 5842 103872 5858 103936
rect 5922 103872 5931 103936
rect 5610 102848 5931 103872
rect 5610 102784 5618 102848
rect 5682 102784 5698 102848
rect 5762 102784 5778 102848
rect 5842 102784 5858 102848
rect 5922 102784 5931 102848
rect 5610 101760 5931 102784
rect 5610 101696 5618 101760
rect 5682 101696 5698 101760
rect 5762 101696 5778 101760
rect 5842 101696 5858 101760
rect 5922 101696 5931 101760
rect 5610 100672 5931 101696
rect 5610 100608 5618 100672
rect 5682 100608 5698 100672
rect 5762 100608 5778 100672
rect 5842 100608 5858 100672
rect 5922 100608 5931 100672
rect 5610 99584 5931 100608
rect 5610 99520 5618 99584
rect 5682 99520 5698 99584
rect 5762 99520 5778 99584
rect 5842 99520 5858 99584
rect 5922 99520 5931 99584
rect 5610 98496 5931 99520
rect 5610 98432 5618 98496
rect 5682 98432 5698 98496
rect 5762 98432 5778 98496
rect 5842 98432 5858 98496
rect 5922 98432 5931 98496
rect 5610 97408 5931 98432
rect 5610 97344 5618 97408
rect 5682 97344 5698 97408
rect 5762 97344 5778 97408
rect 5842 97344 5858 97408
rect 5922 97344 5931 97408
rect 5610 96320 5931 97344
rect 5610 96256 5618 96320
rect 5682 96256 5698 96320
rect 5762 96256 5778 96320
rect 5842 96256 5858 96320
rect 5922 96256 5931 96320
rect 5610 95232 5931 96256
rect 5610 95168 5618 95232
rect 5682 95168 5698 95232
rect 5762 95168 5778 95232
rect 5842 95168 5858 95232
rect 5922 95168 5931 95232
rect 5610 94144 5931 95168
rect 5610 94080 5618 94144
rect 5682 94080 5698 94144
rect 5762 94080 5778 94144
rect 5842 94080 5858 94144
rect 5922 94080 5931 94144
rect 5610 93056 5931 94080
rect 5610 92992 5618 93056
rect 5682 92992 5698 93056
rect 5762 92992 5778 93056
rect 5842 92992 5858 93056
rect 5922 92992 5931 93056
rect 5610 91968 5931 92992
rect 5610 91904 5618 91968
rect 5682 91904 5698 91968
rect 5762 91904 5778 91968
rect 5842 91904 5858 91968
rect 5922 91904 5931 91968
rect 5610 90880 5931 91904
rect 5610 90816 5618 90880
rect 5682 90816 5698 90880
rect 5762 90816 5778 90880
rect 5842 90816 5858 90880
rect 5922 90816 5931 90880
rect 5610 89792 5931 90816
rect 5610 89728 5618 89792
rect 5682 89728 5698 89792
rect 5762 89728 5778 89792
rect 5842 89728 5858 89792
rect 5922 89728 5931 89792
rect 5610 88704 5931 89728
rect 5610 88640 5618 88704
rect 5682 88640 5698 88704
rect 5762 88640 5778 88704
rect 5842 88640 5858 88704
rect 5922 88640 5931 88704
rect 5610 87616 5931 88640
rect 5610 87552 5618 87616
rect 5682 87552 5698 87616
rect 5762 87552 5778 87616
rect 5842 87552 5858 87616
rect 5922 87552 5931 87616
rect 5610 86528 5931 87552
rect 5610 86464 5618 86528
rect 5682 86464 5698 86528
rect 5762 86464 5778 86528
rect 5842 86464 5858 86528
rect 5922 86464 5931 86528
rect 5610 85440 5931 86464
rect 5610 85376 5618 85440
rect 5682 85376 5698 85440
rect 5762 85376 5778 85440
rect 5842 85376 5858 85440
rect 5922 85376 5931 85440
rect 5610 84352 5931 85376
rect 5610 84288 5618 84352
rect 5682 84288 5698 84352
rect 5762 84288 5778 84352
rect 5842 84288 5858 84352
rect 5922 84288 5931 84352
rect 5610 83264 5931 84288
rect 5610 83200 5618 83264
rect 5682 83200 5698 83264
rect 5762 83200 5778 83264
rect 5842 83200 5858 83264
rect 5922 83200 5931 83264
rect 5610 82176 5931 83200
rect 5610 82112 5618 82176
rect 5682 82112 5698 82176
rect 5762 82112 5778 82176
rect 5842 82112 5858 82176
rect 5922 82112 5931 82176
rect 5610 81088 5931 82112
rect 5610 81024 5618 81088
rect 5682 81024 5698 81088
rect 5762 81024 5778 81088
rect 5842 81024 5858 81088
rect 5922 81024 5931 81088
rect 5610 80000 5931 81024
rect 5610 79936 5618 80000
rect 5682 79936 5698 80000
rect 5762 79936 5778 80000
rect 5842 79936 5858 80000
rect 5922 79936 5931 80000
rect 5610 78912 5931 79936
rect 5610 78848 5618 78912
rect 5682 78848 5698 78912
rect 5762 78848 5778 78912
rect 5842 78848 5858 78912
rect 5922 78848 5931 78912
rect 5610 77824 5931 78848
rect 5610 77760 5618 77824
rect 5682 77760 5698 77824
rect 5762 77760 5778 77824
rect 5842 77760 5858 77824
rect 5922 77760 5931 77824
rect 5610 76736 5931 77760
rect 5610 76672 5618 76736
rect 5682 76672 5698 76736
rect 5762 76672 5778 76736
rect 5842 76672 5858 76736
rect 5922 76672 5931 76736
rect 5610 75648 5931 76672
rect 5610 75584 5618 75648
rect 5682 75584 5698 75648
rect 5762 75584 5778 75648
rect 5842 75584 5858 75648
rect 5922 75584 5931 75648
rect 5610 74560 5931 75584
rect 5610 74496 5618 74560
rect 5682 74496 5698 74560
rect 5762 74496 5778 74560
rect 5842 74496 5858 74560
rect 5922 74496 5931 74560
rect 5610 73472 5931 74496
rect 5610 73408 5618 73472
rect 5682 73408 5698 73472
rect 5762 73408 5778 73472
rect 5842 73408 5858 73472
rect 5922 73408 5931 73472
rect 5610 72384 5931 73408
rect 5610 72320 5618 72384
rect 5682 72320 5698 72384
rect 5762 72320 5778 72384
rect 5842 72320 5858 72384
rect 5922 72320 5931 72384
rect 5610 71296 5931 72320
rect 5610 71232 5618 71296
rect 5682 71232 5698 71296
rect 5762 71232 5778 71296
rect 5842 71232 5858 71296
rect 5922 71232 5931 71296
rect 5610 70208 5931 71232
rect 5610 70144 5618 70208
rect 5682 70144 5698 70208
rect 5762 70144 5778 70208
rect 5842 70144 5858 70208
rect 5922 70144 5931 70208
rect 5610 69120 5931 70144
rect 5610 69056 5618 69120
rect 5682 69056 5698 69120
rect 5762 69056 5778 69120
rect 5842 69056 5858 69120
rect 5922 69056 5931 69120
rect 5610 68032 5931 69056
rect 5610 67968 5618 68032
rect 5682 67968 5698 68032
rect 5762 67968 5778 68032
rect 5842 67968 5858 68032
rect 5922 67968 5931 68032
rect 5610 66944 5931 67968
rect 5610 66880 5618 66944
rect 5682 66880 5698 66944
rect 5762 66880 5778 66944
rect 5842 66880 5858 66944
rect 5922 66880 5931 66944
rect 5610 65856 5931 66880
rect 5610 65792 5618 65856
rect 5682 65792 5698 65856
rect 5762 65792 5778 65856
rect 5842 65792 5858 65856
rect 5922 65792 5931 65856
rect 5610 64768 5931 65792
rect 5610 64704 5618 64768
rect 5682 64704 5698 64768
rect 5762 64704 5778 64768
rect 5842 64704 5858 64768
rect 5922 64704 5931 64768
rect 5610 63680 5931 64704
rect 5610 63616 5618 63680
rect 5682 63616 5698 63680
rect 5762 63616 5778 63680
rect 5842 63616 5858 63680
rect 5922 63616 5931 63680
rect 5610 62592 5931 63616
rect 5610 62528 5618 62592
rect 5682 62528 5698 62592
rect 5762 62528 5778 62592
rect 5842 62528 5858 62592
rect 5922 62528 5931 62592
rect 5610 61504 5931 62528
rect 5610 61440 5618 61504
rect 5682 61440 5698 61504
rect 5762 61440 5778 61504
rect 5842 61440 5858 61504
rect 5922 61440 5931 61504
rect 5610 60416 5931 61440
rect 5610 60352 5618 60416
rect 5682 60352 5698 60416
rect 5762 60352 5778 60416
rect 5842 60352 5858 60416
rect 5922 60352 5931 60416
rect 5610 59328 5931 60352
rect 5610 59264 5618 59328
rect 5682 59264 5698 59328
rect 5762 59264 5778 59328
rect 5842 59264 5858 59328
rect 5922 59264 5931 59328
rect 5610 58240 5931 59264
rect 5610 58176 5618 58240
rect 5682 58176 5698 58240
rect 5762 58176 5778 58240
rect 5842 58176 5858 58240
rect 5922 58176 5931 58240
rect 5610 57152 5931 58176
rect 5610 57088 5618 57152
rect 5682 57088 5698 57152
rect 5762 57088 5778 57152
rect 5842 57088 5858 57152
rect 5922 57088 5931 57152
rect 5610 56064 5931 57088
rect 5610 56000 5618 56064
rect 5682 56000 5698 56064
rect 5762 56000 5778 56064
rect 5842 56000 5858 56064
rect 5922 56000 5931 56064
rect 5610 54976 5931 56000
rect 5610 54912 5618 54976
rect 5682 54912 5698 54976
rect 5762 54912 5778 54976
rect 5842 54912 5858 54976
rect 5922 54912 5931 54976
rect 5610 53888 5931 54912
rect 5610 53824 5618 53888
rect 5682 53824 5698 53888
rect 5762 53824 5778 53888
rect 5842 53824 5858 53888
rect 5922 53824 5931 53888
rect 5610 52800 5931 53824
rect 5610 52736 5618 52800
rect 5682 52736 5698 52800
rect 5762 52736 5778 52800
rect 5842 52736 5858 52800
rect 5922 52736 5931 52800
rect 5610 51712 5931 52736
rect 5610 51648 5618 51712
rect 5682 51648 5698 51712
rect 5762 51648 5778 51712
rect 5842 51648 5858 51712
rect 5922 51648 5931 51712
rect 5610 50624 5931 51648
rect 5610 50560 5618 50624
rect 5682 50560 5698 50624
rect 5762 50560 5778 50624
rect 5842 50560 5858 50624
rect 5922 50560 5931 50624
rect 5610 49536 5931 50560
rect 5610 49472 5618 49536
rect 5682 49472 5698 49536
rect 5762 49472 5778 49536
rect 5842 49472 5858 49536
rect 5922 49472 5931 49536
rect 5610 48448 5931 49472
rect 5610 48384 5618 48448
rect 5682 48384 5698 48448
rect 5762 48384 5778 48448
rect 5842 48384 5858 48448
rect 5922 48384 5931 48448
rect 5610 47360 5931 48384
rect 5610 47296 5618 47360
rect 5682 47296 5698 47360
rect 5762 47296 5778 47360
rect 5842 47296 5858 47360
rect 5922 47296 5931 47360
rect 5610 46272 5931 47296
rect 5610 46208 5618 46272
rect 5682 46208 5698 46272
rect 5762 46208 5778 46272
rect 5842 46208 5858 46272
rect 5922 46208 5931 46272
rect 5610 45184 5931 46208
rect 5610 45120 5618 45184
rect 5682 45120 5698 45184
rect 5762 45120 5778 45184
rect 5842 45120 5858 45184
rect 5922 45120 5931 45184
rect 5610 44096 5931 45120
rect 5610 44032 5618 44096
rect 5682 44032 5698 44096
rect 5762 44032 5778 44096
rect 5842 44032 5858 44096
rect 5922 44032 5931 44096
rect 5610 43008 5931 44032
rect 5610 42944 5618 43008
rect 5682 42944 5698 43008
rect 5762 42944 5778 43008
rect 5842 42944 5858 43008
rect 5922 42944 5931 43008
rect 5610 41920 5931 42944
rect 5610 41856 5618 41920
rect 5682 41856 5698 41920
rect 5762 41856 5778 41920
rect 5842 41856 5858 41920
rect 5922 41856 5931 41920
rect 5610 40832 5931 41856
rect 5610 40768 5618 40832
rect 5682 40768 5698 40832
rect 5762 40768 5778 40832
rect 5842 40768 5858 40832
rect 5922 40768 5931 40832
rect 5610 39744 5931 40768
rect 5610 39680 5618 39744
rect 5682 39680 5698 39744
rect 5762 39680 5778 39744
rect 5842 39680 5858 39744
rect 5922 39680 5931 39744
rect 5610 38656 5931 39680
rect 5610 38592 5618 38656
rect 5682 38592 5698 38656
rect 5762 38592 5778 38656
rect 5842 38592 5858 38656
rect 5922 38592 5931 38656
rect 5610 37568 5931 38592
rect 5610 37504 5618 37568
rect 5682 37504 5698 37568
rect 5762 37504 5778 37568
rect 5842 37504 5858 37568
rect 5922 37504 5931 37568
rect 5610 36480 5931 37504
rect 5610 36416 5618 36480
rect 5682 36416 5698 36480
rect 5762 36416 5778 36480
rect 5842 36416 5858 36480
rect 5922 36416 5931 36480
rect 5610 35392 5931 36416
rect 5610 35328 5618 35392
rect 5682 35328 5698 35392
rect 5762 35328 5778 35392
rect 5842 35328 5858 35392
rect 5922 35328 5931 35392
rect 5610 34304 5931 35328
rect 5610 34240 5618 34304
rect 5682 34240 5698 34304
rect 5762 34240 5778 34304
rect 5842 34240 5858 34304
rect 5922 34240 5931 34304
rect 5610 33216 5931 34240
rect 5610 33152 5618 33216
rect 5682 33152 5698 33216
rect 5762 33152 5778 33216
rect 5842 33152 5858 33216
rect 5922 33152 5931 33216
rect 5610 32128 5931 33152
rect 5610 32064 5618 32128
rect 5682 32064 5698 32128
rect 5762 32064 5778 32128
rect 5842 32064 5858 32128
rect 5922 32064 5931 32128
rect 5610 31040 5931 32064
rect 5610 30976 5618 31040
rect 5682 30976 5698 31040
rect 5762 30976 5778 31040
rect 5842 30976 5858 31040
rect 5922 30976 5931 31040
rect 5610 29952 5931 30976
rect 5610 29888 5618 29952
rect 5682 29888 5698 29952
rect 5762 29888 5778 29952
rect 5842 29888 5858 29952
rect 5922 29888 5931 29952
rect 5610 28864 5931 29888
rect 5610 28800 5618 28864
rect 5682 28800 5698 28864
rect 5762 28800 5778 28864
rect 5842 28800 5858 28864
rect 5922 28800 5931 28864
rect 5610 27776 5931 28800
rect 5610 27712 5618 27776
rect 5682 27712 5698 27776
rect 5762 27712 5778 27776
rect 5842 27712 5858 27776
rect 5922 27712 5931 27776
rect 5610 26688 5931 27712
rect 5610 26624 5618 26688
rect 5682 26624 5698 26688
rect 5762 26624 5778 26688
rect 5842 26624 5858 26688
rect 5922 26624 5931 26688
rect 5610 25600 5931 26624
rect 5610 25536 5618 25600
rect 5682 25536 5698 25600
rect 5762 25536 5778 25600
rect 5842 25536 5858 25600
rect 5922 25536 5931 25600
rect 5610 24512 5931 25536
rect 5610 24448 5618 24512
rect 5682 24448 5698 24512
rect 5762 24448 5778 24512
rect 5842 24448 5858 24512
rect 5922 24448 5931 24512
rect 5610 23424 5931 24448
rect 5610 23360 5618 23424
rect 5682 23360 5698 23424
rect 5762 23360 5778 23424
rect 5842 23360 5858 23424
rect 5922 23360 5931 23424
rect 5610 22336 5931 23360
rect 5610 22272 5618 22336
rect 5682 22272 5698 22336
rect 5762 22272 5778 22336
rect 5842 22272 5858 22336
rect 5922 22272 5931 22336
rect 5610 21248 5931 22272
rect 5610 21184 5618 21248
rect 5682 21184 5698 21248
rect 5762 21184 5778 21248
rect 5842 21184 5858 21248
rect 5922 21184 5931 21248
rect 5610 20160 5931 21184
rect 5610 20096 5618 20160
rect 5682 20096 5698 20160
rect 5762 20096 5778 20160
rect 5842 20096 5858 20160
rect 5922 20096 5931 20160
rect 5610 19072 5931 20096
rect 5610 19008 5618 19072
rect 5682 19008 5698 19072
rect 5762 19008 5778 19072
rect 5842 19008 5858 19072
rect 5922 19008 5931 19072
rect 5610 17984 5931 19008
rect 5610 17920 5618 17984
rect 5682 17920 5698 17984
rect 5762 17920 5778 17984
rect 5842 17920 5858 17984
rect 5922 17920 5931 17984
rect 5610 16896 5931 17920
rect 5610 16832 5618 16896
rect 5682 16832 5698 16896
rect 5762 16832 5778 16896
rect 5842 16832 5858 16896
rect 5922 16832 5931 16896
rect 5610 15808 5931 16832
rect 5610 15744 5618 15808
rect 5682 15744 5698 15808
rect 5762 15744 5778 15808
rect 5842 15744 5858 15808
rect 5922 15744 5931 15808
rect 5610 14720 5931 15744
rect 5610 14656 5618 14720
rect 5682 14656 5698 14720
rect 5762 14656 5778 14720
rect 5842 14656 5858 14720
rect 5922 14656 5931 14720
rect 5610 13632 5931 14656
rect 5610 13568 5618 13632
rect 5682 13568 5698 13632
rect 5762 13568 5778 13632
rect 5842 13568 5858 13632
rect 5922 13568 5931 13632
rect 5610 12544 5931 13568
rect 5610 12480 5618 12544
rect 5682 12480 5698 12544
rect 5762 12480 5778 12544
rect 5842 12480 5858 12544
rect 5922 12480 5931 12544
rect 5610 11456 5931 12480
rect 5610 11392 5618 11456
rect 5682 11392 5698 11456
rect 5762 11392 5778 11456
rect 5842 11392 5858 11456
rect 5922 11392 5931 11456
rect 5610 10368 5931 11392
rect 5610 10304 5618 10368
rect 5682 10304 5698 10368
rect 5762 10304 5778 10368
rect 5842 10304 5858 10368
rect 5922 10304 5931 10368
rect 5610 9280 5931 10304
rect 5610 9216 5618 9280
rect 5682 9216 5698 9280
rect 5762 9216 5778 9280
rect 5842 9216 5858 9280
rect 5922 9216 5931 9280
rect 5610 8192 5931 9216
rect 5610 8128 5618 8192
rect 5682 8128 5698 8192
rect 5762 8128 5778 8192
rect 5842 8128 5858 8192
rect 5922 8128 5931 8192
rect 5610 7104 5931 8128
rect 5610 7040 5618 7104
rect 5682 7040 5698 7104
rect 5762 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5931 7104
rect 5610 6016 5931 7040
rect 5610 5952 5618 6016
rect 5682 5952 5698 6016
rect 5762 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5931 6016
rect 5610 4928 5931 5952
rect 5610 4864 5618 4928
rect 5682 4864 5698 4928
rect 5762 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5931 4928
rect 5610 3840 5931 4864
rect 5610 3776 5618 3840
rect 5682 3776 5698 3840
rect 5762 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5931 3840
rect 5610 2752 5931 3776
rect 5610 2688 5618 2752
rect 5682 2688 5698 2752
rect 5762 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5931 2752
rect 5610 2128 5931 2688
rect 7944 106656 8264 106672
rect 7944 106592 7952 106656
rect 8016 106592 8032 106656
rect 8096 106592 8112 106656
rect 8176 106592 8192 106656
rect 8256 106592 8264 106656
rect 7944 105568 8264 106592
rect 7944 105504 7952 105568
rect 8016 105504 8032 105568
rect 8096 105504 8112 105568
rect 8176 105504 8192 105568
rect 8256 105504 8264 105568
rect 7944 104480 8264 105504
rect 7944 104416 7952 104480
rect 8016 104416 8032 104480
rect 8096 104416 8112 104480
rect 8176 104416 8192 104480
rect 8256 104416 8264 104480
rect 7944 103392 8264 104416
rect 7944 103328 7952 103392
rect 8016 103328 8032 103392
rect 8096 103328 8112 103392
rect 8176 103328 8192 103392
rect 8256 103328 8264 103392
rect 7944 102304 8264 103328
rect 7944 102240 7952 102304
rect 8016 102240 8032 102304
rect 8096 102240 8112 102304
rect 8176 102240 8192 102304
rect 8256 102240 8264 102304
rect 7944 101216 8264 102240
rect 7944 101152 7952 101216
rect 8016 101152 8032 101216
rect 8096 101152 8112 101216
rect 8176 101152 8192 101216
rect 8256 101152 8264 101216
rect 7944 100128 8264 101152
rect 7944 100064 7952 100128
rect 8016 100064 8032 100128
rect 8096 100064 8112 100128
rect 8176 100064 8192 100128
rect 8256 100064 8264 100128
rect 7944 99040 8264 100064
rect 7944 98976 7952 99040
rect 8016 98976 8032 99040
rect 8096 98976 8112 99040
rect 8176 98976 8192 99040
rect 8256 98976 8264 99040
rect 7944 97952 8264 98976
rect 7944 97888 7952 97952
rect 8016 97888 8032 97952
rect 8096 97888 8112 97952
rect 8176 97888 8192 97952
rect 8256 97888 8264 97952
rect 7944 96864 8264 97888
rect 7944 96800 7952 96864
rect 8016 96800 8032 96864
rect 8096 96800 8112 96864
rect 8176 96800 8192 96864
rect 8256 96800 8264 96864
rect 7944 95776 8264 96800
rect 7944 95712 7952 95776
rect 8016 95712 8032 95776
rect 8096 95712 8112 95776
rect 8176 95712 8192 95776
rect 8256 95712 8264 95776
rect 7944 94688 8264 95712
rect 7944 94624 7952 94688
rect 8016 94624 8032 94688
rect 8096 94624 8112 94688
rect 8176 94624 8192 94688
rect 8256 94624 8264 94688
rect 7944 93600 8264 94624
rect 7944 93536 7952 93600
rect 8016 93536 8032 93600
rect 8096 93536 8112 93600
rect 8176 93536 8192 93600
rect 8256 93536 8264 93600
rect 7944 92512 8264 93536
rect 7944 92448 7952 92512
rect 8016 92448 8032 92512
rect 8096 92448 8112 92512
rect 8176 92448 8192 92512
rect 8256 92448 8264 92512
rect 7944 91424 8264 92448
rect 7944 91360 7952 91424
rect 8016 91360 8032 91424
rect 8096 91360 8112 91424
rect 8176 91360 8192 91424
rect 8256 91360 8264 91424
rect 7944 90336 8264 91360
rect 7944 90272 7952 90336
rect 8016 90272 8032 90336
rect 8096 90272 8112 90336
rect 8176 90272 8192 90336
rect 8256 90272 8264 90336
rect 7944 89248 8264 90272
rect 7944 89184 7952 89248
rect 8016 89184 8032 89248
rect 8096 89184 8112 89248
rect 8176 89184 8192 89248
rect 8256 89184 8264 89248
rect 7944 88160 8264 89184
rect 7944 88096 7952 88160
rect 8016 88096 8032 88160
rect 8096 88096 8112 88160
rect 8176 88096 8192 88160
rect 8256 88096 8264 88160
rect 7944 87072 8264 88096
rect 7944 87008 7952 87072
rect 8016 87008 8032 87072
rect 8096 87008 8112 87072
rect 8176 87008 8192 87072
rect 8256 87008 8264 87072
rect 7944 85984 8264 87008
rect 7944 85920 7952 85984
rect 8016 85920 8032 85984
rect 8096 85920 8112 85984
rect 8176 85920 8192 85984
rect 8256 85920 8264 85984
rect 7944 84896 8264 85920
rect 7944 84832 7952 84896
rect 8016 84832 8032 84896
rect 8096 84832 8112 84896
rect 8176 84832 8192 84896
rect 8256 84832 8264 84896
rect 7944 83808 8264 84832
rect 7944 83744 7952 83808
rect 8016 83744 8032 83808
rect 8096 83744 8112 83808
rect 8176 83744 8192 83808
rect 8256 83744 8264 83808
rect 7944 82720 8264 83744
rect 7944 82656 7952 82720
rect 8016 82656 8032 82720
rect 8096 82656 8112 82720
rect 8176 82656 8192 82720
rect 8256 82656 8264 82720
rect 7944 81632 8264 82656
rect 7944 81568 7952 81632
rect 8016 81568 8032 81632
rect 8096 81568 8112 81632
rect 8176 81568 8192 81632
rect 8256 81568 8264 81632
rect 7944 80544 8264 81568
rect 7944 80480 7952 80544
rect 8016 80480 8032 80544
rect 8096 80480 8112 80544
rect 8176 80480 8192 80544
rect 8256 80480 8264 80544
rect 7944 79456 8264 80480
rect 7944 79392 7952 79456
rect 8016 79392 8032 79456
rect 8096 79392 8112 79456
rect 8176 79392 8192 79456
rect 8256 79392 8264 79456
rect 7944 78368 8264 79392
rect 7944 78304 7952 78368
rect 8016 78304 8032 78368
rect 8096 78304 8112 78368
rect 8176 78304 8192 78368
rect 8256 78304 8264 78368
rect 7944 77280 8264 78304
rect 7944 77216 7952 77280
rect 8016 77216 8032 77280
rect 8096 77216 8112 77280
rect 8176 77216 8192 77280
rect 8256 77216 8264 77280
rect 7944 76192 8264 77216
rect 7944 76128 7952 76192
rect 8016 76128 8032 76192
rect 8096 76128 8112 76192
rect 8176 76128 8192 76192
rect 8256 76128 8264 76192
rect 7944 75104 8264 76128
rect 7944 75040 7952 75104
rect 8016 75040 8032 75104
rect 8096 75040 8112 75104
rect 8176 75040 8192 75104
rect 8256 75040 8264 75104
rect 7944 74016 8264 75040
rect 7944 73952 7952 74016
rect 8016 73952 8032 74016
rect 8096 73952 8112 74016
rect 8176 73952 8192 74016
rect 8256 73952 8264 74016
rect 7944 72928 8264 73952
rect 7944 72864 7952 72928
rect 8016 72864 8032 72928
rect 8096 72864 8112 72928
rect 8176 72864 8192 72928
rect 8256 72864 8264 72928
rect 7944 71840 8264 72864
rect 7944 71776 7952 71840
rect 8016 71776 8032 71840
rect 8096 71776 8112 71840
rect 8176 71776 8192 71840
rect 8256 71776 8264 71840
rect 7944 70752 8264 71776
rect 7944 70688 7952 70752
rect 8016 70688 8032 70752
rect 8096 70688 8112 70752
rect 8176 70688 8192 70752
rect 8256 70688 8264 70752
rect 7944 69664 8264 70688
rect 7944 69600 7952 69664
rect 8016 69600 8032 69664
rect 8096 69600 8112 69664
rect 8176 69600 8192 69664
rect 8256 69600 8264 69664
rect 7944 68576 8264 69600
rect 7944 68512 7952 68576
rect 8016 68512 8032 68576
rect 8096 68512 8112 68576
rect 8176 68512 8192 68576
rect 8256 68512 8264 68576
rect 7944 67488 8264 68512
rect 7944 67424 7952 67488
rect 8016 67424 8032 67488
rect 8096 67424 8112 67488
rect 8176 67424 8192 67488
rect 8256 67424 8264 67488
rect 7944 66400 8264 67424
rect 7944 66336 7952 66400
rect 8016 66336 8032 66400
rect 8096 66336 8112 66400
rect 8176 66336 8192 66400
rect 8256 66336 8264 66400
rect 7944 65312 8264 66336
rect 7944 65248 7952 65312
rect 8016 65248 8032 65312
rect 8096 65248 8112 65312
rect 8176 65248 8192 65312
rect 8256 65248 8264 65312
rect 7944 64224 8264 65248
rect 7944 64160 7952 64224
rect 8016 64160 8032 64224
rect 8096 64160 8112 64224
rect 8176 64160 8192 64224
rect 8256 64160 8264 64224
rect 7944 63136 8264 64160
rect 7944 63072 7952 63136
rect 8016 63072 8032 63136
rect 8096 63072 8112 63136
rect 8176 63072 8192 63136
rect 8256 63072 8264 63136
rect 7944 62048 8264 63072
rect 7944 61984 7952 62048
rect 8016 61984 8032 62048
rect 8096 61984 8112 62048
rect 8176 61984 8192 62048
rect 8256 61984 8264 62048
rect 7944 60960 8264 61984
rect 7944 60896 7952 60960
rect 8016 60896 8032 60960
rect 8096 60896 8112 60960
rect 8176 60896 8192 60960
rect 8256 60896 8264 60960
rect 7944 59872 8264 60896
rect 7944 59808 7952 59872
rect 8016 59808 8032 59872
rect 8096 59808 8112 59872
rect 8176 59808 8192 59872
rect 8256 59808 8264 59872
rect 7944 58784 8264 59808
rect 7944 58720 7952 58784
rect 8016 58720 8032 58784
rect 8096 58720 8112 58784
rect 8176 58720 8192 58784
rect 8256 58720 8264 58784
rect 7944 57696 8264 58720
rect 7944 57632 7952 57696
rect 8016 57632 8032 57696
rect 8096 57632 8112 57696
rect 8176 57632 8192 57696
rect 8256 57632 8264 57696
rect 7944 56608 8264 57632
rect 7944 56544 7952 56608
rect 8016 56544 8032 56608
rect 8096 56544 8112 56608
rect 8176 56544 8192 56608
rect 8256 56544 8264 56608
rect 7944 55520 8264 56544
rect 7944 55456 7952 55520
rect 8016 55456 8032 55520
rect 8096 55456 8112 55520
rect 8176 55456 8192 55520
rect 8256 55456 8264 55520
rect 7944 54432 8264 55456
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 10277 106112 10597 106672
rect 10277 106048 10285 106112
rect 10349 106048 10365 106112
rect 10429 106048 10445 106112
rect 10509 106048 10525 106112
rect 10589 106048 10597 106112
rect 10277 105024 10597 106048
rect 10277 104960 10285 105024
rect 10349 104960 10365 105024
rect 10429 104960 10445 105024
rect 10509 104960 10525 105024
rect 10589 104960 10597 105024
rect 10277 103936 10597 104960
rect 10277 103872 10285 103936
rect 10349 103872 10365 103936
rect 10429 103872 10445 103936
rect 10509 103872 10525 103936
rect 10589 103872 10597 103936
rect 10277 102848 10597 103872
rect 10277 102784 10285 102848
rect 10349 102784 10365 102848
rect 10429 102784 10445 102848
rect 10509 102784 10525 102848
rect 10589 102784 10597 102848
rect 10277 101760 10597 102784
rect 10277 101696 10285 101760
rect 10349 101696 10365 101760
rect 10429 101696 10445 101760
rect 10509 101696 10525 101760
rect 10589 101696 10597 101760
rect 10277 100672 10597 101696
rect 10277 100608 10285 100672
rect 10349 100608 10365 100672
rect 10429 100608 10445 100672
rect 10509 100608 10525 100672
rect 10589 100608 10597 100672
rect 10277 99584 10597 100608
rect 10277 99520 10285 99584
rect 10349 99520 10365 99584
rect 10429 99520 10445 99584
rect 10509 99520 10525 99584
rect 10589 99520 10597 99584
rect 10277 98496 10597 99520
rect 10277 98432 10285 98496
rect 10349 98432 10365 98496
rect 10429 98432 10445 98496
rect 10509 98432 10525 98496
rect 10589 98432 10597 98496
rect 10277 97408 10597 98432
rect 10277 97344 10285 97408
rect 10349 97344 10365 97408
rect 10429 97344 10445 97408
rect 10509 97344 10525 97408
rect 10589 97344 10597 97408
rect 10277 96320 10597 97344
rect 10277 96256 10285 96320
rect 10349 96256 10365 96320
rect 10429 96256 10445 96320
rect 10509 96256 10525 96320
rect 10589 96256 10597 96320
rect 10277 95232 10597 96256
rect 10277 95168 10285 95232
rect 10349 95168 10365 95232
rect 10429 95168 10445 95232
rect 10509 95168 10525 95232
rect 10589 95168 10597 95232
rect 10277 94144 10597 95168
rect 10277 94080 10285 94144
rect 10349 94080 10365 94144
rect 10429 94080 10445 94144
rect 10509 94080 10525 94144
rect 10589 94080 10597 94144
rect 10277 93056 10597 94080
rect 10277 92992 10285 93056
rect 10349 92992 10365 93056
rect 10429 92992 10445 93056
rect 10509 92992 10525 93056
rect 10589 92992 10597 93056
rect 10277 91968 10597 92992
rect 10277 91904 10285 91968
rect 10349 91904 10365 91968
rect 10429 91904 10445 91968
rect 10509 91904 10525 91968
rect 10589 91904 10597 91968
rect 10277 90880 10597 91904
rect 10277 90816 10285 90880
rect 10349 90816 10365 90880
rect 10429 90816 10445 90880
rect 10509 90816 10525 90880
rect 10589 90816 10597 90880
rect 10277 89792 10597 90816
rect 10277 89728 10285 89792
rect 10349 89728 10365 89792
rect 10429 89728 10445 89792
rect 10509 89728 10525 89792
rect 10589 89728 10597 89792
rect 10277 88704 10597 89728
rect 10277 88640 10285 88704
rect 10349 88640 10365 88704
rect 10429 88640 10445 88704
rect 10509 88640 10525 88704
rect 10589 88640 10597 88704
rect 10277 87616 10597 88640
rect 10277 87552 10285 87616
rect 10349 87552 10365 87616
rect 10429 87552 10445 87616
rect 10509 87552 10525 87616
rect 10589 87552 10597 87616
rect 10277 86528 10597 87552
rect 10277 86464 10285 86528
rect 10349 86464 10365 86528
rect 10429 86464 10445 86528
rect 10509 86464 10525 86528
rect 10589 86464 10597 86528
rect 10277 85440 10597 86464
rect 10277 85376 10285 85440
rect 10349 85376 10365 85440
rect 10429 85376 10445 85440
rect 10509 85376 10525 85440
rect 10589 85376 10597 85440
rect 10277 84352 10597 85376
rect 10277 84288 10285 84352
rect 10349 84288 10365 84352
rect 10429 84288 10445 84352
rect 10509 84288 10525 84352
rect 10589 84288 10597 84352
rect 10277 83264 10597 84288
rect 10277 83200 10285 83264
rect 10349 83200 10365 83264
rect 10429 83200 10445 83264
rect 10509 83200 10525 83264
rect 10589 83200 10597 83264
rect 10277 82176 10597 83200
rect 10277 82112 10285 82176
rect 10349 82112 10365 82176
rect 10429 82112 10445 82176
rect 10509 82112 10525 82176
rect 10589 82112 10597 82176
rect 10277 81088 10597 82112
rect 10277 81024 10285 81088
rect 10349 81024 10365 81088
rect 10429 81024 10445 81088
rect 10509 81024 10525 81088
rect 10589 81024 10597 81088
rect 10277 80000 10597 81024
rect 10277 79936 10285 80000
rect 10349 79936 10365 80000
rect 10429 79936 10445 80000
rect 10509 79936 10525 80000
rect 10589 79936 10597 80000
rect 10277 78912 10597 79936
rect 10277 78848 10285 78912
rect 10349 78848 10365 78912
rect 10429 78848 10445 78912
rect 10509 78848 10525 78912
rect 10589 78848 10597 78912
rect 10277 77824 10597 78848
rect 10277 77760 10285 77824
rect 10349 77760 10365 77824
rect 10429 77760 10445 77824
rect 10509 77760 10525 77824
rect 10589 77760 10597 77824
rect 10277 76736 10597 77760
rect 10277 76672 10285 76736
rect 10349 76672 10365 76736
rect 10429 76672 10445 76736
rect 10509 76672 10525 76736
rect 10589 76672 10597 76736
rect 10277 75648 10597 76672
rect 10277 75584 10285 75648
rect 10349 75584 10365 75648
rect 10429 75584 10445 75648
rect 10509 75584 10525 75648
rect 10589 75584 10597 75648
rect 10277 74560 10597 75584
rect 10277 74496 10285 74560
rect 10349 74496 10365 74560
rect 10429 74496 10445 74560
rect 10509 74496 10525 74560
rect 10589 74496 10597 74560
rect 10277 73472 10597 74496
rect 10277 73408 10285 73472
rect 10349 73408 10365 73472
rect 10429 73408 10445 73472
rect 10509 73408 10525 73472
rect 10589 73408 10597 73472
rect 10277 72384 10597 73408
rect 10277 72320 10285 72384
rect 10349 72320 10365 72384
rect 10429 72320 10445 72384
rect 10509 72320 10525 72384
rect 10589 72320 10597 72384
rect 10277 71296 10597 72320
rect 10277 71232 10285 71296
rect 10349 71232 10365 71296
rect 10429 71232 10445 71296
rect 10509 71232 10525 71296
rect 10589 71232 10597 71296
rect 10277 70208 10597 71232
rect 10277 70144 10285 70208
rect 10349 70144 10365 70208
rect 10429 70144 10445 70208
rect 10509 70144 10525 70208
rect 10589 70144 10597 70208
rect 10277 69120 10597 70144
rect 10277 69056 10285 69120
rect 10349 69056 10365 69120
rect 10429 69056 10445 69120
rect 10509 69056 10525 69120
rect 10589 69056 10597 69120
rect 10277 68032 10597 69056
rect 10277 67968 10285 68032
rect 10349 67968 10365 68032
rect 10429 67968 10445 68032
rect 10509 67968 10525 68032
rect 10589 67968 10597 68032
rect 10277 66944 10597 67968
rect 10277 66880 10285 66944
rect 10349 66880 10365 66944
rect 10429 66880 10445 66944
rect 10509 66880 10525 66944
rect 10589 66880 10597 66944
rect 10277 65856 10597 66880
rect 10277 65792 10285 65856
rect 10349 65792 10365 65856
rect 10429 65792 10445 65856
rect 10509 65792 10525 65856
rect 10589 65792 10597 65856
rect 10277 64768 10597 65792
rect 10277 64704 10285 64768
rect 10349 64704 10365 64768
rect 10429 64704 10445 64768
rect 10509 64704 10525 64768
rect 10589 64704 10597 64768
rect 10277 63680 10597 64704
rect 10277 63616 10285 63680
rect 10349 63616 10365 63680
rect 10429 63616 10445 63680
rect 10509 63616 10525 63680
rect 10589 63616 10597 63680
rect 10277 62592 10597 63616
rect 10277 62528 10285 62592
rect 10349 62528 10365 62592
rect 10429 62528 10445 62592
rect 10509 62528 10525 62592
rect 10589 62528 10597 62592
rect 10277 61504 10597 62528
rect 10277 61440 10285 61504
rect 10349 61440 10365 61504
rect 10429 61440 10445 61504
rect 10509 61440 10525 61504
rect 10589 61440 10597 61504
rect 10277 60416 10597 61440
rect 10277 60352 10285 60416
rect 10349 60352 10365 60416
rect 10429 60352 10445 60416
rect 10509 60352 10525 60416
rect 10589 60352 10597 60416
rect 10277 59328 10597 60352
rect 10277 59264 10285 59328
rect 10349 59264 10365 59328
rect 10429 59264 10445 59328
rect 10509 59264 10525 59328
rect 10589 59264 10597 59328
rect 10277 58240 10597 59264
rect 10277 58176 10285 58240
rect 10349 58176 10365 58240
rect 10429 58176 10445 58240
rect 10509 58176 10525 58240
rect 10589 58176 10597 58240
rect 10277 57152 10597 58176
rect 10277 57088 10285 57152
rect 10349 57088 10365 57152
rect 10429 57088 10445 57152
rect 10509 57088 10525 57152
rect 10589 57088 10597 57152
rect 10277 56064 10597 57088
rect 10277 56000 10285 56064
rect 10349 56000 10365 56064
rect 10429 56000 10445 56064
rect 10509 56000 10525 56064
rect 10589 56000 10597 56064
rect 10277 54976 10597 56000
rect 10277 54912 10285 54976
rect 10349 54912 10365 54976
rect 10429 54912 10445 54976
rect 10509 54912 10525 54976
rect 10589 54912 10597 54976
rect 10277 53888 10597 54912
rect 10277 53824 10285 53888
rect 10349 53824 10365 53888
rect 10429 53824 10445 53888
rect 10509 53824 10525 53888
rect 10589 53824 10597 53888
rect 10277 52800 10597 53824
rect 10277 52736 10285 52800
rect 10349 52736 10365 52800
rect 10429 52736 10445 52800
rect 10509 52736 10525 52800
rect 10589 52736 10597 52800
rect 10277 51712 10597 52736
rect 10277 51648 10285 51712
rect 10349 51648 10365 51712
rect 10429 51648 10445 51712
rect 10509 51648 10525 51712
rect 10589 51648 10597 51712
rect 10277 50624 10597 51648
rect 10277 50560 10285 50624
rect 10349 50560 10365 50624
rect 10429 50560 10445 50624
rect 10509 50560 10525 50624
rect 10589 50560 10597 50624
rect 10277 49536 10597 50560
rect 10277 49472 10285 49536
rect 10349 49472 10365 49536
rect 10429 49472 10445 49536
rect 10509 49472 10525 49536
rect 10589 49472 10597 49536
rect 10277 48448 10597 49472
rect 10277 48384 10285 48448
rect 10349 48384 10365 48448
rect 10429 48384 10445 48448
rect 10509 48384 10525 48448
rect 10589 48384 10597 48448
rect 10277 47360 10597 48384
rect 10277 47296 10285 47360
rect 10349 47296 10365 47360
rect 10429 47296 10445 47360
rect 10509 47296 10525 47360
rect 10589 47296 10597 47360
rect 10277 46272 10597 47296
rect 10277 46208 10285 46272
rect 10349 46208 10365 46272
rect 10429 46208 10445 46272
rect 10509 46208 10525 46272
rect 10589 46208 10597 46272
rect 10277 45184 10597 46208
rect 10277 45120 10285 45184
rect 10349 45120 10365 45184
rect 10429 45120 10445 45184
rect 10509 45120 10525 45184
rect 10589 45120 10597 45184
rect 10277 44096 10597 45120
rect 10277 44032 10285 44096
rect 10349 44032 10365 44096
rect 10429 44032 10445 44096
rect 10509 44032 10525 44096
rect 10589 44032 10597 44096
rect 10277 43008 10597 44032
rect 10277 42944 10285 43008
rect 10349 42944 10365 43008
rect 10429 42944 10445 43008
rect 10509 42944 10525 43008
rect 10589 42944 10597 43008
rect 10277 41920 10597 42944
rect 10277 41856 10285 41920
rect 10349 41856 10365 41920
rect 10429 41856 10445 41920
rect 10509 41856 10525 41920
rect 10589 41856 10597 41920
rect 10277 40832 10597 41856
rect 10277 40768 10285 40832
rect 10349 40768 10365 40832
rect 10429 40768 10445 40832
rect 10509 40768 10525 40832
rect 10589 40768 10597 40832
rect 10277 39744 10597 40768
rect 10277 39680 10285 39744
rect 10349 39680 10365 39744
rect 10429 39680 10445 39744
rect 10509 39680 10525 39744
rect 10589 39680 10597 39744
rect 10277 38656 10597 39680
rect 10277 38592 10285 38656
rect 10349 38592 10365 38656
rect 10429 38592 10445 38656
rect 10509 38592 10525 38656
rect 10589 38592 10597 38656
rect 10277 37568 10597 38592
rect 10277 37504 10285 37568
rect 10349 37504 10365 37568
rect 10429 37504 10445 37568
rect 10509 37504 10525 37568
rect 10589 37504 10597 37568
rect 10277 36480 10597 37504
rect 10277 36416 10285 36480
rect 10349 36416 10365 36480
rect 10429 36416 10445 36480
rect 10509 36416 10525 36480
rect 10589 36416 10597 36480
rect 10277 35392 10597 36416
rect 10277 35328 10285 35392
rect 10349 35328 10365 35392
rect 10429 35328 10445 35392
rect 10509 35328 10525 35392
rect 10589 35328 10597 35392
rect 10277 34304 10597 35328
rect 10277 34240 10285 34304
rect 10349 34240 10365 34304
rect 10429 34240 10445 34304
rect 10509 34240 10525 34304
rect 10589 34240 10597 34304
rect 10277 33216 10597 34240
rect 10277 33152 10285 33216
rect 10349 33152 10365 33216
rect 10429 33152 10445 33216
rect 10509 33152 10525 33216
rect 10589 33152 10597 33216
rect 10277 32128 10597 33152
rect 10277 32064 10285 32128
rect 10349 32064 10365 32128
rect 10429 32064 10445 32128
rect 10509 32064 10525 32128
rect 10589 32064 10597 32128
rect 10277 31040 10597 32064
rect 10277 30976 10285 31040
rect 10349 30976 10365 31040
rect 10429 30976 10445 31040
rect 10509 30976 10525 31040
rect 10589 30976 10597 31040
rect 10277 29952 10597 30976
rect 10277 29888 10285 29952
rect 10349 29888 10365 29952
rect 10429 29888 10445 29952
rect 10509 29888 10525 29952
rect 10589 29888 10597 29952
rect 10277 28864 10597 29888
rect 10277 28800 10285 28864
rect 10349 28800 10365 28864
rect 10429 28800 10445 28864
rect 10509 28800 10525 28864
rect 10589 28800 10597 28864
rect 10277 27776 10597 28800
rect 10277 27712 10285 27776
rect 10349 27712 10365 27776
rect 10429 27712 10445 27776
rect 10509 27712 10525 27776
rect 10589 27712 10597 27776
rect 10277 26688 10597 27712
rect 10277 26624 10285 26688
rect 10349 26624 10365 26688
rect 10429 26624 10445 26688
rect 10509 26624 10525 26688
rect 10589 26624 10597 26688
rect 10277 25600 10597 26624
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_384 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_nor4_4  _15_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__15__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__D
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__B
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_74 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_91
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_104
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 12880 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 12880 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__15__C
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_109
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 12880 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_1  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _19_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 12880 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 12880 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 12880 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 12880 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 12880 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 12880 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 12880 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 12880 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 12880 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 12880 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 12880 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 12880 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_102
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_106
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 12880 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__14__C
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_85
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_99
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_111
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_123
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 12880 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_nor4_4  _14_
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__14__D
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__B
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 12880 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 12880 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _11_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 12880 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 12880 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_111
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 12880 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 590 592
use scs8hd_inv_8  _06_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _08_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__05__B
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_124
timestamp 1586364061
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 12880 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_69
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use scs8hd_and4_4  _07_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_and4_4  _09_
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__C
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_94
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_115
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 12880 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 590 592
use scs8hd_and4_4  _10_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_and4_4  _05_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__D
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_118
timestamp 1586364061
transform 1 0 11960 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_124
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 12880 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_106
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 12880 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_78
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_nor4_4  _13_
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_103
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 314 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_115
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 12880 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 12880 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_109
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 12880 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 12880 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_82
timestamp 1586364061
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_90
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_99
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_115
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_123
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 12880 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 12880 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 12880 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 12880 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 12880 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 12880 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 12880 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 12880 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 12880 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 12880 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 12880 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 12880 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_117
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 12880 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 12880 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_44
timestamp 1586364061
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_56
timestamp 1586364061
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_108
timestamp 1586364061
transform 1 0 11040 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_120
timestamp 1586364061
transform 1 0 12144 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_124
timestamp 1586364061
transform 1 0 12512 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 12880 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 10672 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_45_114
timestamp 1586364061
transform 1 0 11592 0 1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 12880 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_12  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 12880 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 12880 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_105
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_117
timestamp 1586364061
transform 1 0 11868 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 12880 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_110
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 12880 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 12880 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_98
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 12880 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_105
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_117
timestamp 1586364061
transform 1 0 11868 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_114
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_118
timestamp 1586364061
transform 1 0 11960 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 12880 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 12880 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_105
timestamp 1586364061
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 12880 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_98
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_110
timestamp 1586364061
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 12880 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 12880 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_110
timestamp 1586364061
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 12880 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 12880 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_98
timestamp 1586364061
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_110
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 12880 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 12880 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 12880 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 12880 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 12880 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_68
timestamp 1586364061
transform 1 0 7360 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_80
timestamp 1586364061
transform 1 0 8464 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_93
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_105
timestamp 1586364061
transform 1 0 10764 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_117
timestamp 1586364061
transform 1 0 11868 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 12880 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_3  PHY_130
timestamp 1586364061
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_65_3
timestamp 1586364061
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_15
timestamp 1586364061
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_27
timestamp 1586364061
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_39
timestamp 1586364061
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_65_51
timestamp 1586364061
transform 1 0 5796 0 1 37536
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_59
timestamp 1586364061
transform 1 0 6532 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_62
timestamp 1586364061
transform 1 0 6808 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_74
timestamp 1586364061
transform 1 0 7912 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_86
timestamp 1586364061
transform 1 0 9016 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_98
timestamp 1586364061
transform 1 0 10120 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_110
timestamp 1586364061
transform 1 0 11224 0 1 37536
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_65_123
timestamp 1586364061
transform 1 0 12420 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  PHY_131
timestamp 1586364061
transform -1 0 12880 0 1 37536
box -38 -48 314 592
use scs8hd_decap_3  PHY_132
timestamp 1586364061
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_134
timestamp 1586364061
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_66_3
timestamp 1586364061
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_15
timestamp 1586364061
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_3
timestamp 1586364061
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_15
timestamp 1586364061
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_27
timestamp 1586364061
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_66_32
timestamp 1586364061
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_27
timestamp 1586364061
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_44
timestamp 1586364061
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_39
timestamp 1586364061
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_67_51
timestamp 1586364061
transform 1 0 5796 0 1 38624
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_56
timestamp 1586364061
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_68
timestamp 1586364061
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_67_59
timestamp 1586364061
transform 1 0 6532 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_67_62
timestamp 1586364061
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_80
timestamp 1586364061
transform 1 0 8464 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_74
timestamp 1586364061
transform 1 0 7912 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_86
timestamp 1586364061
transform 1 0 9016 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_93
timestamp 1586364061
transform 1 0 9660 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_105
timestamp 1586364061
transform 1 0 10764 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_98
timestamp 1586364061
transform 1 0 10120 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use scs8hd_decap_8  FILLER_66_117
timestamp 1586364061
transform 1 0 11868 0 -1 38624
box -38 -48 774 592
use scs8hd_decap_12  FILLER_67_110
timestamp 1586364061
transform 1 0 11224 0 1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_67_123
timestamp 1586364061
transform 1 0 12420 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  PHY_133
timestamp 1586364061
transform -1 0 12880 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_135
timestamp 1586364061
transform -1 0 12880 0 1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_136
timestamp 1586364061
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_68_3
timestamp 1586364061
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_15
timestamp 1586364061
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_27
timestamp 1586364061
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_68_32
timestamp 1586364061
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_44
timestamp 1586364061
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_56
timestamp 1586364061
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_68
timestamp 1586364061
transform 1 0 7360 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_80
timestamp 1586364061
transform 1 0 8464 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_68_93
timestamp 1586364061
transform 1 0 9660 0 -1 39712
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_68_105
timestamp 1586364061
transform 1 0 10764 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_108
timestamp 1586364061
transform 1 0 11040 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_68_120
timestamp 1586364061
transform 1 0 12144 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_68_124
timestamp 1586364061
transform 1 0 12512 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  PHY_137
timestamp 1586364061
transform -1 0 12880 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_3  PHY_138
timestamp 1586364061
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_3
timestamp 1586364061
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_15
timestamp 1586364061
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_27
timestamp 1586364061
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_39
timestamp 1586364061
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_51
timestamp 1586364061
transform 1 0 5796 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_59
timestamp 1586364061
transform 1 0 6532 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_62
timestamp 1586364061
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_74
timestamp 1586364061
transform 1 0 7912 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_86
timestamp 1586364061
transform 1 0 9016 0 1 39712
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 10856 0 1 39712
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 10672 0 1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_69_98
timestamp 1586364061
transform 1 0 10120 0 1 39712
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use scs8hd_decap_8  FILLER_69_114
timestamp 1586364061
transform 1 0 11592 0 1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_69_123
timestamp 1586364061
transform 1 0 12420 0 1 39712
box -38 -48 222 592
use scs8hd_decap_3  PHY_139
timestamp 1586364061
transform -1 0 12880 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  PHY_140
timestamp 1586364061
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_70_3
timestamp 1586364061
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_15
timestamp 1586364061
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_27
timestamp 1586364061
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_70_32
timestamp 1586364061
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_44
timestamp 1586364061
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_56
timestamp 1586364061
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_68
timestamp 1586364061
transform 1 0 7360 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_80
timestamp 1586364061
transform 1 0 8464 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_93
timestamp 1586364061
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_105
timestamp 1586364061
transform 1 0 10764 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_70_117
timestamp 1586364061
transform 1 0 11868 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_3  PHY_141
timestamp 1586364061
transform -1 0 12880 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_3  PHY_142
timestamp 1586364061
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_3
timestamp 1586364061
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_15
timestamp 1586364061
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_27
timestamp 1586364061
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_39
timestamp 1586364061
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_71_51
timestamp 1586364061
transform 1 0 5796 0 1 40800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_59
timestamp 1586364061
transform 1 0 6532 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_62
timestamp 1586364061
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_74
timestamp 1586364061
transform 1 0 7912 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_86
timestamp 1586364061
transform 1 0 9016 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_98
timestamp 1586364061
transform 1 0 10120 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_110
timestamp 1586364061
transform 1 0 11224 0 1 40800
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_71_123
timestamp 1586364061
transform 1 0 12420 0 1 40800
box -38 -48 222 592
use scs8hd_decap_3  PHY_143
timestamp 1586364061
transform -1 0 12880 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  PHY_144
timestamp 1586364061
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_146
timestamp 1586364061
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_72_3
timestamp 1586364061
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_15
timestamp 1586364061
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_3
timestamp 1586364061
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_15
timestamp 1586364061
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_27
timestamp 1586364061
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_72_32
timestamp 1586364061
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_27
timestamp 1586364061
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_44
timestamp 1586364061
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_39
timestamp 1586364061
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_51
timestamp 1586364061
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_56
timestamp 1586364061
transform 1 0 6256 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_68
timestamp 1586364061
transform 1 0 7360 0 -1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_73_59
timestamp 1586364061
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_73_62
timestamp 1586364061
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_80
timestamp 1586364061
transform 1 0 8464 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_74
timestamp 1586364061
transform 1 0 7912 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_86
timestamp 1586364061
transform 1 0 9016 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_93
timestamp 1586364061
transform 1 0 9660 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_105
timestamp 1586364061
transform 1 0 10764 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_98
timestamp 1586364061
transform 1 0 10120 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use scs8hd_decap_8  FILLER_72_117
timestamp 1586364061
transform 1 0 11868 0 -1 41888
box -38 -48 774 592
use scs8hd_decap_12  FILLER_73_110
timestamp 1586364061
transform 1 0 11224 0 1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_73_123
timestamp 1586364061
transform 1 0 12420 0 1 41888
box -38 -48 222 592
use scs8hd_decap_3  PHY_145
timestamp 1586364061
transform -1 0 12880 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_147
timestamp 1586364061
transform -1 0 12880 0 1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_148
timestamp 1586364061
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_74_3
timestamp 1586364061
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_15
timestamp 1586364061
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_27
timestamp 1586364061
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_74_32
timestamp 1586364061
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_44
timestamp 1586364061
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_56
timestamp 1586364061
transform 1 0 6256 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_68
timestamp 1586364061
transform 1 0 7360 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_80
timestamp 1586364061
transform 1 0 8464 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_93
timestamp 1586364061
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_105
timestamp 1586364061
transform 1 0 10764 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_74_117
timestamp 1586364061
transform 1 0 11868 0 -1 42976
box -38 -48 774 592
use scs8hd_decap_3  PHY_149
timestamp 1586364061
transform -1 0 12880 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_3  PHY_150
timestamp 1586364061
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_3
timestamp 1586364061
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_15
timestamp 1586364061
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_27
timestamp 1586364061
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_39
timestamp 1586364061
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_75_51
timestamp 1586364061
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_75_59
timestamp 1586364061
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_62
timestamp 1586364061
transform 1 0 6808 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_74
timestamp 1586364061
transform 1 0 7912 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_86
timestamp 1586364061
transform 1 0 9016 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_98
timestamp 1586364061
transform 1 0 10120 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_110
timestamp 1586364061
transform 1 0 11224 0 1 42976
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_75_123
timestamp 1586364061
transform 1 0 12420 0 1 42976
box -38 -48 222 592
use scs8hd_decap_3  PHY_151
timestamp 1586364061
transform -1 0 12880 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  PHY_152
timestamp 1586364061
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_3
timestamp 1586364061
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_15
timestamp 1586364061
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_76_27
timestamp 1586364061
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_76_32
timestamp 1586364061
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_44
timestamp 1586364061
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_56
timestamp 1586364061
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_68
timestamp 1586364061
transform 1 0 7360 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_80
timestamp 1586364061
transform 1 0 8464 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_93
timestamp 1586364061
transform 1 0 9660 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_105
timestamp 1586364061
transform 1 0 10764 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_76_117
timestamp 1586364061
transform 1 0 11868 0 -1 44064
box -38 -48 774 592
use scs8hd_decap_3  PHY_153
timestamp 1586364061
transform -1 0 12880 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_3  PHY_154
timestamp 1586364061
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_77_3
timestamp 1586364061
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_15
timestamp 1586364061
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_27
timestamp 1586364061
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_39
timestamp 1586364061
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_77_51
timestamp 1586364061
transform 1 0 5796 0 1 44064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_59
timestamp 1586364061
transform 1 0 6532 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_62
timestamp 1586364061
transform 1 0 6808 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_74
timestamp 1586364061
transform 1 0 7912 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_86
timestamp 1586364061
transform 1 0 9016 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_98
timestamp 1586364061
transform 1 0 10120 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 11500 0 1 44064
box -38 -48 222 592
use scs8hd_decap_3  FILLER_77_110
timestamp 1586364061
transform 1 0 11224 0 1 44064
box -38 -48 314 592
use scs8hd_decap_6  FILLER_77_115
timestamp 1586364061
transform 1 0 11684 0 1 44064
box -38 -48 590 592
use scs8hd_fill_1  FILLER_77_121
timestamp 1586364061
transform 1 0 12236 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_123
timestamp 1586364061
transform 1 0 12420 0 1 44064
box -38 -48 222 592
use scs8hd_decap_3  PHY_155
timestamp 1586364061
transform -1 0 12880 0 1 44064
box -38 -48 314 592
use scs8hd_decap_3  PHY_156
timestamp 1586364061
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_78_3
timestamp 1586364061
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_15
timestamp 1586364061
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_27
timestamp 1586364061
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_78_32
timestamp 1586364061
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_44
timestamp 1586364061
transform 1 0 5152 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_56
timestamp 1586364061
transform 1 0 6256 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_68
timestamp 1586364061
transform 1 0 7360 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_80
timestamp 1586364061
transform 1 0 8464 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_93
timestamp 1586364061
transform 1 0 9660 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_78_105
timestamp 1586364061
transform 1 0 10764 0 -1 45152
box -38 -48 774 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 11500 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_8  FILLER_78_117
timestamp 1586364061
transform 1 0 11868 0 -1 45152
box -38 -48 774 592
use scs8hd_decap_3  PHY_157
timestamp 1586364061
transform -1 0 12880 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_158
timestamp 1586364061
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_160
timestamp 1586364061
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_79_3
timestamp 1586364061
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_15
timestamp 1586364061
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_3
timestamp 1586364061
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_15
timestamp 1586364061
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_27
timestamp 1586364061
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_80_27
timestamp 1586364061
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_80_32
timestamp 1586364061
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_39
timestamp 1586364061
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_79_51
timestamp 1586364061
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use scs8hd_decap_12  FILLER_80_44
timestamp 1586364061
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_79_59
timestamp 1586364061
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_62
timestamp 1586364061
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_56
timestamp 1586364061
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_68
timestamp 1586364061
transform 1 0 7360 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_74
timestamp 1586364061
transform 1 0 7912 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_86
timestamp 1586364061
transform 1 0 9016 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_80
timestamp 1586364061
transform 1 0 8464 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_98
timestamp 1586364061
transform 1 0 10120 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_93
timestamp 1586364061
transform 1 0 9660 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_105
timestamp 1586364061
transform 1 0 10764 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_110
timestamp 1586364061
transform 1 0 11224 0 1 45152
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_79_123
timestamp 1586364061
transform 1 0 12420 0 1 45152
box -38 -48 222 592
use scs8hd_decap_8  FILLER_80_117
timestamp 1586364061
transform 1 0 11868 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_3  PHY_159
timestamp 1586364061
transform -1 0 12880 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_161
timestamp 1586364061
transform -1 0 12880 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_3  PHY_162
timestamp 1586364061
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_3
timestamp 1586364061
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_15
timestamp 1586364061
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_27
timestamp 1586364061
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_39
timestamp 1586364061
transform 1 0 4692 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_81_51
timestamp 1586364061
transform 1 0 5796 0 1 46240
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_81_59
timestamp 1586364061
transform 1 0 6532 0 1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_81_62
timestamp 1586364061
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_74
timestamp 1586364061
transform 1 0 7912 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_86
timestamp 1586364061
transform 1 0 9016 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_98
timestamp 1586364061
transform 1 0 10120 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_110
timestamp 1586364061
transform 1 0 11224 0 1 46240
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_81_123
timestamp 1586364061
transform 1 0 12420 0 1 46240
box -38 -48 222 592
use scs8hd_decap_3  PHY_163
timestamp 1586364061
transform -1 0 12880 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  PHY_164
timestamp 1586364061
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_3
timestamp 1586364061
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_15
timestamp 1586364061
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_4  FILLER_82_27
timestamp 1586364061
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_82_32
timestamp 1586364061
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_44
timestamp 1586364061
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_56
timestamp 1586364061
transform 1 0 6256 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_68
timestamp 1586364061
transform 1 0 7360 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_80
timestamp 1586364061
transform 1 0 8464 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 9568 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_93
timestamp 1586364061
transform 1 0 9660 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_105
timestamp 1586364061
transform 1 0 10764 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_82_117
timestamp 1586364061
transform 1 0 11868 0 -1 47328
box -38 -48 774 592
use scs8hd_decap_3  PHY_165
timestamp 1586364061
transform -1 0 12880 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_3  PHY_166
timestamp 1586364061
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_83_3
timestamp 1586364061
transform 1 0 1380 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_15
timestamp 1586364061
transform 1 0 2484 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_27
timestamp 1586364061
transform 1 0 3588 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_39
timestamp 1586364061
transform 1 0 4692 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_83_51
timestamp 1586364061
transform 1 0 5796 0 1 47328
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 6716 0 1 47328
box -38 -48 130 592
use scs8hd_fill_2  FILLER_83_59
timestamp 1586364061
transform 1 0 6532 0 1 47328
box -38 -48 222 592
use scs8hd_decap_12  FILLER_83_62
timestamp 1586364061
transform 1 0 6808 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_74
timestamp 1586364061
transform 1 0 7912 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_86
timestamp 1586364061
transform 1 0 9016 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_98
timestamp 1586364061
transform 1 0 10120 0 1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 12328 0 1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_83_110
timestamp 1586364061
transform 1 0 11224 0 1 47328
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_83_123
timestamp 1586364061
transform 1 0 12420 0 1 47328
box -38 -48 222 592
use scs8hd_decap_3  PHY_167
timestamp 1586364061
transform -1 0 12880 0 1 47328
box -38 -48 314 592
use scs8hd_decap_3  PHY_168
timestamp 1586364061
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use scs8hd_decap_12  FILLER_84_3
timestamp 1586364061
transform 1 0 1380 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_15
timestamp 1586364061
transform 1 0 2484 0 -1 48416
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 3956 0 -1 48416
box -38 -48 130 592
use scs8hd_decap_4  FILLER_84_27
timestamp 1586364061
transform 1 0 3588 0 -1 48416
box -38 -48 406 592
use scs8hd_decap_12  FILLER_84_32
timestamp 1586364061
transform 1 0 4048 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_44
timestamp 1586364061
transform 1 0 5152 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_56
timestamp 1586364061
transform 1 0 6256 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_68
timestamp 1586364061
transform 1 0 7360 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_80
timestamp 1586364061
transform 1 0 8464 0 -1 48416
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 9568 0 -1 48416
box -38 -48 130 592
use scs8hd_decap_12  FILLER_84_93
timestamp 1586364061
transform 1 0 9660 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_105
timestamp 1586364061
transform 1 0 10764 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_84_117
timestamp 1586364061
transform 1 0 11868 0 -1 48416
box -38 -48 774 592
use scs8hd_decap_3  PHY_169
timestamp 1586364061
transform -1 0 12880 0 -1 48416
box -38 -48 314 592
use scs8hd_decap_3  PHY_170
timestamp 1586364061
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use scs8hd_decap_3  PHY_172
timestamp 1586364061
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use scs8hd_decap_12  FILLER_85_3
timestamp 1586364061
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_85_15
timestamp 1586364061
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_3
timestamp 1586364061
transform 1 0 1380 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_15
timestamp 1586364061
transform 1 0 2484 0 -1 49504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 3956 0 -1 49504
box -38 -48 130 592
use scs8hd_decap_12  FILLER_85_27
timestamp 1586364061
transform 1 0 3588 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_86_27
timestamp 1586364061
transform 1 0 3588 0 -1 49504
box -38 -48 406 592
use scs8hd_decap_12  FILLER_86_32
timestamp 1586364061
transform 1 0 4048 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_85_39
timestamp 1586364061
transform 1 0 4692 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_85_51
timestamp 1586364061
transform 1 0 5796 0 1 48416
box -38 -48 774 592
use scs8hd_decap_12  FILLER_86_44
timestamp 1586364061
transform 1 0 5152 0 -1 49504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 6716 0 1 48416
box -38 -48 130 592
use scs8hd_fill_2  FILLER_85_59
timestamp 1586364061
transform 1 0 6532 0 1 48416
box -38 -48 222 592
use scs8hd_decap_12  FILLER_85_62
timestamp 1586364061
transform 1 0 6808 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_56
timestamp 1586364061
transform 1 0 6256 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_68
timestamp 1586364061
transform 1 0 7360 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_85_74
timestamp 1586364061
transform 1 0 7912 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_85_86
timestamp 1586364061
transform 1 0 9016 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_80
timestamp 1586364061
transform 1 0 8464 0 -1 49504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 9568 0 -1 49504
box -38 -48 130 592
use scs8hd_decap_12  FILLER_85_98
timestamp 1586364061
transform 1 0 10120 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_93
timestamp 1586364061
transform 1 0 9660 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_105
timestamp 1586364061
transform 1 0 10764 0 -1 49504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 12328 0 1 48416
box -38 -48 130 592
use scs8hd_decap_12  FILLER_85_110
timestamp 1586364061
transform 1 0 11224 0 1 48416
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_85_123
timestamp 1586364061
transform 1 0 12420 0 1 48416
box -38 -48 222 592
use scs8hd_decap_8  FILLER_86_117
timestamp 1586364061
transform 1 0 11868 0 -1 49504
box -38 -48 774 592
use scs8hd_decap_3  PHY_171
timestamp 1586364061
transform -1 0 12880 0 1 48416
box -38 -48 314 592
use scs8hd_decap_3  PHY_173
timestamp 1586364061
transform -1 0 12880 0 -1 49504
box -38 -48 314 592
use scs8hd_decap_3  PHY_174
timestamp 1586364061
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use scs8hd_decap_12  FILLER_87_3
timestamp 1586364061
transform 1 0 1380 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_15
timestamp 1586364061
transform 1 0 2484 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_27
timestamp 1586364061
transform 1 0 3588 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_39
timestamp 1586364061
transform 1 0 4692 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_87_51
timestamp 1586364061
transform 1 0 5796 0 1 49504
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 6716 0 1 49504
box -38 -48 130 592
use scs8hd_fill_2  FILLER_87_59
timestamp 1586364061
transform 1 0 6532 0 1 49504
box -38 -48 222 592
use scs8hd_decap_12  FILLER_87_62
timestamp 1586364061
transform 1 0 6808 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_74
timestamp 1586364061
transform 1 0 7912 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_86
timestamp 1586364061
transform 1 0 9016 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_98
timestamp 1586364061
transform 1 0 10120 0 1 49504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 12328 0 1 49504
box -38 -48 130 592
use scs8hd_decap_12  FILLER_87_110
timestamp 1586364061
transform 1 0 11224 0 1 49504
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_87_123
timestamp 1586364061
transform 1 0 12420 0 1 49504
box -38 -48 222 592
use scs8hd_decap_3  PHY_175
timestamp 1586364061
transform -1 0 12880 0 1 49504
box -38 -48 314 592
use scs8hd_decap_3  PHY_176
timestamp 1586364061
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use scs8hd_decap_12  FILLER_88_3
timestamp 1586364061
transform 1 0 1380 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_15
timestamp 1586364061
transform 1 0 2484 0 -1 50592
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 3956 0 -1 50592
box -38 -48 130 592
use scs8hd_decap_4  FILLER_88_27
timestamp 1586364061
transform 1 0 3588 0 -1 50592
box -38 -48 406 592
use scs8hd_decap_12  FILLER_88_32
timestamp 1586364061
transform 1 0 4048 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_44
timestamp 1586364061
transform 1 0 5152 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_56
timestamp 1586364061
transform 1 0 6256 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_68
timestamp 1586364061
transform 1 0 7360 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_80
timestamp 1586364061
transform 1 0 8464 0 -1 50592
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 9568 0 -1 50592
box -38 -48 130 592
use scs8hd_decap_12  FILLER_88_93
timestamp 1586364061
transform 1 0 9660 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_105
timestamp 1586364061
transform 1 0 10764 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_88_117
timestamp 1586364061
transform 1 0 11868 0 -1 50592
box -38 -48 774 592
use scs8hd_decap_3  PHY_177
timestamp 1586364061
transform -1 0 12880 0 -1 50592
box -38 -48 314 592
use scs8hd_decap_3  PHY_178
timestamp 1586364061
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use scs8hd_decap_12  FILLER_89_3
timestamp 1586364061
transform 1 0 1380 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_15
timestamp 1586364061
transform 1 0 2484 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_27
timestamp 1586364061
transform 1 0 3588 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_39
timestamp 1586364061
transform 1 0 4692 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_89_51
timestamp 1586364061
transform 1 0 5796 0 1 50592
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 6716 0 1 50592
box -38 -48 130 592
use scs8hd_fill_2  FILLER_89_59
timestamp 1586364061
transform 1 0 6532 0 1 50592
box -38 -48 222 592
use scs8hd_decap_12  FILLER_89_62
timestamp 1586364061
transform 1 0 6808 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_74
timestamp 1586364061
transform 1 0 7912 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_86
timestamp 1586364061
transform 1 0 9016 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_98
timestamp 1586364061
transform 1 0 10120 0 1 50592
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_565
timestamp 1586364061
transform 1 0 12328 0 1 50592
box -38 -48 130 592
use scs8hd_decap_12  FILLER_89_110
timestamp 1586364061
transform 1 0 11224 0 1 50592
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_89_123
timestamp 1586364061
transform 1 0 12420 0 1 50592
box -38 -48 222 592
use scs8hd_decap_3  PHY_179
timestamp 1586364061
transform -1 0 12880 0 1 50592
box -38 -48 314 592
use scs8hd_decap_3  PHY_180
timestamp 1586364061
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_90_3
timestamp 1586364061
transform 1 0 1380 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_15
timestamp 1586364061
transform 1 0 2484 0 -1 51680
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_566
timestamp 1586364061
transform 1 0 3956 0 -1 51680
box -38 -48 130 592
use scs8hd_decap_4  FILLER_90_27
timestamp 1586364061
transform 1 0 3588 0 -1 51680
box -38 -48 406 592
use scs8hd_decap_12  FILLER_90_32
timestamp 1586364061
transform 1 0 4048 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_44
timestamp 1586364061
transform 1 0 5152 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_56
timestamp 1586364061
transform 1 0 6256 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_68
timestamp 1586364061
transform 1 0 7360 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_80
timestamp 1586364061
transform 1 0 8464 0 -1 51680
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_567
timestamp 1586364061
transform 1 0 9568 0 -1 51680
box -38 -48 130 592
use scs8hd_decap_12  FILLER_90_93
timestamp 1586364061
transform 1 0 9660 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_105
timestamp 1586364061
transform 1 0 10764 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_90_117
timestamp 1586364061
transform 1 0 11868 0 -1 51680
box -38 -48 774 592
use scs8hd_decap_3  PHY_181
timestamp 1586364061
transform -1 0 12880 0 -1 51680
box -38 -48 314 592
use scs8hd_decap_3  PHY_182
timestamp 1586364061
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_91_3
timestamp 1586364061
transform 1 0 1380 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_15
timestamp 1586364061
transform 1 0 2484 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_27
timestamp 1586364061
transform 1 0 3588 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_39
timestamp 1586364061
transform 1 0 4692 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_91_51
timestamp 1586364061
transform 1 0 5796 0 1 51680
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_568
timestamp 1586364061
transform 1 0 6716 0 1 51680
box -38 -48 130 592
use scs8hd_fill_2  FILLER_91_59
timestamp 1586364061
transform 1 0 6532 0 1 51680
box -38 -48 222 592
use scs8hd_decap_12  FILLER_91_62
timestamp 1586364061
transform 1 0 6808 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_74
timestamp 1586364061
transform 1 0 7912 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_86
timestamp 1586364061
transform 1 0 9016 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_98
timestamp 1586364061
transform 1 0 10120 0 1 51680
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_569
timestamp 1586364061
transform 1 0 12328 0 1 51680
box -38 -48 130 592
use scs8hd_decap_12  FILLER_91_110
timestamp 1586364061
transform 1 0 11224 0 1 51680
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_91_123
timestamp 1586364061
transform 1 0 12420 0 1 51680
box -38 -48 222 592
use scs8hd_decap_3  PHY_183
timestamp 1586364061
transform -1 0 12880 0 1 51680
box -38 -48 314 592
use scs8hd_decap_3  PHY_184
timestamp 1586364061
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use scs8hd_decap_3  PHY_186
timestamp 1586364061
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use scs8hd_decap_12  FILLER_92_3
timestamp 1586364061
transform 1 0 1380 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_15
timestamp 1586364061
transform 1 0 2484 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_3
timestamp 1586364061
transform 1 0 1380 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_15
timestamp 1586364061
transform 1 0 2484 0 1 52768
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_570
timestamp 1586364061
transform 1 0 3956 0 -1 52768
box -38 -48 130 592
use scs8hd_decap_4  FILLER_92_27
timestamp 1586364061
transform 1 0 3588 0 -1 52768
box -38 -48 406 592
use scs8hd_decap_12  FILLER_92_32
timestamp 1586364061
transform 1 0 4048 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_27
timestamp 1586364061
transform 1 0 3588 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_44
timestamp 1586364061
transform 1 0 5152 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_39
timestamp 1586364061
transform 1 0 4692 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_93_51
timestamp 1586364061
transform 1 0 5796 0 1 52768
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_572
timestamp 1586364061
transform 1 0 6716 0 1 52768
box -38 -48 130 592
use scs8hd_decap_12  FILLER_92_56
timestamp 1586364061
transform 1 0 6256 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_68
timestamp 1586364061
transform 1 0 7360 0 -1 52768
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_93_59
timestamp 1586364061
transform 1 0 6532 0 1 52768
box -38 -48 222 592
use scs8hd_decap_12  FILLER_93_62
timestamp 1586364061
transform 1 0 6808 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_80
timestamp 1586364061
transform 1 0 8464 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_74
timestamp 1586364061
transform 1 0 7912 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_86
timestamp 1586364061
transform 1 0 9016 0 1 52768
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_571
timestamp 1586364061
transform 1 0 9568 0 -1 52768
box -38 -48 130 592
use scs8hd_decap_12  FILLER_92_93
timestamp 1586364061
transform 1 0 9660 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_105
timestamp 1586364061
transform 1 0 10764 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_93_98
timestamp 1586364061
transform 1 0 10120 0 1 52768
box -38 -48 774 592
use scs8hd_decap_3  FILLER_93_106
timestamp 1586364061
transform 1 0 10856 0 1 52768
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_573
timestamp 1586364061
transform 1 0 12328 0 1 52768
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 11132 0 1 52768
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 11500 0 1 52768
box -38 -48 222 592
use scs8hd_decap_8  FILLER_92_117
timestamp 1586364061
transform 1 0 11868 0 -1 52768
box -38 -48 774 592
use scs8hd_fill_2  FILLER_93_111
timestamp 1586364061
transform 1 0 11316 0 1 52768
box -38 -48 222 592
use scs8hd_decap_6  FILLER_93_115
timestamp 1586364061
transform 1 0 11684 0 1 52768
box -38 -48 590 592
use scs8hd_fill_1  FILLER_93_121
timestamp 1586364061
transform 1 0 12236 0 1 52768
box -38 -48 130 592
use scs8hd_fill_2  FILLER_93_123
timestamp 1586364061
transform 1 0 12420 0 1 52768
box -38 -48 222 592
use scs8hd_decap_3  PHY_185
timestamp 1586364061
transform -1 0 12880 0 -1 52768
box -38 -48 314 592
use scs8hd_decap_3  PHY_187
timestamp 1586364061
transform -1 0 12880 0 1 52768
box -38 -48 314 592
use scs8hd_decap_3  PHY_188
timestamp 1586364061
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use scs8hd_decap_12  FILLER_94_3
timestamp 1586364061
transform 1 0 1380 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_15
timestamp 1586364061
transform 1 0 2484 0 -1 53856
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_574
timestamp 1586364061
transform 1 0 3956 0 -1 53856
box -38 -48 130 592
use scs8hd_decap_4  FILLER_94_27
timestamp 1586364061
transform 1 0 3588 0 -1 53856
box -38 -48 406 592
use scs8hd_decap_12  FILLER_94_32
timestamp 1586364061
transform 1 0 4048 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_44
timestamp 1586364061
transform 1 0 5152 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_56
timestamp 1586364061
transform 1 0 6256 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_68
timestamp 1586364061
transform 1 0 7360 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_80
timestamp 1586364061
transform 1 0 8464 0 -1 53856
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_575
timestamp 1586364061
transform 1 0 9568 0 -1 53856
box -38 -48 130 592
use scs8hd_decap_12  FILLER_94_93
timestamp 1586364061
transform 1 0 9660 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_94_105
timestamp 1586364061
transform 1 0 10764 0 -1 53856
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 11132 0 -1 53856
box -38 -48 774 592
use scs8hd_decap_8  FILLER_94_117
timestamp 1586364061
transform 1 0 11868 0 -1 53856
box -38 -48 774 592
use scs8hd_decap_3  PHY_189
timestamp 1586364061
transform -1 0 12880 0 -1 53856
box -38 -48 314 592
use scs8hd_decap_3  PHY_190
timestamp 1586364061
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use scs8hd_decap_12  FILLER_95_3
timestamp 1586364061
transform 1 0 1380 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_15
timestamp 1586364061
transform 1 0 2484 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_27
timestamp 1586364061
transform 1 0 3588 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_39
timestamp 1586364061
transform 1 0 4692 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_95_51
timestamp 1586364061
transform 1 0 5796 0 1 53856
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_576
timestamp 1586364061
transform 1 0 6716 0 1 53856
box -38 -48 130 592
use scs8hd_fill_2  FILLER_95_59
timestamp 1586364061
transform 1 0 6532 0 1 53856
box -38 -48 222 592
use scs8hd_decap_12  FILLER_95_62
timestamp 1586364061
transform 1 0 6808 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_74
timestamp 1586364061
transform 1 0 7912 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_86
timestamp 1586364061
transform 1 0 9016 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_98
timestamp 1586364061
transform 1 0 10120 0 1 53856
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_577
timestamp 1586364061
transform 1 0 12328 0 1 53856
box -38 -48 130 592
use scs8hd_decap_12  FILLER_95_110
timestamp 1586364061
transform 1 0 11224 0 1 53856
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_95_123
timestamp 1586364061
transform 1 0 12420 0 1 53856
box -38 -48 222 592
use scs8hd_decap_3  PHY_191
timestamp 1586364061
transform -1 0 12880 0 1 53856
box -38 -48 314 592
use scs8hd_decap_3  PHY_192
timestamp 1586364061
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_96_3
timestamp 1586364061
transform 1 0 1380 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_15
timestamp 1586364061
transform 1 0 2484 0 -1 54944
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_578
timestamp 1586364061
transform 1 0 3956 0 -1 54944
box -38 -48 130 592
use scs8hd_decap_4  FILLER_96_27
timestamp 1586364061
transform 1 0 3588 0 -1 54944
box -38 -48 406 592
use scs8hd_decap_12  FILLER_96_32
timestamp 1586364061
transform 1 0 4048 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_44
timestamp 1586364061
transform 1 0 5152 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_56
timestamp 1586364061
transform 1 0 6256 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_68
timestamp 1586364061
transform 1 0 7360 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_80
timestamp 1586364061
transform 1 0 8464 0 -1 54944
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_579
timestamp 1586364061
transform 1 0 9568 0 -1 54944
box -38 -48 130 592
use scs8hd_decap_12  FILLER_96_93
timestamp 1586364061
transform 1 0 9660 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_105
timestamp 1586364061
transform 1 0 10764 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_96_117
timestamp 1586364061
transform 1 0 11868 0 -1 54944
box -38 -48 774 592
use scs8hd_decap_3  PHY_193
timestamp 1586364061
transform -1 0 12880 0 -1 54944
box -38 -48 314 592
use scs8hd_decap_3  PHY_194
timestamp 1586364061
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_97_3
timestamp 1586364061
transform 1 0 1380 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_15
timestamp 1586364061
transform 1 0 2484 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_27
timestamp 1586364061
transform 1 0 3588 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_39
timestamp 1586364061
transform 1 0 4692 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_97_51
timestamp 1586364061
transform 1 0 5796 0 1 54944
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_580
timestamp 1586364061
transform 1 0 6716 0 1 54944
box -38 -48 130 592
use scs8hd_fill_2  FILLER_97_59
timestamp 1586364061
transform 1 0 6532 0 1 54944
box -38 -48 222 592
use scs8hd_decap_12  FILLER_97_62
timestamp 1586364061
transform 1 0 6808 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_74
timestamp 1586364061
transform 1 0 7912 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_86
timestamp 1586364061
transform 1 0 9016 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_98
timestamp 1586364061
transform 1 0 10120 0 1 54944
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_581
timestamp 1586364061
transform 1 0 12328 0 1 54944
box -38 -48 130 592
use scs8hd_decap_12  FILLER_97_110
timestamp 1586364061
transform 1 0 11224 0 1 54944
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_97_123
timestamp 1586364061
transform 1 0 12420 0 1 54944
box -38 -48 222 592
use scs8hd_decap_3  PHY_195
timestamp 1586364061
transform -1 0 12880 0 1 54944
box -38 -48 314 592
use scs8hd_decap_3  PHY_196
timestamp 1586364061
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use scs8hd_decap_12  FILLER_98_3
timestamp 1586364061
transform 1 0 1380 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_15
timestamp 1586364061
transform 1 0 2484 0 -1 56032
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_582
timestamp 1586364061
transform 1 0 3956 0 -1 56032
box -38 -48 130 592
use scs8hd_decap_4  FILLER_98_27
timestamp 1586364061
transform 1 0 3588 0 -1 56032
box -38 -48 406 592
use scs8hd_decap_12  FILLER_98_32
timestamp 1586364061
transform 1 0 4048 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_44
timestamp 1586364061
transform 1 0 5152 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_56
timestamp 1586364061
transform 1 0 6256 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_68
timestamp 1586364061
transform 1 0 7360 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_80
timestamp 1586364061
transform 1 0 8464 0 -1 56032
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_583
timestamp 1586364061
transform 1 0 9568 0 -1 56032
box -38 -48 130 592
use scs8hd_decap_12  FILLER_98_93
timestamp 1586364061
transform 1 0 9660 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_105
timestamp 1586364061
transform 1 0 10764 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_98_117
timestamp 1586364061
transform 1 0 11868 0 -1 56032
box -38 -48 774 592
use scs8hd_decap_3  PHY_197
timestamp 1586364061
transform -1 0 12880 0 -1 56032
box -38 -48 314 592
use scs8hd_decap_3  PHY_198
timestamp 1586364061
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use scs8hd_decap_3  PHY_200
timestamp 1586364061
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use scs8hd_decap_12  FILLER_99_3
timestamp 1586364061
transform 1 0 1380 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_99_15
timestamp 1586364061
transform 1 0 2484 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_3
timestamp 1586364061
transform 1 0 1380 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_15
timestamp 1586364061
transform 1 0 2484 0 -1 57120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_586
timestamp 1586364061
transform 1 0 3956 0 -1 57120
box -38 -48 130 592
use scs8hd_decap_12  FILLER_99_27
timestamp 1586364061
transform 1 0 3588 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_100_27
timestamp 1586364061
transform 1 0 3588 0 -1 57120
box -38 -48 406 592
use scs8hd_decap_12  FILLER_100_32
timestamp 1586364061
transform 1 0 4048 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_99_39
timestamp 1586364061
transform 1 0 4692 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_99_51
timestamp 1586364061
transform 1 0 5796 0 1 56032
box -38 -48 774 592
use scs8hd_decap_12  FILLER_100_44
timestamp 1586364061
transform 1 0 5152 0 -1 57120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_584
timestamp 1586364061
transform 1 0 6716 0 1 56032
box -38 -48 130 592
use scs8hd_fill_2  FILLER_99_59
timestamp 1586364061
transform 1 0 6532 0 1 56032
box -38 -48 222 592
use scs8hd_decap_12  FILLER_99_62
timestamp 1586364061
transform 1 0 6808 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_56
timestamp 1586364061
transform 1 0 6256 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_68
timestamp 1586364061
transform 1 0 7360 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_99_74
timestamp 1586364061
transform 1 0 7912 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_99_86
timestamp 1586364061
transform 1 0 9016 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_80
timestamp 1586364061
transform 1 0 8464 0 -1 57120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_587
timestamp 1586364061
transform 1 0 9568 0 -1 57120
box -38 -48 130 592
use scs8hd_decap_12  FILLER_99_98
timestamp 1586364061
transform 1 0 10120 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_93
timestamp 1586364061
transform 1 0 9660 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_105
timestamp 1586364061
transform 1 0 10764 0 -1 57120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_585
timestamp 1586364061
transform 1 0 12328 0 1 56032
box -38 -48 130 592
use scs8hd_decap_12  FILLER_99_110
timestamp 1586364061
transform 1 0 11224 0 1 56032
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_99_123
timestamp 1586364061
transform 1 0 12420 0 1 56032
box -38 -48 222 592
use scs8hd_decap_8  FILLER_100_117
timestamp 1586364061
transform 1 0 11868 0 -1 57120
box -38 -48 774 592
use scs8hd_decap_3  PHY_199
timestamp 1586364061
transform -1 0 12880 0 1 56032
box -38 -48 314 592
use scs8hd_decap_3  PHY_201
timestamp 1586364061
transform -1 0 12880 0 -1 57120
box -38 -48 314 592
use scs8hd_decap_3  PHY_202
timestamp 1586364061
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use scs8hd_decap_12  FILLER_101_3
timestamp 1586364061
transform 1 0 1380 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_15
timestamp 1586364061
transform 1 0 2484 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_27
timestamp 1586364061
transform 1 0 3588 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_39
timestamp 1586364061
transform 1 0 4692 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_101_51
timestamp 1586364061
transform 1 0 5796 0 1 57120
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_588
timestamp 1586364061
transform 1 0 6716 0 1 57120
box -38 -48 130 592
use scs8hd_fill_2  FILLER_101_59
timestamp 1586364061
transform 1 0 6532 0 1 57120
box -38 -48 222 592
use scs8hd_decap_12  FILLER_101_62
timestamp 1586364061
transform 1 0 6808 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_74
timestamp 1586364061
transform 1 0 7912 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_86
timestamp 1586364061
transform 1 0 9016 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_98
timestamp 1586364061
transform 1 0 10120 0 1 57120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_589
timestamp 1586364061
transform 1 0 12328 0 1 57120
box -38 -48 130 592
use scs8hd_decap_12  FILLER_101_110
timestamp 1586364061
transform 1 0 11224 0 1 57120
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_101_123
timestamp 1586364061
transform 1 0 12420 0 1 57120
box -38 -48 222 592
use scs8hd_decap_3  PHY_203
timestamp 1586364061
transform -1 0 12880 0 1 57120
box -38 -48 314 592
use scs8hd_decap_3  PHY_204
timestamp 1586364061
transform 1 0 1104 0 -1 58208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_102_3
timestamp 1586364061
transform 1 0 1380 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_15
timestamp 1586364061
transform 1 0 2484 0 -1 58208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_590
timestamp 1586364061
transform 1 0 3956 0 -1 58208
box -38 -48 130 592
use scs8hd_decap_4  FILLER_102_27
timestamp 1586364061
transform 1 0 3588 0 -1 58208
box -38 -48 406 592
use scs8hd_decap_12  FILLER_102_32
timestamp 1586364061
transform 1 0 4048 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_44
timestamp 1586364061
transform 1 0 5152 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_56
timestamp 1586364061
transform 1 0 6256 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_68
timestamp 1586364061
transform 1 0 7360 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_80
timestamp 1586364061
transform 1 0 8464 0 -1 58208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_591
timestamp 1586364061
transform 1 0 9568 0 -1 58208
box -38 -48 130 592
use scs8hd_decap_12  FILLER_102_93
timestamp 1586364061
transform 1 0 9660 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_105
timestamp 1586364061
transform 1 0 10764 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_102_117
timestamp 1586364061
transform 1 0 11868 0 -1 58208
box -38 -48 774 592
use scs8hd_decap_3  PHY_205
timestamp 1586364061
transform -1 0 12880 0 -1 58208
box -38 -48 314 592
use scs8hd_decap_3  PHY_206
timestamp 1586364061
transform 1 0 1104 0 1 58208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_103_3
timestamp 1586364061
transform 1 0 1380 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_15
timestamp 1586364061
transform 1 0 2484 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_27
timestamp 1586364061
transform 1 0 3588 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_39
timestamp 1586364061
transform 1 0 4692 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_103_51
timestamp 1586364061
transform 1 0 5796 0 1 58208
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_592
timestamp 1586364061
transform 1 0 6716 0 1 58208
box -38 -48 130 592
use scs8hd_fill_2  FILLER_103_59
timestamp 1586364061
transform 1 0 6532 0 1 58208
box -38 -48 222 592
use scs8hd_decap_12  FILLER_103_62
timestamp 1586364061
transform 1 0 6808 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_74
timestamp 1586364061
transform 1 0 7912 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_86
timestamp 1586364061
transform 1 0 9016 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_98
timestamp 1586364061
transform 1 0 10120 0 1 58208
box -38 -48 1142 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 11224 0 1 58208
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_593
timestamp 1586364061
transform 1 0 12328 0 1 58208
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 11776 0 1 58208
box -38 -48 222 592
use scs8hd_fill_2  FILLER_103_114
timestamp 1586364061
transform 1 0 11592 0 1 58208
box -38 -48 222 592
use scs8hd_decap_4  FILLER_103_118
timestamp 1586364061
transform 1 0 11960 0 1 58208
box -38 -48 406 592
use scs8hd_fill_2  FILLER_103_123
timestamp 1586364061
transform 1 0 12420 0 1 58208
box -38 -48 222 592
use scs8hd_decap_3  PHY_207
timestamp 1586364061
transform -1 0 12880 0 1 58208
box -38 -48 314 592
use scs8hd_decap_3  PHY_208
timestamp 1586364061
transform 1 0 1104 0 -1 59296
box -38 -48 314 592
use scs8hd_decap_12  FILLER_104_3
timestamp 1586364061
transform 1 0 1380 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_15
timestamp 1586364061
transform 1 0 2484 0 -1 59296
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_594
timestamp 1586364061
transform 1 0 3956 0 -1 59296
box -38 -48 130 592
use scs8hd_decap_4  FILLER_104_27
timestamp 1586364061
transform 1 0 3588 0 -1 59296
box -38 -48 406 592
use scs8hd_decap_12  FILLER_104_32
timestamp 1586364061
transform 1 0 4048 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_44
timestamp 1586364061
transform 1 0 5152 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_56
timestamp 1586364061
transform 1 0 6256 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_68
timestamp 1586364061
transform 1 0 7360 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_80
timestamp 1586364061
transform 1 0 8464 0 -1 59296
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_595
timestamp 1586364061
transform 1 0 9568 0 -1 59296
box -38 -48 130 592
use scs8hd_decap_12  FILLER_104_93
timestamp 1586364061
transform 1 0 9660 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_105
timestamp 1586364061
transform 1 0 10764 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_104_117
timestamp 1586364061
transform 1 0 11868 0 -1 59296
box -38 -48 774 592
use scs8hd_decap_3  PHY_209
timestamp 1586364061
transform -1 0 12880 0 -1 59296
box -38 -48 314 592
use scs8hd_decap_3  PHY_210
timestamp 1586364061
transform 1 0 1104 0 1 59296
box -38 -48 314 592
use scs8hd_decap_3  PHY_212
timestamp 1586364061
transform 1 0 1104 0 -1 60384
box -38 -48 314 592
use scs8hd_decap_12  FILLER_105_3
timestamp 1586364061
transform 1 0 1380 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_105_15
timestamp 1586364061
transform 1 0 2484 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_3
timestamp 1586364061
transform 1 0 1380 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_15
timestamp 1586364061
transform 1 0 2484 0 -1 60384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_598
timestamp 1586364061
transform 1 0 3956 0 -1 60384
box -38 -48 130 592
use scs8hd_decap_12  FILLER_105_27
timestamp 1586364061
transform 1 0 3588 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_106_27
timestamp 1586364061
transform 1 0 3588 0 -1 60384
box -38 -48 406 592
use scs8hd_decap_12  FILLER_106_32
timestamp 1586364061
transform 1 0 4048 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_105_39
timestamp 1586364061
transform 1 0 4692 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_105_51
timestamp 1586364061
transform 1 0 5796 0 1 59296
box -38 -48 774 592
use scs8hd_decap_12  FILLER_106_44
timestamp 1586364061
transform 1 0 5152 0 -1 60384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_596
timestamp 1586364061
transform 1 0 6716 0 1 59296
box -38 -48 130 592
use scs8hd_fill_2  FILLER_105_59
timestamp 1586364061
transform 1 0 6532 0 1 59296
box -38 -48 222 592
use scs8hd_decap_12  FILLER_105_62
timestamp 1586364061
transform 1 0 6808 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_56
timestamp 1586364061
transform 1 0 6256 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_68
timestamp 1586364061
transform 1 0 7360 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_105_74
timestamp 1586364061
transform 1 0 7912 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_105_86
timestamp 1586364061
transform 1 0 9016 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_80
timestamp 1586364061
transform 1 0 8464 0 -1 60384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_599
timestamp 1586364061
transform 1 0 9568 0 -1 60384
box -38 -48 130 592
use scs8hd_decap_12  FILLER_105_98
timestamp 1586364061
transform 1 0 10120 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_93
timestamp 1586364061
transform 1 0 9660 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_105
timestamp 1586364061
transform 1 0 10764 0 -1 60384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_597
timestamp 1586364061
transform 1 0 12328 0 1 59296
box -38 -48 130 592
use scs8hd_decap_12  FILLER_105_110
timestamp 1586364061
transform 1 0 11224 0 1 59296
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_105_123
timestamp 1586364061
transform 1 0 12420 0 1 59296
box -38 -48 222 592
use scs8hd_decap_8  FILLER_106_117
timestamp 1586364061
transform 1 0 11868 0 -1 60384
box -38 -48 774 592
use scs8hd_decap_3  PHY_211
timestamp 1586364061
transform -1 0 12880 0 1 59296
box -38 -48 314 592
use scs8hd_decap_3  PHY_213
timestamp 1586364061
transform -1 0 12880 0 -1 60384
box -38 -48 314 592
use scs8hd_decap_3  PHY_214
timestamp 1586364061
transform 1 0 1104 0 1 60384
box -38 -48 314 592
use scs8hd_decap_12  FILLER_107_3
timestamp 1586364061
transform 1 0 1380 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_15
timestamp 1586364061
transform 1 0 2484 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_27
timestamp 1586364061
transform 1 0 3588 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_39
timestamp 1586364061
transform 1 0 4692 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_107_51
timestamp 1586364061
transform 1 0 5796 0 1 60384
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_600
timestamp 1586364061
transform 1 0 6716 0 1 60384
box -38 -48 130 592
use scs8hd_fill_2  FILLER_107_59
timestamp 1586364061
transform 1 0 6532 0 1 60384
box -38 -48 222 592
use scs8hd_decap_12  FILLER_107_62
timestamp 1586364061
transform 1 0 6808 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_74
timestamp 1586364061
transform 1 0 7912 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_86
timestamp 1586364061
transform 1 0 9016 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_98
timestamp 1586364061
transform 1 0 10120 0 1 60384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_601
timestamp 1586364061
transform 1 0 12328 0 1 60384
box -38 -48 130 592
use scs8hd_decap_12  FILLER_107_110
timestamp 1586364061
transform 1 0 11224 0 1 60384
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_107_123
timestamp 1586364061
transform 1 0 12420 0 1 60384
box -38 -48 222 592
use scs8hd_decap_3  PHY_215
timestamp 1586364061
transform -1 0 12880 0 1 60384
box -38 -48 314 592
use scs8hd_decap_3  PHY_216
timestamp 1586364061
transform 1 0 1104 0 -1 61472
box -38 -48 314 592
use scs8hd_decap_12  FILLER_108_3
timestamp 1586364061
transform 1 0 1380 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_15
timestamp 1586364061
transform 1 0 2484 0 -1 61472
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_602
timestamp 1586364061
transform 1 0 3956 0 -1 61472
box -38 -48 130 592
use scs8hd_decap_4  FILLER_108_27
timestamp 1586364061
transform 1 0 3588 0 -1 61472
box -38 -48 406 592
use scs8hd_decap_12  FILLER_108_32
timestamp 1586364061
transform 1 0 4048 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_44
timestamp 1586364061
transform 1 0 5152 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_56
timestamp 1586364061
transform 1 0 6256 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_68
timestamp 1586364061
transform 1 0 7360 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_80
timestamp 1586364061
transform 1 0 8464 0 -1 61472
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_603
timestamp 1586364061
transform 1 0 9568 0 -1 61472
box -38 -48 130 592
use scs8hd_decap_12  FILLER_108_93
timestamp 1586364061
transform 1 0 9660 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_105
timestamp 1586364061
transform 1 0 10764 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_108_117
timestamp 1586364061
transform 1 0 11868 0 -1 61472
box -38 -48 774 592
use scs8hd_decap_3  PHY_217
timestamp 1586364061
transform -1 0 12880 0 -1 61472
box -38 -48 314 592
use scs8hd_decap_3  PHY_218
timestamp 1586364061
transform 1 0 1104 0 1 61472
box -38 -48 314 592
use scs8hd_decap_12  FILLER_109_3
timestamp 1586364061
transform 1 0 1380 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_15
timestamp 1586364061
transform 1 0 2484 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_27
timestamp 1586364061
transform 1 0 3588 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_39
timestamp 1586364061
transform 1 0 4692 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_109_51
timestamp 1586364061
transform 1 0 5796 0 1 61472
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_604
timestamp 1586364061
transform 1 0 6716 0 1 61472
box -38 -48 130 592
use scs8hd_fill_2  FILLER_109_59
timestamp 1586364061
transform 1 0 6532 0 1 61472
box -38 -48 222 592
use scs8hd_decap_12  FILLER_109_62
timestamp 1586364061
transform 1 0 6808 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_74
timestamp 1586364061
transform 1 0 7912 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_86
timestamp 1586364061
transform 1 0 9016 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_98
timestamp 1586364061
transform 1 0 10120 0 1 61472
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_605
timestamp 1586364061
transform 1 0 12328 0 1 61472
box -38 -48 130 592
use scs8hd_decap_12  FILLER_109_110
timestamp 1586364061
transform 1 0 11224 0 1 61472
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_109_123
timestamp 1586364061
transform 1 0 12420 0 1 61472
box -38 -48 222 592
use scs8hd_decap_3  PHY_219
timestamp 1586364061
transform -1 0 12880 0 1 61472
box -38 -48 314 592
use scs8hd_decap_3  PHY_220
timestamp 1586364061
transform 1 0 1104 0 -1 62560
box -38 -48 314 592
use scs8hd_decap_12  FILLER_110_3
timestamp 1586364061
transform 1 0 1380 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_15
timestamp 1586364061
transform 1 0 2484 0 -1 62560
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_606
timestamp 1586364061
transform 1 0 3956 0 -1 62560
box -38 -48 130 592
use scs8hd_decap_4  FILLER_110_27
timestamp 1586364061
transform 1 0 3588 0 -1 62560
box -38 -48 406 592
use scs8hd_decap_12  FILLER_110_32
timestamp 1586364061
transform 1 0 4048 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_44
timestamp 1586364061
transform 1 0 5152 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_56
timestamp 1586364061
transform 1 0 6256 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_68
timestamp 1586364061
transform 1 0 7360 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_80
timestamp 1586364061
transform 1 0 8464 0 -1 62560
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_607
timestamp 1586364061
transform 1 0 9568 0 -1 62560
box -38 -48 130 592
use scs8hd_decap_12  FILLER_110_93
timestamp 1586364061
transform 1 0 9660 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_105
timestamp 1586364061
transform 1 0 10764 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_110_117
timestamp 1586364061
transform 1 0 11868 0 -1 62560
box -38 -48 774 592
use scs8hd_decap_3  PHY_221
timestamp 1586364061
transform -1 0 12880 0 -1 62560
box -38 -48 314 592
use scs8hd_decap_3  PHY_222
timestamp 1586364061
transform 1 0 1104 0 1 62560
box -38 -48 314 592
use scs8hd_decap_12  FILLER_111_3
timestamp 1586364061
transform 1 0 1380 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_15
timestamp 1586364061
transform 1 0 2484 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_27
timestamp 1586364061
transform 1 0 3588 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_39
timestamp 1586364061
transform 1 0 4692 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_111_51
timestamp 1586364061
transform 1 0 5796 0 1 62560
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_608
timestamp 1586364061
transform 1 0 6716 0 1 62560
box -38 -48 130 592
use scs8hd_fill_2  FILLER_111_59
timestamp 1586364061
transform 1 0 6532 0 1 62560
box -38 -48 222 592
use scs8hd_decap_12  FILLER_111_62
timestamp 1586364061
transform 1 0 6808 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_74
timestamp 1586364061
transform 1 0 7912 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_86
timestamp 1586364061
transform 1 0 9016 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_98
timestamp 1586364061
transform 1 0 10120 0 1 62560
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_609
timestamp 1586364061
transform 1 0 12328 0 1 62560
box -38 -48 130 592
use scs8hd_decap_12  FILLER_111_110
timestamp 1586364061
transform 1 0 11224 0 1 62560
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_111_123
timestamp 1586364061
transform 1 0 12420 0 1 62560
box -38 -48 222 592
use scs8hd_decap_3  PHY_223
timestamp 1586364061
transform -1 0 12880 0 1 62560
box -38 -48 314 592
use scs8hd_decap_3  PHY_224
timestamp 1586364061
transform 1 0 1104 0 -1 63648
box -38 -48 314 592
use scs8hd_decap_3  PHY_226
timestamp 1586364061
transform 1 0 1104 0 1 63648
box -38 -48 314 592
use scs8hd_decap_12  FILLER_112_3
timestamp 1586364061
transform 1 0 1380 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_15
timestamp 1586364061
transform 1 0 2484 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_3
timestamp 1586364061
transform 1 0 1380 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_15
timestamp 1586364061
transform 1 0 2484 0 1 63648
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_610
timestamp 1586364061
transform 1 0 3956 0 -1 63648
box -38 -48 130 592
use scs8hd_decap_4  FILLER_112_27
timestamp 1586364061
transform 1 0 3588 0 -1 63648
box -38 -48 406 592
use scs8hd_decap_12  FILLER_112_32
timestamp 1586364061
transform 1 0 4048 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_27
timestamp 1586364061
transform 1 0 3588 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_44
timestamp 1586364061
transform 1 0 5152 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_39
timestamp 1586364061
transform 1 0 4692 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_113_51
timestamp 1586364061
transform 1 0 5796 0 1 63648
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_612
timestamp 1586364061
transform 1 0 6716 0 1 63648
box -38 -48 130 592
use scs8hd_decap_12  FILLER_112_56
timestamp 1586364061
transform 1 0 6256 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_68
timestamp 1586364061
transform 1 0 7360 0 -1 63648
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_113_59
timestamp 1586364061
transform 1 0 6532 0 1 63648
box -38 -48 222 592
use scs8hd_decap_12  FILLER_113_62
timestamp 1586364061
transform 1 0 6808 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_80
timestamp 1586364061
transform 1 0 8464 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_74
timestamp 1586364061
transform 1 0 7912 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_86
timestamp 1586364061
transform 1 0 9016 0 1 63648
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_611
timestamp 1586364061
transform 1 0 9568 0 -1 63648
box -38 -48 130 592
use scs8hd_decap_12  FILLER_112_93
timestamp 1586364061
transform 1 0 9660 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_105
timestamp 1586364061
transform 1 0 10764 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_98
timestamp 1586364061
transform 1 0 10120 0 1 63648
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_613
timestamp 1586364061
transform 1 0 12328 0 1 63648
box -38 -48 130 592
use scs8hd_decap_8  FILLER_112_117
timestamp 1586364061
transform 1 0 11868 0 -1 63648
box -38 -48 774 592
use scs8hd_decap_12  FILLER_113_110
timestamp 1586364061
transform 1 0 11224 0 1 63648
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_113_123
timestamp 1586364061
transform 1 0 12420 0 1 63648
box -38 -48 222 592
use scs8hd_decap_3  PHY_225
timestamp 1586364061
transform -1 0 12880 0 -1 63648
box -38 -48 314 592
use scs8hd_decap_3  PHY_227
timestamp 1586364061
transform -1 0 12880 0 1 63648
box -38 -48 314 592
use scs8hd_decap_3  PHY_228
timestamp 1586364061
transform 1 0 1104 0 -1 64736
box -38 -48 314 592
use scs8hd_decap_12  FILLER_114_3
timestamp 1586364061
transform 1 0 1380 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_15
timestamp 1586364061
transform 1 0 2484 0 -1 64736
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_614
timestamp 1586364061
transform 1 0 3956 0 -1 64736
box -38 -48 130 592
use scs8hd_decap_4  FILLER_114_27
timestamp 1586364061
transform 1 0 3588 0 -1 64736
box -38 -48 406 592
use scs8hd_decap_12  FILLER_114_32
timestamp 1586364061
transform 1 0 4048 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_44
timestamp 1586364061
transform 1 0 5152 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_56
timestamp 1586364061
transform 1 0 6256 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_68
timestamp 1586364061
transform 1 0 7360 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_80
timestamp 1586364061
transform 1 0 8464 0 -1 64736
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_615
timestamp 1586364061
transform 1 0 9568 0 -1 64736
box -38 -48 130 592
use scs8hd_decap_12  FILLER_114_93
timestamp 1586364061
transform 1 0 9660 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_105
timestamp 1586364061
transform 1 0 10764 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_114_117
timestamp 1586364061
transform 1 0 11868 0 -1 64736
box -38 -48 774 592
use scs8hd_decap_3  PHY_229
timestamp 1586364061
transform -1 0 12880 0 -1 64736
box -38 -48 314 592
use scs8hd_decap_3  PHY_230
timestamp 1586364061
transform 1 0 1104 0 1 64736
box -38 -48 314 592
use scs8hd_decap_12  FILLER_115_3
timestamp 1586364061
transform 1 0 1380 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_15
timestamp 1586364061
transform 1 0 2484 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_27
timestamp 1586364061
transform 1 0 3588 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_39
timestamp 1586364061
transform 1 0 4692 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_115_51
timestamp 1586364061
transform 1 0 5796 0 1 64736
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_616
timestamp 1586364061
transform 1 0 6716 0 1 64736
box -38 -48 130 592
use scs8hd_fill_2  FILLER_115_59
timestamp 1586364061
transform 1 0 6532 0 1 64736
box -38 -48 222 592
use scs8hd_decap_12  FILLER_115_62
timestamp 1586364061
transform 1 0 6808 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_74
timestamp 1586364061
transform 1 0 7912 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_86
timestamp 1586364061
transform 1 0 9016 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_98
timestamp 1586364061
transform 1 0 10120 0 1 64736
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_617
timestamp 1586364061
transform 1 0 12328 0 1 64736
box -38 -48 130 592
use scs8hd_decap_12  FILLER_115_110
timestamp 1586364061
transform 1 0 11224 0 1 64736
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_115_123
timestamp 1586364061
transform 1 0 12420 0 1 64736
box -38 -48 222 592
use scs8hd_decap_3  PHY_231
timestamp 1586364061
transform -1 0 12880 0 1 64736
box -38 -48 314 592
use scs8hd_decap_3  PHY_232
timestamp 1586364061
transform 1 0 1104 0 -1 65824
box -38 -48 314 592
use scs8hd_decap_12  FILLER_116_3
timestamp 1586364061
transform 1 0 1380 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_15
timestamp 1586364061
transform 1 0 2484 0 -1 65824
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_618
timestamp 1586364061
transform 1 0 3956 0 -1 65824
box -38 -48 130 592
use scs8hd_decap_4  FILLER_116_27
timestamp 1586364061
transform 1 0 3588 0 -1 65824
box -38 -48 406 592
use scs8hd_decap_12  FILLER_116_32
timestamp 1586364061
transform 1 0 4048 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_44
timestamp 1586364061
transform 1 0 5152 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_56
timestamp 1586364061
transform 1 0 6256 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_68
timestamp 1586364061
transform 1 0 7360 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_80
timestamp 1586364061
transform 1 0 8464 0 -1 65824
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_619
timestamp 1586364061
transform 1 0 9568 0 -1 65824
box -38 -48 130 592
use scs8hd_decap_12  FILLER_116_93
timestamp 1586364061
transform 1 0 9660 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_105
timestamp 1586364061
transform 1 0 10764 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_116_117
timestamp 1586364061
transform 1 0 11868 0 -1 65824
box -38 -48 774 592
use scs8hd_decap_3  PHY_233
timestamp 1586364061
transform -1 0 12880 0 -1 65824
box -38 -48 314 592
use scs8hd_decap_3  PHY_234
timestamp 1586364061
transform 1 0 1104 0 1 65824
box -38 -48 314 592
use scs8hd_decap_12  FILLER_117_3
timestamp 1586364061
transform 1 0 1380 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_15
timestamp 1586364061
transform 1 0 2484 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_27
timestamp 1586364061
transform 1 0 3588 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_39
timestamp 1586364061
transform 1 0 4692 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_117_51
timestamp 1586364061
transform 1 0 5796 0 1 65824
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_620
timestamp 1586364061
transform 1 0 6716 0 1 65824
box -38 -48 130 592
use scs8hd_fill_2  FILLER_117_59
timestamp 1586364061
transform 1 0 6532 0 1 65824
box -38 -48 222 592
use scs8hd_decap_12  FILLER_117_62
timestamp 1586364061
transform 1 0 6808 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_74
timestamp 1586364061
transform 1 0 7912 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_86
timestamp 1586364061
transform 1 0 9016 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_117_98
timestamp 1586364061
transform 1 0 10120 0 1 65824
box -38 -48 774 592
use scs8hd_decap_3  FILLER_117_106
timestamp 1586364061
transform 1 0 10856 0 1 65824
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_621
timestamp 1586364061
transform 1 0 12328 0 1 65824
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 11132 0 1 65824
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 11500 0 1 65824
box -38 -48 222 592
use scs8hd_fill_2  FILLER_117_111
timestamp 1586364061
transform 1 0 11316 0 1 65824
box -38 -48 222 592
use scs8hd_decap_6  FILLER_117_115
timestamp 1586364061
transform 1 0 11684 0 1 65824
box -38 -48 590 592
use scs8hd_fill_1  FILLER_117_121
timestamp 1586364061
transform 1 0 12236 0 1 65824
box -38 -48 130 592
use scs8hd_fill_2  FILLER_117_123
timestamp 1586364061
transform 1 0 12420 0 1 65824
box -38 -48 222 592
use scs8hd_decap_3  PHY_235
timestamp 1586364061
transform -1 0 12880 0 1 65824
box -38 -48 314 592
use scs8hd_decap_3  PHY_236
timestamp 1586364061
transform 1 0 1104 0 -1 66912
box -38 -48 314 592
use scs8hd_decap_3  PHY_238
timestamp 1586364061
transform 1 0 1104 0 1 66912
box -38 -48 314 592
use scs8hd_decap_12  FILLER_118_3
timestamp 1586364061
transform 1 0 1380 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_118_15
timestamp 1586364061
transform 1 0 2484 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_3
timestamp 1586364061
transform 1 0 1380 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_15
timestamp 1586364061
transform 1 0 2484 0 1 66912
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_622
timestamp 1586364061
transform 1 0 3956 0 -1 66912
box -38 -48 130 592
use scs8hd_decap_4  FILLER_118_27
timestamp 1586364061
transform 1 0 3588 0 -1 66912
box -38 -48 406 592
use scs8hd_decap_12  FILLER_118_32
timestamp 1586364061
transform 1 0 4048 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_27
timestamp 1586364061
transform 1 0 3588 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_118_44
timestamp 1586364061
transform 1 0 5152 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_39
timestamp 1586364061
transform 1 0 4692 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_119_51
timestamp 1586364061
transform 1 0 5796 0 1 66912
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_624
timestamp 1586364061
transform 1 0 6716 0 1 66912
box -38 -48 130 592
use scs8hd_decap_12  FILLER_118_56
timestamp 1586364061
transform 1 0 6256 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_118_68
timestamp 1586364061
transform 1 0 7360 0 -1 66912
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_119_59
timestamp 1586364061
transform 1 0 6532 0 1 66912
box -38 -48 222 592
use scs8hd_decap_12  FILLER_119_62
timestamp 1586364061
transform 1 0 6808 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_118_80
timestamp 1586364061
transform 1 0 8464 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_74
timestamp 1586364061
transform 1 0 7912 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_86
timestamp 1586364061
transform 1 0 9016 0 1 66912
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_623
timestamp 1586364061
transform 1 0 9568 0 -1 66912
box -38 -48 130 592
use scs8hd_decap_12  FILLER_118_93
timestamp 1586364061
transform 1 0 9660 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_118_105
timestamp 1586364061
transform 1 0 10764 0 -1 66912
box -38 -48 406 592
use scs8hd_decap_12  FILLER_119_98
timestamp 1586364061
transform 1 0 10120 0 1 66912
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 11132 0 -1 66912
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_625
timestamp 1586364061
transform 1 0 12328 0 1 66912
box -38 -48 130 592
use scs8hd_decap_8  FILLER_118_117
timestamp 1586364061
transform 1 0 11868 0 -1 66912
box -38 -48 774 592
use scs8hd_decap_12  FILLER_119_110
timestamp 1586364061
transform 1 0 11224 0 1 66912
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_119_123
timestamp 1586364061
transform 1 0 12420 0 1 66912
box -38 -48 222 592
use scs8hd_decap_3  PHY_237
timestamp 1586364061
transform -1 0 12880 0 -1 66912
box -38 -48 314 592
use scs8hd_decap_3  PHY_239
timestamp 1586364061
transform -1 0 12880 0 1 66912
box -38 -48 314 592
use scs8hd_decap_3  PHY_240
timestamp 1586364061
transform 1 0 1104 0 -1 68000
box -38 -48 314 592
use scs8hd_decap_12  FILLER_120_3
timestamp 1586364061
transform 1 0 1380 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_15
timestamp 1586364061
transform 1 0 2484 0 -1 68000
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_626
timestamp 1586364061
transform 1 0 3956 0 -1 68000
box -38 -48 130 592
use scs8hd_decap_4  FILLER_120_27
timestamp 1586364061
transform 1 0 3588 0 -1 68000
box -38 -48 406 592
use scs8hd_decap_12  FILLER_120_32
timestamp 1586364061
transform 1 0 4048 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_44
timestamp 1586364061
transform 1 0 5152 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_56
timestamp 1586364061
transform 1 0 6256 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_68
timestamp 1586364061
transform 1 0 7360 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_80
timestamp 1586364061
transform 1 0 8464 0 -1 68000
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_627
timestamp 1586364061
transform 1 0 9568 0 -1 68000
box -38 -48 130 592
use scs8hd_decap_12  FILLER_120_93
timestamp 1586364061
transform 1 0 9660 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_105
timestamp 1586364061
transform 1 0 10764 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_120_117
timestamp 1586364061
transform 1 0 11868 0 -1 68000
box -38 -48 774 592
use scs8hd_decap_3  PHY_241
timestamp 1586364061
transform -1 0 12880 0 -1 68000
box -38 -48 314 592
use scs8hd_decap_3  PHY_242
timestamp 1586364061
transform 1 0 1104 0 1 68000
box -38 -48 314 592
use scs8hd_decap_12  FILLER_121_3
timestamp 1586364061
transform 1 0 1380 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_15
timestamp 1586364061
transform 1 0 2484 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_27
timestamp 1586364061
transform 1 0 3588 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_39
timestamp 1586364061
transform 1 0 4692 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_121_51
timestamp 1586364061
transform 1 0 5796 0 1 68000
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_628
timestamp 1586364061
transform 1 0 6716 0 1 68000
box -38 -48 130 592
use scs8hd_fill_2  FILLER_121_59
timestamp 1586364061
transform 1 0 6532 0 1 68000
box -38 -48 222 592
use scs8hd_decap_12  FILLER_121_62
timestamp 1586364061
transform 1 0 6808 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_74
timestamp 1586364061
transform 1 0 7912 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_86
timestamp 1586364061
transform 1 0 9016 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_98
timestamp 1586364061
transform 1 0 10120 0 1 68000
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_629
timestamp 1586364061
transform 1 0 12328 0 1 68000
box -38 -48 130 592
use scs8hd_decap_12  FILLER_121_110
timestamp 1586364061
transform 1 0 11224 0 1 68000
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_121_123
timestamp 1586364061
transform 1 0 12420 0 1 68000
box -38 -48 222 592
use scs8hd_decap_3  PHY_243
timestamp 1586364061
transform -1 0 12880 0 1 68000
box -38 -48 314 592
use scs8hd_decap_3  PHY_244
timestamp 1586364061
transform 1 0 1104 0 -1 69088
box -38 -48 314 592
use scs8hd_decap_12  FILLER_122_3
timestamp 1586364061
transform 1 0 1380 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_15
timestamp 1586364061
transform 1 0 2484 0 -1 69088
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_630
timestamp 1586364061
transform 1 0 3956 0 -1 69088
box -38 -48 130 592
use scs8hd_decap_4  FILLER_122_27
timestamp 1586364061
transform 1 0 3588 0 -1 69088
box -38 -48 406 592
use scs8hd_decap_12  FILLER_122_32
timestamp 1586364061
transform 1 0 4048 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_44
timestamp 1586364061
transform 1 0 5152 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_56
timestamp 1586364061
transform 1 0 6256 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_68
timestamp 1586364061
transform 1 0 7360 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_80
timestamp 1586364061
transform 1 0 8464 0 -1 69088
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_631
timestamp 1586364061
transform 1 0 9568 0 -1 69088
box -38 -48 130 592
use scs8hd_decap_12  FILLER_122_93
timestamp 1586364061
transform 1 0 9660 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_105
timestamp 1586364061
transform 1 0 10764 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_122_117
timestamp 1586364061
transform 1 0 11868 0 -1 69088
box -38 -48 774 592
use scs8hd_decap_3  PHY_245
timestamp 1586364061
transform -1 0 12880 0 -1 69088
box -38 -48 314 592
use scs8hd_decap_3  PHY_246
timestamp 1586364061
transform 1 0 1104 0 1 69088
box -38 -48 314 592
use scs8hd_decap_12  FILLER_123_3
timestamp 1586364061
transform 1 0 1380 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_15
timestamp 1586364061
transform 1 0 2484 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_27
timestamp 1586364061
transform 1 0 3588 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_39
timestamp 1586364061
transform 1 0 4692 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_123_51
timestamp 1586364061
transform 1 0 5796 0 1 69088
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_632
timestamp 1586364061
transform 1 0 6716 0 1 69088
box -38 -48 130 592
use scs8hd_fill_2  FILLER_123_59
timestamp 1586364061
transform 1 0 6532 0 1 69088
box -38 -48 222 592
use scs8hd_decap_12  FILLER_123_62
timestamp 1586364061
transform 1 0 6808 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_74
timestamp 1586364061
transform 1 0 7912 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_86
timestamp 1586364061
transform 1 0 9016 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_98
timestamp 1586364061
transform 1 0 10120 0 1 69088
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_633
timestamp 1586364061
transform 1 0 12328 0 1 69088
box -38 -48 130 592
use scs8hd_decap_12  FILLER_123_110
timestamp 1586364061
transform 1 0 11224 0 1 69088
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_123_123
timestamp 1586364061
transform 1 0 12420 0 1 69088
box -38 -48 222 592
use scs8hd_decap_3  PHY_247
timestamp 1586364061
transform -1 0 12880 0 1 69088
box -38 -48 314 592
use scs8hd_decap_3  PHY_248
timestamp 1586364061
transform 1 0 1104 0 -1 70176
box -38 -48 314 592
use scs8hd_decap_12  FILLER_124_3
timestamp 1586364061
transform 1 0 1380 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_15
timestamp 1586364061
transform 1 0 2484 0 -1 70176
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_634
timestamp 1586364061
transform 1 0 3956 0 -1 70176
box -38 -48 130 592
use scs8hd_decap_4  FILLER_124_27
timestamp 1586364061
transform 1 0 3588 0 -1 70176
box -38 -48 406 592
use scs8hd_decap_12  FILLER_124_32
timestamp 1586364061
transform 1 0 4048 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_44
timestamp 1586364061
transform 1 0 5152 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_56
timestamp 1586364061
transform 1 0 6256 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_68
timestamp 1586364061
transform 1 0 7360 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_80
timestamp 1586364061
transform 1 0 8464 0 -1 70176
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_635
timestamp 1586364061
transform 1 0 9568 0 -1 70176
box -38 -48 130 592
use scs8hd_decap_12  FILLER_124_93
timestamp 1586364061
transform 1 0 9660 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_105
timestamp 1586364061
transform 1 0 10764 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_124_117
timestamp 1586364061
transform 1 0 11868 0 -1 70176
box -38 -48 774 592
use scs8hd_decap_3  PHY_249
timestamp 1586364061
transform -1 0 12880 0 -1 70176
box -38 -48 314 592
use scs8hd_decap_3  PHY_250
timestamp 1586364061
transform 1 0 1104 0 1 70176
box -38 -48 314 592
use scs8hd_decap_3  PHY_252
timestamp 1586364061
transform 1 0 1104 0 -1 71264
box -38 -48 314 592
use scs8hd_decap_12  FILLER_125_3
timestamp 1586364061
transform 1 0 1380 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_125_15
timestamp 1586364061
transform 1 0 2484 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_3
timestamp 1586364061
transform 1 0 1380 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_15
timestamp 1586364061
transform 1 0 2484 0 -1 71264
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_638
timestamp 1586364061
transform 1 0 3956 0 -1 71264
box -38 -48 130 592
use scs8hd_decap_12  FILLER_125_27
timestamp 1586364061
transform 1 0 3588 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_126_27
timestamp 1586364061
transform 1 0 3588 0 -1 71264
box -38 -48 406 592
use scs8hd_decap_12  FILLER_126_32
timestamp 1586364061
transform 1 0 4048 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_125_39
timestamp 1586364061
transform 1 0 4692 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_125_51
timestamp 1586364061
transform 1 0 5796 0 1 70176
box -38 -48 774 592
use scs8hd_decap_12  FILLER_126_44
timestamp 1586364061
transform 1 0 5152 0 -1 71264
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_636
timestamp 1586364061
transform 1 0 6716 0 1 70176
box -38 -48 130 592
use scs8hd_fill_2  FILLER_125_59
timestamp 1586364061
transform 1 0 6532 0 1 70176
box -38 -48 222 592
use scs8hd_decap_12  FILLER_125_62
timestamp 1586364061
transform 1 0 6808 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_56
timestamp 1586364061
transform 1 0 6256 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_68
timestamp 1586364061
transform 1 0 7360 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_125_74
timestamp 1586364061
transform 1 0 7912 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_125_86
timestamp 1586364061
transform 1 0 9016 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_80
timestamp 1586364061
transform 1 0 8464 0 -1 71264
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_639
timestamp 1586364061
transform 1 0 9568 0 -1 71264
box -38 -48 130 592
use scs8hd_decap_12  FILLER_125_98
timestamp 1586364061
transform 1 0 10120 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_93
timestamp 1586364061
transform 1 0 9660 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_105
timestamp 1586364061
transform 1 0 10764 0 -1 71264
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_637
timestamp 1586364061
transform 1 0 12328 0 1 70176
box -38 -48 130 592
use scs8hd_decap_12  FILLER_125_110
timestamp 1586364061
transform 1 0 11224 0 1 70176
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_125_123
timestamp 1586364061
transform 1 0 12420 0 1 70176
box -38 -48 222 592
use scs8hd_decap_8  FILLER_126_117
timestamp 1586364061
transform 1 0 11868 0 -1 71264
box -38 -48 774 592
use scs8hd_decap_3  PHY_251
timestamp 1586364061
transform -1 0 12880 0 1 70176
box -38 -48 314 592
use scs8hd_decap_3  PHY_253
timestamp 1586364061
transform -1 0 12880 0 -1 71264
box -38 -48 314 592
use scs8hd_decap_3  PHY_254
timestamp 1586364061
transform 1 0 1104 0 1 71264
box -38 -48 314 592
use scs8hd_decap_12  FILLER_127_3
timestamp 1586364061
transform 1 0 1380 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_15
timestamp 1586364061
transform 1 0 2484 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_27
timestamp 1586364061
transform 1 0 3588 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_39
timestamp 1586364061
transform 1 0 4692 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_127_51
timestamp 1586364061
transform 1 0 5796 0 1 71264
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_640
timestamp 1586364061
transform 1 0 6716 0 1 71264
box -38 -48 130 592
use scs8hd_fill_2  FILLER_127_59
timestamp 1586364061
transform 1 0 6532 0 1 71264
box -38 -48 222 592
use scs8hd_decap_12  FILLER_127_62
timestamp 1586364061
transform 1 0 6808 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_74
timestamp 1586364061
transform 1 0 7912 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_86
timestamp 1586364061
transform 1 0 9016 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_98
timestamp 1586364061
transform 1 0 10120 0 1 71264
box -38 -48 1142 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 11224 0 1 71264
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_641
timestamp 1586364061
transform 1 0 12328 0 1 71264
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 11776 0 1 71264
box -38 -48 222 592
use scs8hd_fill_2  FILLER_127_114
timestamp 1586364061
transform 1 0 11592 0 1 71264
box -38 -48 222 592
use scs8hd_decap_4  FILLER_127_118
timestamp 1586364061
transform 1 0 11960 0 1 71264
box -38 -48 406 592
use scs8hd_fill_2  FILLER_127_123
timestamp 1586364061
transform 1 0 12420 0 1 71264
box -38 -48 222 592
use scs8hd_decap_3  PHY_255
timestamp 1586364061
transform -1 0 12880 0 1 71264
box -38 -48 314 592
use scs8hd_decap_3  PHY_256
timestamp 1586364061
transform 1 0 1104 0 -1 72352
box -38 -48 314 592
use scs8hd_decap_12  FILLER_128_3
timestamp 1586364061
transform 1 0 1380 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_15
timestamp 1586364061
transform 1 0 2484 0 -1 72352
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_642
timestamp 1586364061
transform 1 0 3956 0 -1 72352
box -38 -48 130 592
use scs8hd_decap_4  FILLER_128_27
timestamp 1586364061
transform 1 0 3588 0 -1 72352
box -38 -48 406 592
use scs8hd_decap_12  FILLER_128_32
timestamp 1586364061
transform 1 0 4048 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_44
timestamp 1586364061
transform 1 0 5152 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_56
timestamp 1586364061
transform 1 0 6256 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_68
timestamp 1586364061
transform 1 0 7360 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_80
timestamp 1586364061
transform 1 0 8464 0 -1 72352
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_643
timestamp 1586364061
transform 1 0 9568 0 -1 72352
box -38 -48 130 592
use scs8hd_decap_12  FILLER_128_93
timestamp 1586364061
transform 1 0 9660 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_105
timestamp 1586364061
transform 1 0 10764 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_128_117
timestamp 1586364061
transform 1 0 11868 0 -1 72352
box -38 -48 774 592
use scs8hd_decap_3  PHY_257
timestamp 1586364061
transform -1 0 12880 0 -1 72352
box -38 -48 314 592
use scs8hd_decap_3  PHY_258
timestamp 1586364061
transform 1 0 1104 0 1 72352
box -38 -48 314 592
use scs8hd_decap_12  FILLER_129_3
timestamp 1586364061
transform 1 0 1380 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_15
timestamp 1586364061
transform 1 0 2484 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_27
timestamp 1586364061
transform 1 0 3588 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_39
timestamp 1586364061
transform 1 0 4692 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_129_51
timestamp 1586364061
transform 1 0 5796 0 1 72352
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_644
timestamp 1586364061
transform 1 0 6716 0 1 72352
box -38 -48 130 592
use scs8hd_fill_2  FILLER_129_59
timestamp 1586364061
transform 1 0 6532 0 1 72352
box -38 -48 222 592
use scs8hd_decap_12  FILLER_129_62
timestamp 1586364061
transform 1 0 6808 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_74
timestamp 1586364061
transform 1 0 7912 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_86
timestamp 1586364061
transform 1 0 9016 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_98
timestamp 1586364061
transform 1 0 10120 0 1 72352
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_645
timestamp 1586364061
transform 1 0 12328 0 1 72352
box -38 -48 130 592
use scs8hd_decap_12  FILLER_129_110
timestamp 1586364061
transform 1 0 11224 0 1 72352
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_129_123
timestamp 1586364061
transform 1 0 12420 0 1 72352
box -38 -48 222 592
use scs8hd_decap_3  PHY_259
timestamp 1586364061
transform -1 0 12880 0 1 72352
box -38 -48 314 592
use scs8hd_decap_3  PHY_260
timestamp 1586364061
transform 1 0 1104 0 -1 73440
box -38 -48 314 592
use scs8hd_decap_12  FILLER_130_3
timestamp 1586364061
transform 1 0 1380 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_15
timestamp 1586364061
transform 1 0 2484 0 -1 73440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_646
timestamp 1586364061
transform 1 0 3956 0 -1 73440
box -38 -48 130 592
use scs8hd_decap_4  FILLER_130_27
timestamp 1586364061
transform 1 0 3588 0 -1 73440
box -38 -48 406 592
use scs8hd_decap_12  FILLER_130_32
timestamp 1586364061
transform 1 0 4048 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_44
timestamp 1586364061
transform 1 0 5152 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_56
timestamp 1586364061
transform 1 0 6256 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_68
timestamp 1586364061
transform 1 0 7360 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_80
timestamp 1586364061
transform 1 0 8464 0 -1 73440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_647
timestamp 1586364061
transform 1 0 9568 0 -1 73440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_130_93
timestamp 1586364061
transform 1 0 9660 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_105
timestamp 1586364061
transform 1 0 10764 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_130_117
timestamp 1586364061
transform 1 0 11868 0 -1 73440
box -38 -48 774 592
use scs8hd_decap_3  PHY_261
timestamp 1586364061
transform -1 0 12880 0 -1 73440
box -38 -48 314 592
use scs8hd_decap_3  PHY_262
timestamp 1586364061
transform 1 0 1104 0 1 73440
box -38 -48 314 592
use scs8hd_decap_12  FILLER_131_3
timestamp 1586364061
transform 1 0 1380 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_15
timestamp 1586364061
transform 1 0 2484 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_27
timestamp 1586364061
transform 1 0 3588 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_39
timestamp 1586364061
transform 1 0 4692 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_131_51
timestamp 1586364061
transform 1 0 5796 0 1 73440
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_648
timestamp 1586364061
transform 1 0 6716 0 1 73440
box -38 -48 130 592
use scs8hd_fill_2  FILLER_131_59
timestamp 1586364061
transform 1 0 6532 0 1 73440
box -38 -48 222 592
use scs8hd_decap_12  FILLER_131_62
timestamp 1586364061
transform 1 0 6808 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_74
timestamp 1586364061
transform 1 0 7912 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_86
timestamp 1586364061
transform 1 0 9016 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_98
timestamp 1586364061
transform 1 0 10120 0 1 73440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_649
timestamp 1586364061
transform 1 0 12328 0 1 73440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_131_110
timestamp 1586364061
transform 1 0 11224 0 1 73440
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_131_123
timestamp 1586364061
transform 1 0 12420 0 1 73440
box -38 -48 222 592
use scs8hd_decap_3  PHY_263
timestamp 1586364061
transform -1 0 12880 0 1 73440
box -38 -48 314 592
use scs8hd_decap_3  PHY_264
timestamp 1586364061
transform 1 0 1104 0 -1 74528
box -38 -48 314 592
use scs8hd_decap_3  PHY_266
timestamp 1586364061
transform 1 0 1104 0 1 74528
box -38 -48 314 592
use scs8hd_decap_12  FILLER_132_3
timestamp 1586364061
transform 1 0 1380 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_15
timestamp 1586364061
transform 1 0 2484 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_3
timestamp 1586364061
transform 1 0 1380 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_15
timestamp 1586364061
transform 1 0 2484 0 1 74528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_650
timestamp 1586364061
transform 1 0 3956 0 -1 74528
box -38 -48 130 592
use scs8hd_decap_4  FILLER_132_27
timestamp 1586364061
transform 1 0 3588 0 -1 74528
box -38 -48 406 592
use scs8hd_decap_12  FILLER_132_32
timestamp 1586364061
transform 1 0 4048 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_27
timestamp 1586364061
transform 1 0 3588 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_44
timestamp 1586364061
transform 1 0 5152 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_39
timestamp 1586364061
transform 1 0 4692 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_133_51
timestamp 1586364061
transform 1 0 5796 0 1 74528
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_652
timestamp 1586364061
transform 1 0 6716 0 1 74528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_132_56
timestamp 1586364061
transform 1 0 6256 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_68
timestamp 1586364061
transform 1 0 7360 0 -1 74528
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_133_59
timestamp 1586364061
transform 1 0 6532 0 1 74528
box -38 -48 222 592
use scs8hd_decap_12  FILLER_133_62
timestamp 1586364061
transform 1 0 6808 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_80
timestamp 1586364061
transform 1 0 8464 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_74
timestamp 1586364061
transform 1 0 7912 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_86
timestamp 1586364061
transform 1 0 9016 0 1 74528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_651
timestamp 1586364061
transform 1 0 9568 0 -1 74528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_132_93
timestamp 1586364061
transform 1 0 9660 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_105
timestamp 1586364061
transform 1 0 10764 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_98
timestamp 1586364061
transform 1 0 10120 0 1 74528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_653
timestamp 1586364061
transform 1 0 12328 0 1 74528
box -38 -48 130 592
use scs8hd_decap_8  FILLER_132_117
timestamp 1586364061
transform 1 0 11868 0 -1 74528
box -38 -48 774 592
use scs8hd_decap_12  FILLER_133_110
timestamp 1586364061
transform 1 0 11224 0 1 74528
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_133_123
timestamp 1586364061
transform 1 0 12420 0 1 74528
box -38 -48 222 592
use scs8hd_decap_3  PHY_265
timestamp 1586364061
transform -1 0 12880 0 -1 74528
box -38 -48 314 592
use scs8hd_decap_3  PHY_267
timestamp 1586364061
transform -1 0 12880 0 1 74528
box -38 -48 314 592
use scs8hd_decap_3  PHY_268
timestamp 1586364061
transform 1 0 1104 0 -1 75616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_134_3
timestamp 1586364061
transform 1 0 1380 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_15
timestamp 1586364061
transform 1 0 2484 0 -1 75616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_654
timestamp 1586364061
transform 1 0 3956 0 -1 75616
box -38 -48 130 592
use scs8hd_decap_4  FILLER_134_27
timestamp 1586364061
transform 1 0 3588 0 -1 75616
box -38 -48 406 592
use scs8hd_decap_12  FILLER_134_32
timestamp 1586364061
transform 1 0 4048 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_44
timestamp 1586364061
transform 1 0 5152 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_56
timestamp 1586364061
transform 1 0 6256 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_68
timestamp 1586364061
transform 1 0 7360 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_80
timestamp 1586364061
transform 1 0 8464 0 -1 75616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_655
timestamp 1586364061
transform 1 0 9568 0 -1 75616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_134_93
timestamp 1586364061
transform 1 0 9660 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_105
timestamp 1586364061
transform 1 0 10764 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_134_117
timestamp 1586364061
transform 1 0 11868 0 -1 75616
box -38 -48 774 592
use scs8hd_decap_3  PHY_269
timestamp 1586364061
transform -1 0 12880 0 -1 75616
box -38 -48 314 592
use scs8hd_decap_3  PHY_270
timestamp 1586364061
transform 1 0 1104 0 1 75616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_135_3
timestamp 1586364061
transform 1 0 1380 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_15
timestamp 1586364061
transform 1 0 2484 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_27
timestamp 1586364061
transform 1 0 3588 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_39
timestamp 1586364061
transform 1 0 4692 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_135_51
timestamp 1586364061
transform 1 0 5796 0 1 75616
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_656
timestamp 1586364061
transform 1 0 6716 0 1 75616
box -38 -48 130 592
use scs8hd_fill_2  FILLER_135_59
timestamp 1586364061
transform 1 0 6532 0 1 75616
box -38 -48 222 592
use scs8hd_decap_12  FILLER_135_62
timestamp 1586364061
transform 1 0 6808 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_74
timestamp 1586364061
transform 1 0 7912 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_86
timestamp 1586364061
transform 1 0 9016 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_98
timestamp 1586364061
transform 1 0 10120 0 1 75616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_657
timestamp 1586364061
transform 1 0 12328 0 1 75616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_135_110
timestamp 1586364061
transform 1 0 11224 0 1 75616
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_135_123
timestamp 1586364061
transform 1 0 12420 0 1 75616
box -38 -48 222 592
use scs8hd_decap_3  PHY_271
timestamp 1586364061
transform -1 0 12880 0 1 75616
box -38 -48 314 592
use scs8hd_decap_3  PHY_272
timestamp 1586364061
transform 1 0 1104 0 -1 76704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_136_3
timestamp 1586364061
transform 1 0 1380 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_15
timestamp 1586364061
transform 1 0 2484 0 -1 76704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_658
timestamp 1586364061
transform 1 0 3956 0 -1 76704
box -38 -48 130 592
use scs8hd_decap_4  FILLER_136_27
timestamp 1586364061
transform 1 0 3588 0 -1 76704
box -38 -48 406 592
use scs8hd_decap_12  FILLER_136_32
timestamp 1586364061
transform 1 0 4048 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_44
timestamp 1586364061
transform 1 0 5152 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_56
timestamp 1586364061
transform 1 0 6256 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_68
timestamp 1586364061
transform 1 0 7360 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_80
timestamp 1586364061
transform 1 0 8464 0 -1 76704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_659
timestamp 1586364061
transform 1 0 9568 0 -1 76704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_136_93
timestamp 1586364061
transform 1 0 9660 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_105
timestamp 1586364061
transform 1 0 10764 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_136_117
timestamp 1586364061
transform 1 0 11868 0 -1 76704
box -38 -48 774 592
use scs8hd_decap_3  PHY_273
timestamp 1586364061
transform -1 0 12880 0 -1 76704
box -38 -48 314 592
use scs8hd_decap_3  PHY_274
timestamp 1586364061
transform 1 0 1104 0 1 76704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_137_3
timestamp 1586364061
transform 1 0 1380 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_15
timestamp 1586364061
transform 1 0 2484 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_27
timestamp 1586364061
transform 1 0 3588 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_39
timestamp 1586364061
transform 1 0 4692 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_137_51
timestamp 1586364061
transform 1 0 5796 0 1 76704
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_660
timestamp 1586364061
transform 1 0 6716 0 1 76704
box -38 -48 130 592
use scs8hd_fill_2  FILLER_137_59
timestamp 1586364061
transform 1 0 6532 0 1 76704
box -38 -48 222 592
use scs8hd_decap_12  FILLER_137_62
timestamp 1586364061
transform 1 0 6808 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_74
timestamp 1586364061
transform 1 0 7912 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_86
timestamp 1586364061
transform 1 0 9016 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_98
timestamp 1586364061
transform 1 0 10120 0 1 76704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_661
timestamp 1586364061
transform 1 0 12328 0 1 76704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_137_110
timestamp 1586364061
transform 1 0 11224 0 1 76704
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_137_123
timestamp 1586364061
transform 1 0 12420 0 1 76704
box -38 -48 222 592
use scs8hd_decap_3  PHY_275
timestamp 1586364061
transform -1 0 12880 0 1 76704
box -38 -48 314 592
use scs8hd_decap_3  PHY_276
timestamp 1586364061
transform 1 0 1104 0 -1 77792
box -38 -48 314 592
use scs8hd_decap_3  PHY_278
timestamp 1586364061
transform 1 0 1104 0 1 77792
box -38 -48 314 592
use scs8hd_decap_12  FILLER_138_3
timestamp 1586364061
transform 1 0 1380 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_15
timestamp 1586364061
transform 1 0 2484 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_3
timestamp 1586364061
transform 1 0 1380 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_15
timestamp 1586364061
transform 1 0 2484 0 1 77792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_662
timestamp 1586364061
transform 1 0 3956 0 -1 77792
box -38 -48 130 592
use scs8hd_decap_4  FILLER_138_27
timestamp 1586364061
transform 1 0 3588 0 -1 77792
box -38 -48 406 592
use scs8hd_decap_12  FILLER_138_32
timestamp 1586364061
transform 1 0 4048 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_27
timestamp 1586364061
transform 1 0 3588 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_44
timestamp 1586364061
transform 1 0 5152 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_39
timestamp 1586364061
transform 1 0 4692 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_139_51
timestamp 1586364061
transform 1 0 5796 0 1 77792
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_664
timestamp 1586364061
transform 1 0 6716 0 1 77792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_138_56
timestamp 1586364061
transform 1 0 6256 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_68
timestamp 1586364061
transform 1 0 7360 0 -1 77792
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_139_59
timestamp 1586364061
transform 1 0 6532 0 1 77792
box -38 -48 222 592
use scs8hd_decap_12  FILLER_139_62
timestamp 1586364061
transform 1 0 6808 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_80
timestamp 1586364061
transform 1 0 8464 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_74
timestamp 1586364061
transform 1 0 7912 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_86
timestamp 1586364061
transform 1 0 9016 0 1 77792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_663
timestamp 1586364061
transform 1 0 9568 0 -1 77792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_138_93
timestamp 1586364061
transform 1 0 9660 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_105
timestamp 1586364061
transform 1 0 10764 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_98
timestamp 1586364061
transform 1 0 10120 0 1 77792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_665
timestamp 1586364061
transform 1 0 12328 0 1 77792
box -38 -48 130 592
use scs8hd_decap_8  FILLER_138_117
timestamp 1586364061
transform 1 0 11868 0 -1 77792
box -38 -48 774 592
use scs8hd_decap_12  FILLER_139_110
timestamp 1586364061
transform 1 0 11224 0 1 77792
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_139_123
timestamp 1586364061
transform 1 0 12420 0 1 77792
box -38 -48 222 592
use scs8hd_decap_3  PHY_277
timestamp 1586364061
transform -1 0 12880 0 -1 77792
box -38 -48 314 592
use scs8hd_decap_3  PHY_279
timestamp 1586364061
transform -1 0 12880 0 1 77792
box -38 -48 314 592
use scs8hd_decap_3  PHY_280
timestamp 1586364061
transform 1 0 1104 0 -1 78880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_140_3
timestamp 1586364061
transform 1 0 1380 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_15
timestamp 1586364061
transform 1 0 2484 0 -1 78880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_666
timestamp 1586364061
transform 1 0 3956 0 -1 78880
box -38 -48 130 592
use scs8hd_decap_4  FILLER_140_27
timestamp 1586364061
transform 1 0 3588 0 -1 78880
box -38 -48 406 592
use scs8hd_decap_12  FILLER_140_32
timestamp 1586364061
transform 1 0 4048 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_44
timestamp 1586364061
transform 1 0 5152 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_56
timestamp 1586364061
transform 1 0 6256 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_68
timestamp 1586364061
transform 1 0 7360 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_80
timestamp 1586364061
transform 1 0 8464 0 -1 78880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_667
timestamp 1586364061
transform 1 0 9568 0 -1 78880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_140_93
timestamp 1586364061
transform 1 0 9660 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_105
timestamp 1586364061
transform 1 0 10764 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_140_117
timestamp 1586364061
transform 1 0 11868 0 -1 78880
box -38 -48 774 592
use scs8hd_decap_3  PHY_281
timestamp 1586364061
transform -1 0 12880 0 -1 78880
box -38 -48 314 592
use scs8hd_decap_3  PHY_282
timestamp 1586364061
transform 1 0 1104 0 1 78880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_141_3
timestamp 1586364061
transform 1 0 1380 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_15
timestamp 1586364061
transform 1 0 2484 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_27
timestamp 1586364061
transform 1 0 3588 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_39
timestamp 1586364061
transform 1 0 4692 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_141_51
timestamp 1586364061
transform 1 0 5796 0 1 78880
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_668
timestamp 1586364061
transform 1 0 6716 0 1 78880
box -38 -48 130 592
use scs8hd_fill_2  FILLER_141_59
timestamp 1586364061
transform 1 0 6532 0 1 78880
box -38 -48 222 592
use scs8hd_decap_12  FILLER_141_62
timestamp 1586364061
transform 1 0 6808 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_74
timestamp 1586364061
transform 1 0 7912 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_86
timestamp 1586364061
transform 1 0 9016 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_98
timestamp 1586364061
transform 1 0 10120 0 1 78880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_669
timestamp 1586364061
transform 1 0 12328 0 1 78880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_141_110
timestamp 1586364061
transform 1 0 11224 0 1 78880
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_141_123
timestamp 1586364061
transform 1 0 12420 0 1 78880
box -38 -48 222 592
use scs8hd_decap_3  PHY_283
timestamp 1586364061
transform -1 0 12880 0 1 78880
box -38 -48 314 592
use scs8hd_decap_3  PHY_284
timestamp 1586364061
transform 1 0 1104 0 -1 79968
box -38 -48 314 592
use scs8hd_decap_12  FILLER_142_3
timestamp 1586364061
transform 1 0 1380 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_15
timestamp 1586364061
transform 1 0 2484 0 -1 79968
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_670
timestamp 1586364061
transform 1 0 3956 0 -1 79968
box -38 -48 130 592
use scs8hd_decap_4  FILLER_142_27
timestamp 1586364061
transform 1 0 3588 0 -1 79968
box -38 -48 406 592
use scs8hd_decap_12  FILLER_142_32
timestamp 1586364061
transform 1 0 4048 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_44
timestamp 1586364061
transform 1 0 5152 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_56
timestamp 1586364061
transform 1 0 6256 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_68
timestamp 1586364061
transform 1 0 7360 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_80
timestamp 1586364061
transform 1 0 8464 0 -1 79968
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_671
timestamp 1586364061
transform 1 0 9568 0 -1 79968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_142_93
timestamp 1586364061
transform 1 0 9660 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_105
timestamp 1586364061
transform 1 0 10764 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_142_117
timestamp 1586364061
transform 1 0 11868 0 -1 79968
box -38 -48 774 592
use scs8hd_decap_3  PHY_285
timestamp 1586364061
transform -1 0 12880 0 -1 79968
box -38 -48 314 592
use scs8hd_decap_3  PHY_286
timestamp 1586364061
transform 1 0 1104 0 1 79968
box -38 -48 314 592
use scs8hd_decap_12  FILLER_143_3
timestamp 1586364061
transform 1 0 1380 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_15
timestamp 1586364061
transform 1 0 2484 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_27
timestamp 1586364061
transform 1 0 3588 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_39
timestamp 1586364061
transform 1 0 4692 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_143_51
timestamp 1586364061
transform 1 0 5796 0 1 79968
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_672
timestamp 1586364061
transform 1 0 6716 0 1 79968
box -38 -48 130 592
use scs8hd_fill_2  FILLER_143_59
timestamp 1586364061
transform 1 0 6532 0 1 79968
box -38 -48 222 592
use scs8hd_decap_12  FILLER_143_62
timestamp 1586364061
transform 1 0 6808 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_74
timestamp 1586364061
transform 1 0 7912 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_86
timestamp 1586364061
transform 1 0 9016 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_143_98
timestamp 1586364061
transform 1 0 10120 0 1 79968
box -38 -48 774 592
use scs8hd_decap_3  FILLER_143_106
timestamp 1586364061
transform 1 0 10856 0 1 79968
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_673
timestamp 1586364061
transform 1 0 12328 0 1 79968
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 11132 0 1 79968
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 11500 0 1 79968
box -38 -48 222 592
use scs8hd_fill_2  FILLER_143_111
timestamp 1586364061
transform 1 0 11316 0 1 79968
box -38 -48 222 592
use scs8hd_decap_6  FILLER_143_115
timestamp 1586364061
transform 1 0 11684 0 1 79968
box -38 -48 590 592
use scs8hd_fill_1  FILLER_143_121
timestamp 1586364061
transform 1 0 12236 0 1 79968
box -38 -48 130 592
use scs8hd_fill_2  FILLER_143_123
timestamp 1586364061
transform 1 0 12420 0 1 79968
box -38 -48 222 592
use scs8hd_decap_3  PHY_287
timestamp 1586364061
transform -1 0 12880 0 1 79968
box -38 -48 314 592
use scs8hd_decap_3  PHY_288
timestamp 1586364061
transform 1 0 1104 0 -1 81056
box -38 -48 314 592
use scs8hd_decap_12  FILLER_144_3
timestamp 1586364061
transform 1 0 1380 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_15
timestamp 1586364061
transform 1 0 2484 0 -1 81056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_674
timestamp 1586364061
transform 1 0 3956 0 -1 81056
box -38 -48 130 592
use scs8hd_decap_4  FILLER_144_27
timestamp 1586364061
transform 1 0 3588 0 -1 81056
box -38 -48 406 592
use scs8hd_decap_12  FILLER_144_32
timestamp 1586364061
transform 1 0 4048 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_44
timestamp 1586364061
transform 1 0 5152 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_56
timestamp 1586364061
transform 1 0 6256 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_68
timestamp 1586364061
transform 1 0 7360 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_80
timestamp 1586364061
transform 1 0 8464 0 -1 81056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_675
timestamp 1586364061
transform 1 0 9568 0 -1 81056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_144_93
timestamp 1586364061
transform 1 0 9660 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_144_105
timestamp 1586364061
transform 1 0 10764 0 -1 81056
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 11132 0 -1 81056
box -38 -48 774 592
use scs8hd_decap_8  FILLER_144_117
timestamp 1586364061
transform 1 0 11868 0 -1 81056
box -38 -48 774 592
use scs8hd_decap_3  PHY_289
timestamp 1586364061
transform -1 0 12880 0 -1 81056
box -38 -48 314 592
use scs8hd_decap_3  PHY_290
timestamp 1586364061
transform 1 0 1104 0 1 81056
box -38 -48 314 592
use scs8hd_decap_3  PHY_292
timestamp 1586364061
transform 1 0 1104 0 -1 82144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_145_3
timestamp 1586364061
transform 1 0 1380 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_145_15
timestamp 1586364061
transform 1 0 2484 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_3
timestamp 1586364061
transform 1 0 1380 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_15
timestamp 1586364061
transform 1 0 2484 0 -1 82144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_678
timestamp 1586364061
transform 1 0 3956 0 -1 82144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_145_27
timestamp 1586364061
transform 1 0 3588 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_146_27
timestamp 1586364061
transform 1 0 3588 0 -1 82144
box -38 -48 406 592
use scs8hd_decap_12  FILLER_146_32
timestamp 1586364061
transform 1 0 4048 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_145_39
timestamp 1586364061
transform 1 0 4692 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_145_51
timestamp 1586364061
transform 1 0 5796 0 1 81056
box -38 -48 774 592
use scs8hd_decap_12  FILLER_146_44
timestamp 1586364061
transform 1 0 5152 0 -1 82144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_676
timestamp 1586364061
transform 1 0 6716 0 1 81056
box -38 -48 130 592
use scs8hd_fill_2  FILLER_145_59
timestamp 1586364061
transform 1 0 6532 0 1 81056
box -38 -48 222 592
use scs8hd_decap_12  FILLER_145_62
timestamp 1586364061
transform 1 0 6808 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_56
timestamp 1586364061
transform 1 0 6256 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_68
timestamp 1586364061
transform 1 0 7360 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_145_74
timestamp 1586364061
transform 1 0 7912 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_145_86
timestamp 1586364061
transform 1 0 9016 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_80
timestamp 1586364061
transform 1 0 8464 0 -1 82144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_679
timestamp 1586364061
transform 1 0 9568 0 -1 82144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_145_98
timestamp 1586364061
transform 1 0 10120 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_93
timestamp 1586364061
transform 1 0 9660 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_105
timestamp 1586364061
transform 1 0 10764 0 -1 82144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_677
timestamp 1586364061
transform 1 0 12328 0 1 81056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_145_110
timestamp 1586364061
transform 1 0 11224 0 1 81056
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_145_123
timestamp 1586364061
transform 1 0 12420 0 1 81056
box -38 -48 222 592
use scs8hd_decap_8  FILLER_146_117
timestamp 1586364061
transform 1 0 11868 0 -1 82144
box -38 -48 774 592
use scs8hd_decap_3  PHY_291
timestamp 1586364061
transform -1 0 12880 0 1 81056
box -38 -48 314 592
use scs8hd_decap_3  PHY_293
timestamp 1586364061
transform -1 0 12880 0 -1 82144
box -38 -48 314 592
use scs8hd_decap_3  PHY_294
timestamp 1586364061
transform 1 0 1104 0 1 82144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_147_3
timestamp 1586364061
transform 1 0 1380 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_15
timestamp 1586364061
transform 1 0 2484 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_27
timestamp 1586364061
transform 1 0 3588 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_39
timestamp 1586364061
transform 1 0 4692 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_147_51
timestamp 1586364061
transform 1 0 5796 0 1 82144
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_680
timestamp 1586364061
transform 1 0 6716 0 1 82144
box -38 -48 130 592
use scs8hd_fill_2  FILLER_147_59
timestamp 1586364061
transform 1 0 6532 0 1 82144
box -38 -48 222 592
use scs8hd_decap_12  FILLER_147_62
timestamp 1586364061
transform 1 0 6808 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_74
timestamp 1586364061
transform 1 0 7912 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_86
timestamp 1586364061
transform 1 0 9016 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_98
timestamp 1586364061
transform 1 0 10120 0 1 82144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_681
timestamp 1586364061
transform 1 0 12328 0 1 82144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_147_110
timestamp 1586364061
transform 1 0 11224 0 1 82144
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_147_123
timestamp 1586364061
transform 1 0 12420 0 1 82144
box -38 -48 222 592
use scs8hd_decap_3  PHY_295
timestamp 1586364061
transform -1 0 12880 0 1 82144
box -38 -48 314 592
use scs8hd_decap_3  PHY_296
timestamp 1586364061
transform 1 0 1104 0 -1 83232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_148_3
timestamp 1586364061
transform 1 0 1380 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_15
timestamp 1586364061
transform 1 0 2484 0 -1 83232
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_682
timestamp 1586364061
transform 1 0 3956 0 -1 83232
box -38 -48 130 592
use scs8hd_decap_4  FILLER_148_27
timestamp 1586364061
transform 1 0 3588 0 -1 83232
box -38 -48 406 592
use scs8hd_decap_12  FILLER_148_32
timestamp 1586364061
transform 1 0 4048 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_44
timestamp 1586364061
transform 1 0 5152 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_56
timestamp 1586364061
transform 1 0 6256 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_68
timestamp 1586364061
transform 1 0 7360 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_80
timestamp 1586364061
transform 1 0 8464 0 -1 83232
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_683
timestamp 1586364061
transform 1 0 9568 0 -1 83232
box -38 -48 130 592
use scs8hd_decap_12  FILLER_148_93
timestamp 1586364061
transform 1 0 9660 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_105
timestamp 1586364061
transform 1 0 10764 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_148_117
timestamp 1586364061
transform 1 0 11868 0 -1 83232
box -38 -48 774 592
use scs8hd_decap_3  PHY_297
timestamp 1586364061
transform -1 0 12880 0 -1 83232
box -38 -48 314 592
use scs8hd_decap_3  PHY_298
timestamp 1586364061
transform 1 0 1104 0 1 83232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_149_3
timestamp 1586364061
transform 1 0 1380 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_15
timestamp 1586364061
transform 1 0 2484 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_27
timestamp 1586364061
transform 1 0 3588 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_39
timestamp 1586364061
transform 1 0 4692 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_149_51
timestamp 1586364061
transform 1 0 5796 0 1 83232
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_684
timestamp 1586364061
transform 1 0 6716 0 1 83232
box -38 -48 130 592
use scs8hd_fill_2  FILLER_149_59
timestamp 1586364061
transform 1 0 6532 0 1 83232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_149_62
timestamp 1586364061
transform 1 0 6808 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_74
timestamp 1586364061
transform 1 0 7912 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_86
timestamp 1586364061
transform 1 0 9016 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_98
timestamp 1586364061
transform 1 0 10120 0 1 83232
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_685
timestamp 1586364061
transform 1 0 12328 0 1 83232
box -38 -48 130 592
use scs8hd_decap_12  FILLER_149_110
timestamp 1586364061
transform 1 0 11224 0 1 83232
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_149_123
timestamp 1586364061
transform 1 0 12420 0 1 83232
box -38 -48 222 592
use scs8hd_decap_3  PHY_299
timestamp 1586364061
transform -1 0 12880 0 1 83232
box -38 -48 314 592
use scs8hd_decap_3  PHY_300
timestamp 1586364061
transform 1 0 1104 0 -1 84320
box -38 -48 314 592
use scs8hd_decap_12  FILLER_150_3
timestamp 1586364061
transform 1 0 1380 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_15
timestamp 1586364061
transform 1 0 2484 0 -1 84320
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_686
timestamp 1586364061
transform 1 0 3956 0 -1 84320
box -38 -48 130 592
use scs8hd_decap_4  FILLER_150_27
timestamp 1586364061
transform 1 0 3588 0 -1 84320
box -38 -48 406 592
use scs8hd_decap_12  FILLER_150_32
timestamp 1586364061
transform 1 0 4048 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_44
timestamp 1586364061
transform 1 0 5152 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_56
timestamp 1586364061
transform 1 0 6256 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_68
timestamp 1586364061
transform 1 0 7360 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_80
timestamp 1586364061
transform 1 0 8464 0 -1 84320
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_687
timestamp 1586364061
transform 1 0 9568 0 -1 84320
box -38 -48 130 592
use scs8hd_decap_12  FILLER_150_93
timestamp 1586364061
transform 1 0 9660 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_105
timestamp 1586364061
transform 1 0 10764 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_150_117
timestamp 1586364061
transform 1 0 11868 0 -1 84320
box -38 -48 774 592
use scs8hd_decap_3  PHY_301
timestamp 1586364061
transform -1 0 12880 0 -1 84320
box -38 -48 314 592
use scs8hd_decap_3  PHY_302
timestamp 1586364061
transform 1 0 1104 0 1 84320
box -38 -48 314 592
use scs8hd_decap_3  PHY_304
timestamp 1586364061
transform 1 0 1104 0 -1 85408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_151_3
timestamp 1586364061
transform 1 0 1380 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_151_15
timestamp 1586364061
transform 1 0 2484 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_3
timestamp 1586364061
transform 1 0 1380 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_15
timestamp 1586364061
transform 1 0 2484 0 -1 85408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_690
timestamp 1586364061
transform 1 0 3956 0 -1 85408
box -38 -48 130 592
use scs8hd_decap_12  FILLER_151_27
timestamp 1586364061
transform 1 0 3588 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_152_27
timestamp 1586364061
transform 1 0 3588 0 -1 85408
box -38 -48 406 592
use scs8hd_decap_12  FILLER_152_32
timestamp 1586364061
transform 1 0 4048 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_151_39
timestamp 1586364061
transform 1 0 4692 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_151_51
timestamp 1586364061
transform 1 0 5796 0 1 84320
box -38 -48 774 592
use scs8hd_decap_12  FILLER_152_44
timestamp 1586364061
transform 1 0 5152 0 -1 85408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_688
timestamp 1586364061
transform 1 0 6716 0 1 84320
box -38 -48 130 592
use scs8hd_fill_2  FILLER_151_59
timestamp 1586364061
transform 1 0 6532 0 1 84320
box -38 -48 222 592
use scs8hd_decap_12  FILLER_151_62
timestamp 1586364061
transform 1 0 6808 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_56
timestamp 1586364061
transform 1 0 6256 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_68
timestamp 1586364061
transform 1 0 7360 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_151_74
timestamp 1586364061
transform 1 0 7912 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_151_86
timestamp 1586364061
transform 1 0 9016 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_80
timestamp 1586364061
transform 1 0 8464 0 -1 85408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_691
timestamp 1586364061
transform 1 0 9568 0 -1 85408
box -38 -48 130 592
use scs8hd_decap_12  FILLER_151_98
timestamp 1586364061
transform 1 0 10120 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_93
timestamp 1586364061
transform 1 0 9660 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_152_105
timestamp 1586364061
transform 1 0 10764 0 -1 85408
box -38 -48 774 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 11500 0 -1 85408
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_689
timestamp 1586364061
transform 1 0 12328 0 1 84320
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 11500 0 1 84320
box -38 -48 222 592
use scs8hd_decap_3  FILLER_151_110
timestamp 1586364061
transform 1 0 11224 0 1 84320
box -38 -48 314 592
use scs8hd_decap_6  FILLER_151_115
timestamp 1586364061
transform 1 0 11684 0 1 84320
box -38 -48 590 592
use scs8hd_fill_1  FILLER_151_121
timestamp 1586364061
transform 1 0 12236 0 1 84320
box -38 -48 130 592
use scs8hd_fill_2  FILLER_151_123
timestamp 1586364061
transform 1 0 12420 0 1 84320
box -38 -48 222 592
use scs8hd_decap_8  FILLER_152_117
timestamp 1586364061
transform 1 0 11868 0 -1 85408
box -38 -48 774 592
use scs8hd_decap_3  PHY_303
timestamp 1586364061
transform -1 0 12880 0 1 84320
box -38 -48 314 592
use scs8hd_decap_3  PHY_305
timestamp 1586364061
transform -1 0 12880 0 -1 85408
box -38 -48 314 592
use scs8hd_decap_3  PHY_306
timestamp 1586364061
transform 1 0 1104 0 1 85408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_153_3
timestamp 1586364061
transform 1 0 1380 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_15
timestamp 1586364061
transform 1 0 2484 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_27
timestamp 1586364061
transform 1 0 3588 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_39
timestamp 1586364061
transform 1 0 4692 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_153_51
timestamp 1586364061
transform 1 0 5796 0 1 85408
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_692
timestamp 1586364061
transform 1 0 6716 0 1 85408
box -38 -48 130 592
use scs8hd_fill_2  FILLER_153_59
timestamp 1586364061
transform 1 0 6532 0 1 85408
box -38 -48 222 592
use scs8hd_decap_12  FILLER_153_62
timestamp 1586364061
transform 1 0 6808 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_74
timestamp 1586364061
transform 1 0 7912 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_86
timestamp 1586364061
transform 1 0 9016 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_98
timestamp 1586364061
transform 1 0 10120 0 1 85408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_693
timestamp 1586364061
transform 1 0 12328 0 1 85408
box -38 -48 130 592
use scs8hd_decap_12  FILLER_153_110
timestamp 1586364061
transform 1 0 11224 0 1 85408
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_153_123
timestamp 1586364061
transform 1 0 12420 0 1 85408
box -38 -48 222 592
use scs8hd_decap_3  PHY_307
timestamp 1586364061
transform -1 0 12880 0 1 85408
box -38 -48 314 592
use scs8hd_decap_3  PHY_308
timestamp 1586364061
transform 1 0 1104 0 -1 86496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_154_3
timestamp 1586364061
transform 1 0 1380 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_15
timestamp 1586364061
transform 1 0 2484 0 -1 86496
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_694
timestamp 1586364061
transform 1 0 3956 0 -1 86496
box -38 -48 130 592
use scs8hd_decap_4  FILLER_154_27
timestamp 1586364061
transform 1 0 3588 0 -1 86496
box -38 -48 406 592
use scs8hd_decap_12  FILLER_154_32
timestamp 1586364061
transform 1 0 4048 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_44
timestamp 1586364061
transform 1 0 5152 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_56
timestamp 1586364061
transform 1 0 6256 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_68
timestamp 1586364061
transform 1 0 7360 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_80
timestamp 1586364061
transform 1 0 8464 0 -1 86496
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_695
timestamp 1586364061
transform 1 0 9568 0 -1 86496
box -38 -48 130 592
use scs8hd_decap_12  FILLER_154_93
timestamp 1586364061
transform 1 0 9660 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_105
timestamp 1586364061
transform 1 0 10764 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_154_117
timestamp 1586364061
transform 1 0 11868 0 -1 86496
box -38 -48 774 592
use scs8hd_decap_3  PHY_309
timestamp 1586364061
transform -1 0 12880 0 -1 86496
box -38 -48 314 592
use scs8hd_decap_3  PHY_310
timestamp 1586364061
transform 1 0 1104 0 1 86496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_155_3
timestamp 1586364061
transform 1 0 1380 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_15
timestamp 1586364061
transform 1 0 2484 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_27
timestamp 1586364061
transform 1 0 3588 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_39
timestamp 1586364061
transform 1 0 4692 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_155_51
timestamp 1586364061
transform 1 0 5796 0 1 86496
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_696
timestamp 1586364061
transform 1 0 6716 0 1 86496
box -38 -48 130 592
use scs8hd_fill_2  FILLER_155_59
timestamp 1586364061
transform 1 0 6532 0 1 86496
box -38 -48 222 592
use scs8hd_decap_12  FILLER_155_62
timestamp 1586364061
transform 1 0 6808 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_74
timestamp 1586364061
transform 1 0 7912 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_86
timestamp 1586364061
transform 1 0 9016 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_98
timestamp 1586364061
transform 1 0 10120 0 1 86496
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_697
timestamp 1586364061
transform 1 0 12328 0 1 86496
box -38 -48 130 592
use scs8hd_decap_12  FILLER_155_110
timestamp 1586364061
transform 1 0 11224 0 1 86496
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_155_123
timestamp 1586364061
transform 1 0 12420 0 1 86496
box -38 -48 222 592
use scs8hd_decap_3  PHY_311
timestamp 1586364061
transform -1 0 12880 0 1 86496
box -38 -48 314 592
use scs8hd_decap_3  PHY_312
timestamp 1586364061
transform 1 0 1104 0 -1 87584
box -38 -48 314 592
use scs8hd_decap_12  FILLER_156_3
timestamp 1586364061
transform 1 0 1380 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_15
timestamp 1586364061
transform 1 0 2484 0 -1 87584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_698
timestamp 1586364061
transform 1 0 3956 0 -1 87584
box -38 -48 130 592
use scs8hd_decap_4  FILLER_156_27
timestamp 1586364061
transform 1 0 3588 0 -1 87584
box -38 -48 406 592
use scs8hd_decap_12  FILLER_156_32
timestamp 1586364061
transform 1 0 4048 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_44
timestamp 1586364061
transform 1 0 5152 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_56
timestamp 1586364061
transform 1 0 6256 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_68
timestamp 1586364061
transform 1 0 7360 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_80
timestamp 1586364061
transform 1 0 8464 0 -1 87584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_699
timestamp 1586364061
transform 1 0 9568 0 -1 87584
box -38 -48 130 592
use scs8hd_decap_12  FILLER_156_93
timestamp 1586364061
transform 1 0 9660 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_105
timestamp 1586364061
transform 1 0 10764 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_156_117
timestamp 1586364061
transform 1 0 11868 0 -1 87584
box -38 -48 774 592
use scs8hd_decap_3  PHY_313
timestamp 1586364061
transform -1 0 12880 0 -1 87584
box -38 -48 314 592
use scs8hd_decap_3  PHY_314
timestamp 1586364061
transform 1 0 1104 0 1 87584
box -38 -48 314 592
use scs8hd_decap_12  FILLER_157_3
timestamp 1586364061
transform 1 0 1380 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_15
timestamp 1586364061
transform 1 0 2484 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_27
timestamp 1586364061
transform 1 0 3588 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_39
timestamp 1586364061
transform 1 0 4692 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_157_51
timestamp 1586364061
transform 1 0 5796 0 1 87584
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_700
timestamp 1586364061
transform 1 0 6716 0 1 87584
box -38 -48 130 592
use scs8hd_fill_2  FILLER_157_59
timestamp 1586364061
transform 1 0 6532 0 1 87584
box -38 -48 222 592
use scs8hd_decap_12  FILLER_157_62
timestamp 1586364061
transform 1 0 6808 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_74
timestamp 1586364061
transform 1 0 7912 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_86
timestamp 1586364061
transform 1 0 9016 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_98
timestamp 1586364061
transform 1 0 10120 0 1 87584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_701
timestamp 1586364061
transform 1 0 12328 0 1 87584
box -38 -48 130 592
use scs8hd_decap_12  FILLER_157_110
timestamp 1586364061
transform 1 0 11224 0 1 87584
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_157_123
timestamp 1586364061
transform 1 0 12420 0 1 87584
box -38 -48 222 592
use scs8hd_decap_3  PHY_315
timestamp 1586364061
transform -1 0 12880 0 1 87584
box -38 -48 314 592
use scs8hd_decap_3  PHY_316
timestamp 1586364061
transform 1 0 1104 0 -1 88672
box -38 -48 314 592
use scs8hd_decap_3  PHY_318
timestamp 1586364061
transform 1 0 1104 0 1 88672
box -38 -48 314 592
use scs8hd_decap_12  FILLER_158_3
timestamp 1586364061
transform 1 0 1380 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_15
timestamp 1586364061
transform 1 0 2484 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_3
timestamp 1586364061
transform 1 0 1380 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_15
timestamp 1586364061
transform 1 0 2484 0 1 88672
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_702
timestamp 1586364061
transform 1 0 3956 0 -1 88672
box -38 -48 130 592
use scs8hd_decap_4  FILLER_158_27
timestamp 1586364061
transform 1 0 3588 0 -1 88672
box -38 -48 406 592
use scs8hd_decap_12  FILLER_158_32
timestamp 1586364061
transform 1 0 4048 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_27
timestamp 1586364061
transform 1 0 3588 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_44
timestamp 1586364061
transform 1 0 5152 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_39
timestamp 1586364061
transform 1 0 4692 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_159_51
timestamp 1586364061
transform 1 0 5796 0 1 88672
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_704
timestamp 1586364061
transform 1 0 6716 0 1 88672
box -38 -48 130 592
use scs8hd_decap_12  FILLER_158_56
timestamp 1586364061
transform 1 0 6256 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_68
timestamp 1586364061
transform 1 0 7360 0 -1 88672
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_159_59
timestamp 1586364061
transform 1 0 6532 0 1 88672
box -38 -48 222 592
use scs8hd_decap_12  FILLER_159_62
timestamp 1586364061
transform 1 0 6808 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_80
timestamp 1586364061
transform 1 0 8464 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_74
timestamp 1586364061
transform 1 0 7912 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_86
timestamp 1586364061
transform 1 0 9016 0 1 88672
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_703
timestamp 1586364061
transform 1 0 9568 0 -1 88672
box -38 -48 130 592
use scs8hd_decap_12  FILLER_158_93
timestamp 1586364061
transform 1 0 9660 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_105
timestamp 1586364061
transform 1 0 10764 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_98
timestamp 1586364061
transform 1 0 10120 0 1 88672
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_705
timestamp 1586364061
transform 1 0 12328 0 1 88672
box -38 -48 130 592
use scs8hd_decap_8  FILLER_158_117
timestamp 1586364061
transform 1 0 11868 0 -1 88672
box -38 -48 774 592
use scs8hd_decap_12  FILLER_159_110
timestamp 1586364061
transform 1 0 11224 0 1 88672
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_159_123
timestamp 1586364061
transform 1 0 12420 0 1 88672
box -38 -48 222 592
use scs8hd_decap_3  PHY_317
timestamp 1586364061
transform -1 0 12880 0 -1 88672
box -38 -48 314 592
use scs8hd_decap_3  PHY_319
timestamp 1586364061
transform -1 0 12880 0 1 88672
box -38 -48 314 592
use scs8hd_decap_3  PHY_320
timestamp 1586364061
transform 1 0 1104 0 -1 89760
box -38 -48 314 592
use scs8hd_decap_12  FILLER_160_3
timestamp 1586364061
transform 1 0 1380 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_15
timestamp 1586364061
transform 1 0 2484 0 -1 89760
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_706
timestamp 1586364061
transform 1 0 3956 0 -1 89760
box -38 -48 130 592
use scs8hd_decap_4  FILLER_160_27
timestamp 1586364061
transform 1 0 3588 0 -1 89760
box -38 -48 406 592
use scs8hd_decap_12  FILLER_160_32
timestamp 1586364061
transform 1 0 4048 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_44
timestamp 1586364061
transform 1 0 5152 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_56
timestamp 1586364061
transform 1 0 6256 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_68
timestamp 1586364061
transform 1 0 7360 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_80
timestamp 1586364061
transform 1 0 8464 0 -1 89760
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_707
timestamp 1586364061
transform 1 0 9568 0 -1 89760
box -38 -48 130 592
use scs8hd_decap_12  FILLER_160_93
timestamp 1586364061
transform 1 0 9660 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_105
timestamp 1586364061
transform 1 0 10764 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_160_117
timestamp 1586364061
transform 1 0 11868 0 -1 89760
box -38 -48 774 592
use scs8hd_decap_3  PHY_321
timestamp 1586364061
transform -1 0 12880 0 -1 89760
box -38 -48 314 592
use scs8hd_decap_3  PHY_322
timestamp 1586364061
transform 1 0 1104 0 1 89760
box -38 -48 314 592
use scs8hd_decap_12  FILLER_161_3
timestamp 1586364061
transform 1 0 1380 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_15
timestamp 1586364061
transform 1 0 2484 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_27
timestamp 1586364061
transform 1 0 3588 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_39
timestamp 1586364061
transform 1 0 4692 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_161_51
timestamp 1586364061
transform 1 0 5796 0 1 89760
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_708
timestamp 1586364061
transform 1 0 6716 0 1 89760
box -38 -48 130 592
use scs8hd_fill_2  FILLER_161_59
timestamp 1586364061
transform 1 0 6532 0 1 89760
box -38 -48 222 592
use scs8hd_decap_12  FILLER_161_62
timestamp 1586364061
transform 1 0 6808 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_74
timestamp 1586364061
transform 1 0 7912 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_86
timestamp 1586364061
transform 1 0 9016 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_98
timestamp 1586364061
transform 1 0 10120 0 1 89760
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_709
timestamp 1586364061
transform 1 0 12328 0 1 89760
box -38 -48 130 592
use scs8hd_decap_12  FILLER_161_110
timestamp 1586364061
transform 1 0 11224 0 1 89760
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_161_123
timestamp 1586364061
transform 1 0 12420 0 1 89760
box -38 -48 222 592
use scs8hd_decap_3  PHY_323
timestamp 1586364061
transform -1 0 12880 0 1 89760
box -38 -48 314 592
use scs8hd_decap_3  PHY_324
timestamp 1586364061
transform 1 0 1104 0 -1 90848
box -38 -48 314 592
use scs8hd_decap_12  FILLER_162_3
timestamp 1586364061
transform 1 0 1380 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_15
timestamp 1586364061
transform 1 0 2484 0 -1 90848
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_710
timestamp 1586364061
transform 1 0 3956 0 -1 90848
box -38 -48 130 592
use scs8hd_decap_4  FILLER_162_27
timestamp 1586364061
transform 1 0 3588 0 -1 90848
box -38 -48 406 592
use scs8hd_decap_12  FILLER_162_32
timestamp 1586364061
transform 1 0 4048 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_44
timestamp 1586364061
transform 1 0 5152 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_56
timestamp 1586364061
transform 1 0 6256 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_68
timestamp 1586364061
transform 1 0 7360 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_80
timestamp 1586364061
transform 1 0 8464 0 -1 90848
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_711
timestamp 1586364061
transform 1 0 9568 0 -1 90848
box -38 -48 130 592
use scs8hd_decap_12  FILLER_162_93
timestamp 1586364061
transform 1 0 9660 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_105
timestamp 1586364061
transform 1 0 10764 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_162_117
timestamp 1586364061
transform 1 0 11868 0 -1 90848
box -38 -48 774 592
use scs8hd_decap_3  PHY_325
timestamp 1586364061
transform -1 0 12880 0 -1 90848
box -38 -48 314 592
use scs8hd_decap_3  PHY_326
timestamp 1586364061
transform 1 0 1104 0 1 90848
box -38 -48 314 592
use scs8hd_decap_12  FILLER_163_3
timestamp 1586364061
transform 1 0 1380 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_15
timestamp 1586364061
transform 1 0 2484 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_27
timestamp 1586364061
transform 1 0 3588 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_39
timestamp 1586364061
transform 1 0 4692 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_163_51
timestamp 1586364061
transform 1 0 5796 0 1 90848
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_712
timestamp 1586364061
transform 1 0 6716 0 1 90848
box -38 -48 130 592
use scs8hd_fill_2  FILLER_163_59
timestamp 1586364061
transform 1 0 6532 0 1 90848
box -38 -48 222 592
use scs8hd_decap_12  FILLER_163_62
timestamp 1586364061
transform 1 0 6808 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_74
timestamp 1586364061
transform 1 0 7912 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_86
timestamp 1586364061
transform 1 0 9016 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_98
timestamp 1586364061
transform 1 0 10120 0 1 90848
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_713
timestamp 1586364061
transform 1 0 12328 0 1 90848
box -38 -48 130 592
use scs8hd_decap_12  FILLER_163_110
timestamp 1586364061
transform 1 0 11224 0 1 90848
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_163_123
timestamp 1586364061
transform 1 0 12420 0 1 90848
box -38 -48 222 592
use scs8hd_decap_3  PHY_327
timestamp 1586364061
transform -1 0 12880 0 1 90848
box -38 -48 314 592
use scs8hd_decap_3  PHY_328
timestamp 1586364061
transform 1 0 1104 0 -1 91936
box -38 -48 314 592
use scs8hd_decap_12  FILLER_164_3
timestamp 1586364061
transform 1 0 1380 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_15
timestamp 1586364061
transform 1 0 2484 0 -1 91936
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_714
timestamp 1586364061
transform 1 0 3956 0 -1 91936
box -38 -48 130 592
use scs8hd_decap_4  FILLER_164_27
timestamp 1586364061
transform 1 0 3588 0 -1 91936
box -38 -48 406 592
use scs8hd_decap_12  FILLER_164_32
timestamp 1586364061
transform 1 0 4048 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_44
timestamp 1586364061
transform 1 0 5152 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_56
timestamp 1586364061
transform 1 0 6256 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_68
timestamp 1586364061
transform 1 0 7360 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_80
timestamp 1586364061
transform 1 0 8464 0 -1 91936
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_715
timestamp 1586364061
transform 1 0 9568 0 -1 91936
box -38 -48 130 592
use scs8hd_decap_12  FILLER_164_93
timestamp 1586364061
transform 1 0 9660 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_105
timestamp 1586364061
transform 1 0 10764 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_164_117
timestamp 1586364061
transform 1 0 11868 0 -1 91936
box -38 -48 774 592
use scs8hd_decap_3  PHY_329
timestamp 1586364061
transform -1 0 12880 0 -1 91936
box -38 -48 314 592
use scs8hd_decap_3  PHY_330
timestamp 1586364061
transform 1 0 1104 0 1 91936
box -38 -48 314 592
use scs8hd_decap_3  PHY_332
timestamp 1586364061
transform 1 0 1104 0 -1 93024
box -38 -48 314 592
use scs8hd_decap_12  FILLER_165_3
timestamp 1586364061
transform 1 0 1380 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_165_15
timestamp 1586364061
transform 1 0 2484 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_3
timestamp 1586364061
transform 1 0 1380 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_15
timestamp 1586364061
transform 1 0 2484 0 -1 93024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_718
timestamp 1586364061
transform 1 0 3956 0 -1 93024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_165_27
timestamp 1586364061
transform 1 0 3588 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_166_27
timestamp 1586364061
transform 1 0 3588 0 -1 93024
box -38 -48 406 592
use scs8hd_decap_12  FILLER_166_32
timestamp 1586364061
transform 1 0 4048 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_165_39
timestamp 1586364061
transform 1 0 4692 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_165_51
timestamp 1586364061
transform 1 0 5796 0 1 91936
box -38 -48 774 592
use scs8hd_decap_12  FILLER_166_44
timestamp 1586364061
transform 1 0 5152 0 -1 93024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_716
timestamp 1586364061
transform 1 0 6716 0 1 91936
box -38 -48 130 592
use scs8hd_fill_2  FILLER_165_59
timestamp 1586364061
transform 1 0 6532 0 1 91936
box -38 -48 222 592
use scs8hd_decap_12  FILLER_165_62
timestamp 1586364061
transform 1 0 6808 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_56
timestamp 1586364061
transform 1 0 6256 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_68
timestamp 1586364061
transform 1 0 7360 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_165_74
timestamp 1586364061
transform 1 0 7912 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_165_86
timestamp 1586364061
transform 1 0 9016 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_80
timestamp 1586364061
transform 1 0 8464 0 -1 93024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_719
timestamp 1586364061
transform 1 0 9568 0 -1 93024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_165_98
timestamp 1586364061
transform 1 0 10120 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_93
timestamp 1586364061
transform 1 0 9660 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_105
timestamp 1586364061
transform 1 0 10764 0 -1 93024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_717
timestamp 1586364061
transform 1 0 12328 0 1 91936
box -38 -48 130 592
use scs8hd_decap_12  FILLER_165_110
timestamp 1586364061
transform 1 0 11224 0 1 91936
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_165_123
timestamp 1586364061
transform 1 0 12420 0 1 91936
box -38 -48 222 592
use scs8hd_decap_8  FILLER_166_117
timestamp 1586364061
transform 1 0 11868 0 -1 93024
box -38 -48 774 592
use scs8hd_decap_3  PHY_331
timestamp 1586364061
transform -1 0 12880 0 1 91936
box -38 -48 314 592
use scs8hd_decap_3  PHY_333
timestamp 1586364061
transform -1 0 12880 0 -1 93024
box -38 -48 314 592
use scs8hd_decap_3  PHY_334
timestamp 1586364061
transform 1 0 1104 0 1 93024
box -38 -48 314 592
use scs8hd_decap_12  FILLER_167_3
timestamp 1586364061
transform 1 0 1380 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_15
timestamp 1586364061
transform 1 0 2484 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_27
timestamp 1586364061
transform 1 0 3588 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_39
timestamp 1586364061
transform 1 0 4692 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_167_51
timestamp 1586364061
transform 1 0 5796 0 1 93024
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_720
timestamp 1586364061
transform 1 0 6716 0 1 93024
box -38 -48 130 592
use scs8hd_fill_2  FILLER_167_59
timestamp 1586364061
transform 1 0 6532 0 1 93024
box -38 -48 222 592
use scs8hd_decap_12  FILLER_167_62
timestamp 1586364061
transform 1 0 6808 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_74
timestamp 1586364061
transform 1 0 7912 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_86
timestamp 1586364061
transform 1 0 9016 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_98
timestamp 1586364061
transform 1 0 10120 0 1 93024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_721
timestamp 1586364061
transform 1 0 12328 0 1 93024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_167_110
timestamp 1586364061
transform 1 0 11224 0 1 93024
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_167_123
timestamp 1586364061
transform 1 0 12420 0 1 93024
box -38 -48 222 592
use scs8hd_decap_3  PHY_335
timestamp 1586364061
transform -1 0 12880 0 1 93024
box -38 -48 314 592
use scs8hd_decap_3  PHY_336
timestamp 1586364061
transform 1 0 1104 0 -1 94112
box -38 -48 314 592
use scs8hd_decap_12  FILLER_168_3
timestamp 1586364061
transform 1 0 1380 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_15
timestamp 1586364061
transform 1 0 2484 0 -1 94112
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_722
timestamp 1586364061
transform 1 0 3956 0 -1 94112
box -38 -48 130 592
use scs8hd_decap_4  FILLER_168_27
timestamp 1586364061
transform 1 0 3588 0 -1 94112
box -38 -48 406 592
use scs8hd_decap_12  FILLER_168_32
timestamp 1586364061
transform 1 0 4048 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_44
timestamp 1586364061
transform 1 0 5152 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_56
timestamp 1586364061
transform 1 0 6256 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_68
timestamp 1586364061
transform 1 0 7360 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_80
timestamp 1586364061
transform 1 0 8464 0 -1 94112
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_723
timestamp 1586364061
transform 1 0 9568 0 -1 94112
box -38 -48 130 592
use scs8hd_decap_12  FILLER_168_93
timestamp 1586364061
transform 1 0 9660 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_105
timestamp 1586364061
transform 1 0 10764 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_168_117
timestamp 1586364061
transform 1 0 11868 0 -1 94112
box -38 -48 774 592
use scs8hd_decap_3  PHY_337
timestamp 1586364061
transform -1 0 12880 0 -1 94112
box -38 -48 314 592
use scs8hd_decap_3  PHY_338
timestamp 1586364061
transform 1 0 1104 0 1 94112
box -38 -48 314 592
use scs8hd_decap_12  FILLER_169_3
timestamp 1586364061
transform 1 0 1380 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_15
timestamp 1586364061
transform 1 0 2484 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_27
timestamp 1586364061
transform 1 0 3588 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_39
timestamp 1586364061
transform 1 0 4692 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_169_51
timestamp 1586364061
transform 1 0 5796 0 1 94112
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_724
timestamp 1586364061
transform 1 0 6716 0 1 94112
box -38 -48 130 592
use scs8hd_fill_2  FILLER_169_59
timestamp 1586364061
transform 1 0 6532 0 1 94112
box -38 -48 222 592
use scs8hd_decap_12  FILLER_169_62
timestamp 1586364061
transform 1 0 6808 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_74
timestamp 1586364061
transform 1 0 7912 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_86
timestamp 1586364061
transform 1 0 9016 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_169_98
timestamp 1586364061
transform 1 0 10120 0 1 94112
box -38 -48 774 592
use scs8hd_decap_3  FILLER_169_106
timestamp 1586364061
transform 1 0 10856 0 1 94112
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_725
timestamp 1586364061
transform 1 0 12328 0 1 94112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 11132 0 1 94112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 11500 0 1 94112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_169_111
timestamp 1586364061
transform 1 0 11316 0 1 94112
box -38 -48 222 592
use scs8hd_decap_6  FILLER_169_115
timestamp 1586364061
transform 1 0 11684 0 1 94112
box -38 -48 590 592
use scs8hd_fill_1  FILLER_169_121
timestamp 1586364061
transform 1 0 12236 0 1 94112
box -38 -48 130 592
use scs8hd_fill_2  FILLER_169_123
timestamp 1586364061
transform 1 0 12420 0 1 94112
box -38 -48 222 592
use scs8hd_decap_3  PHY_339
timestamp 1586364061
transform -1 0 12880 0 1 94112
box -38 -48 314 592
use scs8hd_decap_3  PHY_340
timestamp 1586364061
transform 1 0 1104 0 -1 95200
box -38 -48 314 592
use scs8hd_decap_12  FILLER_170_3
timestamp 1586364061
transform 1 0 1380 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_15
timestamp 1586364061
transform 1 0 2484 0 -1 95200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_726
timestamp 1586364061
transform 1 0 3956 0 -1 95200
box -38 -48 130 592
use scs8hd_decap_4  FILLER_170_27
timestamp 1586364061
transform 1 0 3588 0 -1 95200
box -38 -48 406 592
use scs8hd_decap_12  FILLER_170_32
timestamp 1586364061
transform 1 0 4048 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_44
timestamp 1586364061
transform 1 0 5152 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_56
timestamp 1586364061
transform 1 0 6256 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_68
timestamp 1586364061
transform 1 0 7360 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_80
timestamp 1586364061
transform 1 0 8464 0 -1 95200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_727
timestamp 1586364061
transform 1 0 9568 0 -1 95200
box -38 -48 130 592
use scs8hd_decap_12  FILLER_170_93
timestamp 1586364061
transform 1 0 9660 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_170_105
timestamp 1586364061
transform 1 0 10764 0 -1 95200
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 11132 0 -1 95200
box -38 -48 774 592
use scs8hd_decap_8  FILLER_170_117
timestamp 1586364061
transform 1 0 11868 0 -1 95200
box -38 -48 774 592
use scs8hd_decap_3  PHY_341
timestamp 1586364061
transform -1 0 12880 0 -1 95200
box -38 -48 314 592
use scs8hd_decap_3  PHY_342
timestamp 1586364061
transform 1 0 1104 0 1 95200
box -38 -48 314 592
use scs8hd_decap_3  PHY_344
timestamp 1586364061
transform 1 0 1104 0 -1 96288
box -38 -48 314 592
use scs8hd_decap_12  FILLER_171_3
timestamp 1586364061
transform 1 0 1380 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_171_15
timestamp 1586364061
transform 1 0 2484 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_3
timestamp 1586364061
transform 1 0 1380 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_15
timestamp 1586364061
transform 1 0 2484 0 -1 96288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_730
timestamp 1586364061
transform 1 0 3956 0 -1 96288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_171_27
timestamp 1586364061
transform 1 0 3588 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_172_27
timestamp 1586364061
transform 1 0 3588 0 -1 96288
box -38 -48 406 592
use scs8hd_decap_12  FILLER_172_32
timestamp 1586364061
transform 1 0 4048 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_171_39
timestamp 1586364061
transform 1 0 4692 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_171_51
timestamp 1586364061
transform 1 0 5796 0 1 95200
box -38 -48 774 592
use scs8hd_decap_12  FILLER_172_44
timestamp 1586364061
transform 1 0 5152 0 -1 96288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_728
timestamp 1586364061
transform 1 0 6716 0 1 95200
box -38 -48 130 592
use scs8hd_fill_2  FILLER_171_59
timestamp 1586364061
transform 1 0 6532 0 1 95200
box -38 -48 222 592
use scs8hd_decap_12  FILLER_171_62
timestamp 1586364061
transform 1 0 6808 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_56
timestamp 1586364061
transform 1 0 6256 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_68
timestamp 1586364061
transform 1 0 7360 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_171_74
timestamp 1586364061
transform 1 0 7912 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_171_86
timestamp 1586364061
transform 1 0 9016 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_80
timestamp 1586364061
transform 1 0 8464 0 -1 96288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_731
timestamp 1586364061
transform 1 0 9568 0 -1 96288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_171_98
timestamp 1586364061
transform 1 0 10120 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_93
timestamp 1586364061
transform 1 0 9660 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_105
timestamp 1586364061
transform 1 0 10764 0 -1 96288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_729
timestamp 1586364061
transform 1 0 12328 0 1 95200
box -38 -48 130 592
use scs8hd_decap_12  FILLER_171_110
timestamp 1586364061
transform 1 0 11224 0 1 95200
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_171_123
timestamp 1586364061
transform 1 0 12420 0 1 95200
box -38 -48 222 592
use scs8hd_decap_8  FILLER_172_117
timestamp 1586364061
transform 1 0 11868 0 -1 96288
box -38 -48 774 592
use scs8hd_decap_3  PHY_343
timestamp 1586364061
transform -1 0 12880 0 1 95200
box -38 -48 314 592
use scs8hd_decap_3  PHY_345
timestamp 1586364061
transform -1 0 12880 0 -1 96288
box -38 -48 314 592
use scs8hd_decap_3  PHY_346
timestamp 1586364061
transform 1 0 1104 0 1 96288
box -38 -48 314 592
use scs8hd_decap_12  FILLER_173_3
timestamp 1586364061
transform 1 0 1380 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_15
timestamp 1586364061
transform 1 0 2484 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_27
timestamp 1586364061
transform 1 0 3588 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_39
timestamp 1586364061
transform 1 0 4692 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_173_51
timestamp 1586364061
transform 1 0 5796 0 1 96288
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_732
timestamp 1586364061
transform 1 0 6716 0 1 96288
box -38 -48 130 592
use scs8hd_fill_2  FILLER_173_59
timestamp 1586364061
transform 1 0 6532 0 1 96288
box -38 -48 222 592
use scs8hd_decap_12  FILLER_173_62
timestamp 1586364061
transform 1 0 6808 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_74
timestamp 1586364061
transform 1 0 7912 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_86
timestamp 1586364061
transform 1 0 9016 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_98
timestamp 1586364061
transform 1 0 10120 0 1 96288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_733
timestamp 1586364061
transform 1 0 12328 0 1 96288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_173_110
timestamp 1586364061
transform 1 0 11224 0 1 96288
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_173_123
timestamp 1586364061
transform 1 0 12420 0 1 96288
box -38 -48 222 592
use scs8hd_decap_3  PHY_347
timestamp 1586364061
transform -1 0 12880 0 1 96288
box -38 -48 314 592
use scs8hd_decap_3  PHY_348
timestamp 1586364061
transform 1 0 1104 0 -1 97376
box -38 -48 314 592
use scs8hd_decap_12  FILLER_174_3
timestamp 1586364061
transform 1 0 1380 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_15
timestamp 1586364061
transform 1 0 2484 0 -1 97376
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_734
timestamp 1586364061
transform 1 0 3956 0 -1 97376
box -38 -48 130 592
use scs8hd_decap_4  FILLER_174_27
timestamp 1586364061
transform 1 0 3588 0 -1 97376
box -38 -48 406 592
use scs8hd_decap_12  FILLER_174_32
timestamp 1586364061
transform 1 0 4048 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_44
timestamp 1586364061
transform 1 0 5152 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_56
timestamp 1586364061
transform 1 0 6256 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_68
timestamp 1586364061
transform 1 0 7360 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_80
timestamp 1586364061
transform 1 0 8464 0 -1 97376
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_735
timestamp 1586364061
transform 1 0 9568 0 -1 97376
box -38 -48 130 592
use scs8hd_decap_12  FILLER_174_93
timestamp 1586364061
transform 1 0 9660 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_105
timestamp 1586364061
transform 1 0 10764 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_174_117
timestamp 1586364061
transform 1 0 11868 0 -1 97376
box -38 -48 774 592
use scs8hd_decap_3  PHY_349
timestamp 1586364061
transform -1 0 12880 0 -1 97376
box -38 -48 314 592
use scs8hd_decap_3  PHY_350
timestamp 1586364061
transform 1 0 1104 0 1 97376
box -38 -48 314 592
use scs8hd_decap_12  FILLER_175_3
timestamp 1586364061
transform 1 0 1380 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_15
timestamp 1586364061
transform 1 0 2484 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_27
timestamp 1586364061
transform 1 0 3588 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_39
timestamp 1586364061
transform 1 0 4692 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_175_51
timestamp 1586364061
transform 1 0 5796 0 1 97376
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_736
timestamp 1586364061
transform 1 0 6716 0 1 97376
box -38 -48 130 592
use scs8hd_fill_2  FILLER_175_59
timestamp 1586364061
transform 1 0 6532 0 1 97376
box -38 -48 222 592
use scs8hd_decap_12  FILLER_175_62
timestamp 1586364061
transform 1 0 6808 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_74
timestamp 1586364061
transform 1 0 7912 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_86
timestamp 1586364061
transform 1 0 9016 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_98
timestamp 1586364061
transform 1 0 10120 0 1 97376
box -38 -48 1142 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 11224 0 1 97376
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_737
timestamp 1586364061
transform 1 0 12328 0 1 97376
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 11776 0 1 97376
box -38 -48 222 592
use scs8hd_fill_2  FILLER_175_114
timestamp 1586364061
transform 1 0 11592 0 1 97376
box -38 -48 222 592
use scs8hd_decap_4  FILLER_175_118
timestamp 1586364061
transform 1 0 11960 0 1 97376
box -38 -48 406 592
use scs8hd_fill_2  FILLER_175_123
timestamp 1586364061
transform 1 0 12420 0 1 97376
box -38 -48 222 592
use scs8hd_decap_3  PHY_351
timestamp 1586364061
transform -1 0 12880 0 1 97376
box -38 -48 314 592
use scs8hd_decap_3  PHY_352
timestamp 1586364061
transform 1 0 1104 0 -1 98464
box -38 -48 314 592
use scs8hd_decap_12  FILLER_176_3
timestamp 1586364061
transform 1 0 1380 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_15
timestamp 1586364061
transform 1 0 2484 0 -1 98464
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_738
timestamp 1586364061
transform 1 0 3956 0 -1 98464
box -38 -48 130 592
use scs8hd_decap_4  FILLER_176_27
timestamp 1586364061
transform 1 0 3588 0 -1 98464
box -38 -48 406 592
use scs8hd_decap_12  FILLER_176_32
timestamp 1586364061
transform 1 0 4048 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_44
timestamp 1586364061
transform 1 0 5152 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_56
timestamp 1586364061
transform 1 0 6256 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_68
timestamp 1586364061
transform 1 0 7360 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_80
timestamp 1586364061
transform 1 0 8464 0 -1 98464
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_739
timestamp 1586364061
transform 1 0 9568 0 -1 98464
box -38 -48 130 592
use scs8hd_decap_12  FILLER_176_93
timestamp 1586364061
transform 1 0 9660 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_105
timestamp 1586364061
transform 1 0 10764 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_176_117
timestamp 1586364061
transform 1 0 11868 0 -1 98464
box -38 -48 774 592
use scs8hd_decap_3  PHY_353
timestamp 1586364061
transform -1 0 12880 0 -1 98464
box -38 -48 314 592
use scs8hd_decap_3  PHY_354
timestamp 1586364061
transform 1 0 1104 0 1 98464
box -38 -48 314 592
use scs8hd_decap_12  FILLER_177_3
timestamp 1586364061
transform 1 0 1380 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_15
timestamp 1586364061
transform 1 0 2484 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_27
timestamp 1586364061
transform 1 0 3588 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_39
timestamp 1586364061
transform 1 0 4692 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_177_51
timestamp 1586364061
transform 1 0 5796 0 1 98464
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_740
timestamp 1586364061
transform 1 0 6716 0 1 98464
box -38 -48 130 592
use scs8hd_fill_2  FILLER_177_59
timestamp 1586364061
transform 1 0 6532 0 1 98464
box -38 -48 222 592
use scs8hd_decap_12  FILLER_177_62
timestamp 1586364061
transform 1 0 6808 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_74
timestamp 1586364061
transform 1 0 7912 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_86
timestamp 1586364061
transform 1 0 9016 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_98
timestamp 1586364061
transform 1 0 10120 0 1 98464
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_741
timestamp 1586364061
transform 1 0 12328 0 1 98464
box -38 -48 130 592
use scs8hd_decap_12  FILLER_177_110
timestamp 1586364061
transform 1 0 11224 0 1 98464
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_177_123
timestamp 1586364061
transform 1 0 12420 0 1 98464
box -38 -48 222 592
use scs8hd_decap_3  PHY_355
timestamp 1586364061
transform -1 0 12880 0 1 98464
box -38 -48 314 592
use scs8hd_decap_3  PHY_356
timestamp 1586364061
transform 1 0 1104 0 -1 99552
box -38 -48 314 592
use scs8hd_decap_3  PHY_358
timestamp 1586364061
transform 1 0 1104 0 1 99552
box -38 -48 314 592
use scs8hd_decap_12  FILLER_178_3
timestamp 1586364061
transform 1 0 1380 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_15
timestamp 1586364061
transform 1 0 2484 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_3
timestamp 1586364061
transform 1 0 1380 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_15
timestamp 1586364061
transform 1 0 2484 0 1 99552
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_742
timestamp 1586364061
transform 1 0 3956 0 -1 99552
box -38 -48 130 592
use scs8hd_decap_4  FILLER_178_27
timestamp 1586364061
transform 1 0 3588 0 -1 99552
box -38 -48 406 592
use scs8hd_decap_12  FILLER_178_32
timestamp 1586364061
transform 1 0 4048 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_27
timestamp 1586364061
transform 1 0 3588 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_44
timestamp 1586364061
transform 1 0 5152 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_39
timestamp 1586364061
transform 1 0 4692 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_179_51
timestamp 1586364061
transform 1 0 5796 0 1 99552
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_744
timestamp 1586364061
transform 1 0 6716 0 1 99552
box -38 -48 130 592
use scs8hd_decap_12  FILLER_178_56
timestamp 1586364061
transform 1 0 6256 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_68
timestamp 1586364061
transform 1 0 7360 0 -1 99552
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_179_59
timestamp 1586364061
transform 1 0 6532 0 1 99552
box -38 -48 222 592
use scs8hd_decap_12  FILLER_179_62
timestamp 1586364061
transform 1 0 6808 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_80
timestamp 1586364061
transform 1 0 8464 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_74
timestamp 1586364061
transform 1 0 7912 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_86
timestamp 1586364061
transform 1 0 9016 0 1 99552
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_743
timestamp 1586364061
transform 1 0 9568 0 -1 99552
box -38 -48 130 592
use scs8hd_decap_12  FILLER_178_93
timestamp 1586364061
transform 1 0 9660 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_105
timestamp 1586364061
transform 1 0 10764 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_98
timestamp 1586364061
transform 1 0 10120 0 1 99552
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_745
timestamp 1586364061
transform 1 0 12328 0 1 99552
box -38 -48 130 592
use scs8hd_decap_8  FILLER_178_117
timestamp 1586364061
transform 1 0 11868 0 -1 99552
box -38 -48 774 592
use scs8hd_decap_12  FILLER_179_110
timestamp 1586364061
transform 1 0 11224 0 1 99552
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_179_123
timestamp 1586364061
transform 1 0 12420 0 1 99552
box -38 -48 222 592
use scs8hd_decap_3  PHY_357
timestamp 1586364061
transform -1 0 12880 0 -1 99552
box -38 -48 314 592
use scs8hd_decap_3  PHY_359
timestamp 1586364061
transform -1 0 12880 0 1 99552
box -38 -48 314 592
use scs8hd_decap_3  PHY_360
timestamp 1586364061
transform 1 0 1104 0 -1 100640
box -38 -48 314 592
use scs8hd_decap_12  FILLER_180_3
timestamp 1586364061
transform 1 0 1380 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_15
timestamp 1586364061
transform 1 0 2484 0 -1 100640
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_746
timestamp 1586364061
transform 1 0 3956 0 -1 100640
box -38 -48 130 592
use scs8hd_decap_4  FILLER_180_27
timestamp 1586364061
transform 1 0 3588 0 -1 100640
box -38 -48 406 592
use scs8hd_decap_12  FILLER_180_32
timestamp 1586364061
transform 1 0 4048 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_44
timestamp 1586364061
transform 1 0 5152 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_56
timestamp 1586364061
transform 1 0 6256 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_68
timestamp 1586364061
transform 1 0 7360 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_80
timestamp 1586364061
transform 1 0 8464 0 -1 100640
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_747
timestamp 1586364061
transform 1 0 9568 0 -1 100640
box -38 -48 130 592
use scs8hd_decap_12  FILLER_180_93
timestamp 1586364061
transform 1 0 9660 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_105
timestamp 1586364061
transform 1 0 10764 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_180_117
timestamp 1586364061
transform 1 0 11868 0 -1 100640
box -38 -48 774 592
use scs8hd_decap_3  PHY_361
timestamp 1586364061
transform -1 0 12880 0 -1 100640
box -38 -48 314 592
use scs8hd_decap_3  PHY_362
timestamp 1586364061
transform 1 0 1104 0 1 100640
box -38 -48 314 592
use scs8hd_decap_12  FILLER_181_3
timestamp 1586364061
transform 1 0 1380 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_15
timestamp 1586364061
transform 1 0 2484 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_27
timestamp 1586364061
transform 1 0 3588 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_39
timestamp 1586364061
transform 1 0 4692 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_181_51
timestamp 1586364061
transform 1 0 5796 0 1 100640
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_748
timestamp 1586364061
transform 1 0 6716 0 1 100640
box -38 -48 130 592
use scs8hd_fill_2  FILLER_181_59
timestamp 1586364061
transform 1 0 6532 0 1 100640
box -38 -48 222 592
use scs8hd_decap_12  FILLER_181_62
timestamp 1586364061
transform 1 0 6808 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_74
timestamp 1586364061
transform 1 0 7912 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_86
timestamp 1586364061
transform 1 0 9016 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_98
timestamp 1586364061
transform 1 0 10120 0 1 100640
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_749
timestamp 1586364061
transform 1 0 12328 0 1 100640
box -38 -48 130 592
use scs8hd_decap_12  FILLER_181_110
timestamp 1586364061
transform 1 0 11224 0 1 100640
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_181_123
timestamp 1586364061
transform 1 0 12420 0 1 100640
box -38 -48 222 592
use scs8hd_decap_3  PHY_363
timestamp 1586364061
transform -1 0 12880 0 1 100640
box -38 -48 314 592
use scs8hd_decap_3  PHY_364
timestamp 1586364061
transform 1 0 1104 0 -1 101728
box -38 -48 314 592
use scs8hd_decap_12  FILLER_182_3
timestamp 1586364061
transform 1 0 1380 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_15
timestamp 1586364061
transform 1 0 2484 0 -1 101728
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_750
timestamp 1586364061
transform 1 0 3956 0 -1 101728
box -38 -48 130 592
use scs8hd_decap_4  FILLER_182_27
timestamp 1586364061
transform 1 0 3588 0 -1 101728
box -38 -48 406 592
use scs8hd_decap_12  FILLER_182_32
timestamp 1586364061
transform 1 0 4048 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_44
timestamp 1586364061
transform 1 0 5152 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_56
timestamp 1586364061
transform 1 0 6256 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_68
timestamp 1586364061
transform 1 0 7360 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_80
timestamp 1586364061
transform 1 0 8464 0 -1 101728
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_751
timestamp 1586364061
transform 1 0 9568 0 -1 101728
box -38 -48 130 592
use scs8hd_decap_12  FILLER_182_93
timestamp 1586364061
transform 1 0 9660 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_105
timestamp 1586364061
transform 1 0 10764 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_182_117
timestamp 1586364061
transform 1 0 11868 0 -1 101728
box -38 -48 774 592
use scs8hd_decap_3  PHY_365
timestamp 1586364061
transform -1 0 12880 0 -1 101728
box -38 -48 314 592
use scs8hd_decap_3  PHY_366
timestamp 1586364061
transform 1 0 1104 0 1 101728
box -38 -48 314 592
use scs8hd_decap_12  FILLER_183_3
timestamp 1586364061
transform 1 0 1380 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_15
timestamp 1586364061
transform 1 0 2484 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_27
timestamp 1586364061
transform 1 0 3588 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_39
timestamp 1586364061
transform 1 0 4692 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_183_51
timestamp 1586364061
transform 1 0 5796 0 1 101728
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_752
timestamp 1586364061
transform 1 0 6716 0 1 101728
box -38 -48 130 592
use scs8hd_fill_2  FILLER_183_59
timestamp 1586364061
transform 1 0 6532 0 1 101728
box -38 -48 222 592
use scs8hd_decap_12  FILLER_183_62
timestamp 1586364061
transform 1 0 6808 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_74
timestamp 1586364061
transform 1 0 7912 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_86
timestamp 1586364061
transform 1 0 9016 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_98
timestamp 1586364061
transform 1 0 10120 0 1 101728
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_753
timestamp 1586364061
transform 1 0 12328 0 1 101728
box -38 -48 130 592
use scs8hd_decap_12  FILLER_183_110
timestamp 1586364061
transform 1 0 11224 0 1 101728
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_183_123
timestamp 1586364061
transform 1 0 12420 0 1 101728
box -38 -48 222 592
use scs8hd_decap_3  PHY_367
timestamp 1586364061
transform -1 0 12880 0 1 101728
box -38 -48 314 592
use scs8hd_decap_3  PHY_368
timestamp 1586364061
transform 1 0 1104 0 -1 102816
box -38 -48 314 592
use scs8hd_decap_12  FILLER_184_3
timestamp 1586364061
transform 1 0 1380 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_15
timestamp 1586364061
transform 1 0 2484 0 -1 102816
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_754
timestamp 1586364061
transform 1 0 3956 0 -1 102816
box -38 -48 130 592
use scs8hd_decap_4  FILLER_184_27
timestamp 1586364061
transform 1 0 3588 0 -1 102816
box -38 -48 406 592
use scs8hd_decap_12  FILLER_184_32
timestamp 1586364061
transform 1 0 4048 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_44
timestamp 1586364061
transform 1 0 5152 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_56
timestamp 1586364061
transform 1 0 6256 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_68
timestamp 1586364061
transform 1 0 7360 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_80
timestamp 1586364061
transform 1 0 8464 0 -1 102816
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_755
timestamp 1586364061
transform 1 0 9568 0 -1 102816
box -38 -48 130 592
use scs8hd_decap_12  FILLER_184_93
timestamp 1586364061
transform 1 0 9660 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_105
timestamp 1586364061
transform 1 0 10764 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_184_117
timestamp 1586364061
transform 1 0 11868 0 -1 102816
box -38 -48 774 592
use scs8hd_decap_3  PHY_369
timestamp 1586364061
transform -1 0 12880 0 -1 102816
box -38 -48 314 592
use scs8hd_decap_3  PHY_370
timestamp 1586364061
transform 1 0 1104 0 1 102816
box -38 -48 314 592
use scs8hd_decap_3  PHY_372
timestamp 1586364061
transform 1 0 1104 0 -1 103904
box -38 -48 314 592
use scs8hd_decap_12  FILLER_185_3
timestamp 1586364061
transform 1 0 1380 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_185_15
timestamp 1586364061
transform 1 0 2484 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_3
timestamp 1586364061
transform 1 0 1380 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_15
timestamp 1586364061
transform 1 0 2484 0 -1 103904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_758
timestamp 1586364061
transform 1 0 3956 0 -1 103904
box -38 -48 130 592
use scs8hd_decap_12  FILLER_185_27
timestamp 1586364061
transform 1 0 3588 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_186_27
timestamp 1586364061
transform 1 0 3588 0 -1 103904
box -38 -48 406 592
use scs8hd_decap_12  FILLER_186_32
timestamp 1586364061
transform 1 0 4048 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_185_39
timestamp 1586364061
transform 1 0 4692 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_185_51
timestamp 1586364061
transform 1 0 5796 0 1 102816
box -38 -48 774 592
use scs8hd_decap_12  FILLER_186_44
timestamp 1586364061
transform 1 0 5152 0 -1 103904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_756
timestamp 1586364061
transform 1 0 6716 0 1 102816
box -38 -48 130 592
use scs8hd_fill_2  FILLER_185_59
timestamp 1586364061
transform 1 0 6532 0 1 102816
box -38 -48 222 592
use scs8hd_decap_12  FILLER_185_62
timestamp 1586364061
transform 1 0 6808 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_56
timestamp 1586364061
transform 1 0 6256 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_68
timestamp 1586364061
transform 1 0 7360 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_185_74
timestamp 1586364061
transform 1 0 7912 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_185_86
timestamp 1586364061
transform 1 0 9016 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_80
timestamp 1586364061
transform 1 0 8464 0 -1 103904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_759
timestamp 1586364061
transform 1 0 9568 0 -1 103904
box -38 -48 130 592
use scs8hd_decap_12  FILLER_185_98
timestamp 1586364061
transform 1 0 10120 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_93
timestamp 1586364061
transform 1 0 9660 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_105
timestamp 1586364061
transform 1 0 10764 0 -1 103904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_757
timestamp 1586364061
transform 1 0 12328 0 1 102816
box -38 -48 130 592
use scs8hd_decap_12  FILLER_185_110
timestamp 1586364061
transform 1 0 11224 0 1 102816
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_185_123
timestamp 1586364061
transform 1 0 12420 0 1 102816
box -38 -48 222 592
use scs8hd_decap_8  FILLER_186_117
timestamp 1586364061
transform 1 0 11868 0 -1 103904
box -38 -48 774 592
use scs8hd_decap_3  PHY_371
timestamp 1586364061
transform -1 0 12880 0 1 102816
box -38 -48 314 592
use scs8hd_decap_3  PHY_373
timestamp 1586364061
transform -1 0 12880 0 -1 103904
box -38 -48 314 592
use scs8hd_decap_3  PHY_374
timestamp 1586364061
transform 1 0 1104 0 1 103904
box -38 -48 314 592
use scs8hd_decap_12  FILLER_187_3
timestamp 1586364061
transform 1 0 1380 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_15
timestamp 1586364061
transform 1 0 2484 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_27
timestamp 1586364061
transform 1 0 3588 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_39
timestamp 1586364061
transform 1 0 4692 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_187_51
timestamp 1586364061
transform 1 0 5796 0 1 103904
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_760
timestamp 1586364061
transform 1 0 6716 0 1 103904
box -38 -48 130 592
use scs8hd_fill_2  FILLER_187_59
timestamp 1586364061
transform 1 0 6532 0 1 103904
box -38 -48 222 592
use scs8hd_decap_12  FILLER_187_62
timestamp 1586364061
transform 1 0 6808 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_74
timestamp 1586364061
transform 1 0 7912 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_86
timestamp 1586364061
transform 1 0 9016 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_98
timestamp 1586364061
transform 1 0 10120 0 1 103904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_761
timestamp 1586364061
transform 1 0 12328 0 1 103904
box -38 -48 130 592
use scs8hd_decap_12  FILLER_187_110
timestamp 1586364061
transform 1 0 11224 0 1 103904
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_187_123
timestamp 1586364061
transform 1 0 12420 0 1 103904
box -38 -48 222 592
use scs8hd_decap_3  PHY_375
timestamp 1586364061
transform -1 0 12880 0 1 103904
box -38 -48 314 592
use scs8hd_decap_3  PHY_376
timestamp 1586364061
transform 1 0 1104 0 -1 104992
box -38 -48 314 592
use scs8hd_decap_12  FILLER_188_3
timestamp 1586364061
transform 1 0 1380 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_15
timestamp 1586364061
transform 1 0 2484 0 -1 104992
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_762
timestamp 1586364061
transform 1 0 3956 0 -1 104992
box -38 -48 130 592
use scs8hd_decap_4  FILLER_188_27
timestamp 1586364061
transform 1 0 3588 0 -1 104992
box -38 -48 406 592
use scs8hd_decap_12  FILLER_188_32
timestamp 1586364061
transform 1 0 4048 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_44
timestamp 1586364061
transform 1 0 5152 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_56
timestamp 1586364061
transform 1 0 6256 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_68
timestamp 1586364061
transform 1 0 7360 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_80
timestamp 1586364061
transform 1 0 8464 0 -1 104992
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_763
timestamp 1586364061
transform 1 0 9568 0 -1 104992
box -38 -48 130 592
use scs8hd_decap_12  FILLER_188_93
timestamp 1586364061
transform 1 0 9660 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_105
timestamp 1586364061
transform 1 0 10764 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_188_117
timestamp 1586364061
transform 1 0 11868 0 -1 104992
box -38 -48 774 592
use scs8hd_decap_3  PHY_377
timestamp 1586364061
transform -1 0 12880 0 -1 104992
box -38 -48 314 592
use scs8hd_decap_3  PHY_378
timestamp 1586364061
transform 1 0 1104 0 1 104992
box -38 -48 314 592
use scs8hd_decap_12  FILLER_189_3
timestamp 1586364061
transform 1 0 1380 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_15
timestamp 1586364061
transform 1 0 2484 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_27
timestamp 1586364061
transform 1 0 3588 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_39
timestamp 1586364061
transform 1 0 4692 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_189_51
timestamp 1586364061
transform 1 0 5796 0 1 104992
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_764
timestamp 1586364061
transform 1 0 6716 0 1 104992
box -38 -48 130 592
use scs8hd_fill_2  FILLER_189_59
timestamp 1586364061
transform 1 0 6532 0 1 104992
box -38 -48 222 592
use scs8hd_decap_12  FILLER_189_62
timestamp 1586364061
transform 1 0 6808 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_74
timestamp 1586364061
transform 1 0 7912 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_86
timestamp 1586364061
transform 1 0 9016 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_98
timestamp 1586364061
transform 1 0 10120 0 1 104992
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_765
timestamp 1586364061
transform 1 0 12328 0 1 104992
box -38 -48 130 592
use scs8hd_decap_12  FILLER_189_110
timestamp 1586364061
transform 1 0 11224 0 1 104992
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_189_123
timestamp 1586364061
transform 1 0 12420 0 1 104992
box -38 -48 222 592
use scs8hd_decap_3  PHY_379
timestamp 1586364061
transform -1 0 12880 0 1 104992
box -38 -48 314 592
use scs8hd_decap_3  PHY_380
timestamp 1586364061
transform 1 0 1104 0 -1 106080
box -38 -48 314 592
use scs8hd_decap_12  FILLER_190_3
timestamp 1586364061
transform 1 0 1380 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_15
timestamp 1586364061
transform 1 0 2484 0 -1 106080
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_766
timestamp 1586364061
transform 1 0 3956 0 -1 106080
box -38 -48 130 592
use scs8hd_decap_4  FILLER_190_27
timestamp 1586364061
transform 1 0 3588 0 -1 106080
box -38 -48 406 592
use scs8hd_decap_12  FILLER_190_32
timestamp 1586364061
transform 1 0 4048 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_44
timestamp 1586364061
transform 1 0 5152 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_56
timestamp 1586364061
transform 1 0 6256 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_68
timestamp 1586364061
transform 1 0 7360 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_80
timestamp 1586364061
transform 1 0 8464 0 -1 106080
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_767
timestamp 1586364061
transform 1 0 9568 0 -1 106080
box -38 -48 130 592
use scs8hd_decap_12  FILLER_190_93
timestamp 1586364061
transform 1 0 9660 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_105
timestamp 1586364061
transform 1 0 10764 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_190_117
timestamp 1586364061
transform 1 0 11868 0 -1 106080
box -38 -48 774 592
use scs8hd_decap_3  PHY_381
timestamp 1586364061
transform -1 0 12880 0 -1 106080
box -38 -48 314 592
use scs8hd_decap_3  PHY_382
timestamp 1586364061
transform 1 0 1104 0 1 106080
box -38 -48 314 592
use scs8hd_decap_12  FILLER_191_3
timestamp 1586364061
transform 1 0 1380 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_191_15
timestamp 1586364061
transform 1 0 2484 0 1 106080
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_768
timestamp 1586364061
transform 1 0 3956 0 1 106080
box -38 -48 130 592
use scs8hd_decap_4  FILLER_191_27
timestamp 1586364061
transform 1 0 3588 0 1 106080
box -38 -48 406 592
use scs8hd_decap_12  FILLER_191_32
timestamp 1586364061
transform 1 0 4048 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_191_44
timestamp 1586364061
transform 1 0 5152 0 1 106080
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_769
timestamp 1586364061
transform 1 0 6808 0 1 106080
box -38 -48 130 592
use scs8hd_decap_6  FILLER_191_56
timestamp 1586364061
transform 1 0 6256 0 1 106080
box -38 -48 590 592
use scs8hd_decap_12  FILLER_191_63
timestamp 1586364061
transform 1 0 6900 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_191_75
timestamp 1586364061
transform 1 0 8004 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_191_87
timestamp 1586364061
transform 1 0 9108 0 1 106080
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_770
timestamp 1586364061
transform 1 0 9660 0 1 106080
box -38 -48 130 592
use scs8hd_decap_12  FILLER_191_94
timestamp 1586364061
transform 1 0 9752 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_191_106
timestamp 1586364061
transform 1 0 10856 0 1 106080
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_771
timestamp 1586364061
transform 1 0 12512 0 1 106080
box -38 -48 130 592
use scs8hd_decap_6  FILLER_191_118
timestamp 1586364061
transform 1 0 11960 0 1 106080
box -38 -48 590 592
use scs8hd_decap_3  PHY_383
timestamp 1586364061
transform -1 0 12880 0 1 106080
box -38 -48 314 592
<< labels >>
rlabel metal2 s 3422 0 3478 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 5722 0 5778 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 8114 0 8170 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 10414 0 10470 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 12714 0 12770 480 6 data_in
port 4 nsew default input
rlabel metal2 s 1122 0 1178 480 6 enable
port 5 nsew default input
rlabel metal3 s 0 6808 480 6928 6 gfpga_pad_GPIO_PAD[0]
port 6 nsew default bidirectional
rlabel metal3 s 0 20408 480 20528 6 gfpga_pad_GPIO_PAD[1]
port 7 nsew default bidirectional
rlabel metal3 s 0 34008 480 34128 6 gfpga_pad_GPIO_PAD[2]
port 8 nsew default bidirectional
rlabel metal3 s 0 47608 480 47728 6 gfpga_pad_GPIO_PAD[3]
port 9 nsew default bidirectional
rlabel metal3 s 0 61208 480 61328 6 gfpga_pad_GPIO_PAD[4]
port 10 nsew default bidirectional
rlabel metal3 s 0 74808 480 74928 6 gfpga_pad_GPIO_PAD[5]
port 11 nsew default bidirectional
rlabel metal3 s 0 88408 480 88528 6 gfpga_pad_GPIO_PAD[6]
port 12 nsew default bidirectional
rlabel metal3 s 0 102008 480 102128 6 gfpga_pad_GPIO_PAD[7]
port 13 nsew default bidirectional
rlabel metal3 s 13520 3408 14000 3528 6 right_width_0_height_0__pin_0_
port 14 nsew default input
rlabel metal3 s 13520 71408 14000 71528 6 right_width_0_height_0__pin_10_
port 15 nsew default input
rlabel metal3 s 13520 78208 14000 78328 6 right_width_0_height_0__pin_11_
port 16 nsew default tristate
rlabel metal3 s 13520 85008 14000 85128 6 right_width_0_height_0__pin_12_
port 17 nsew default input
rlabel metal3 s 13520 91808 14000 91928 6 right_width_0_height_0__pin_13_
port 18 nsew default tristate
rlabel metal3 s 13520 98608 14000 98728 6 right_width_0_height_0__pin_14_
port 19 nsew default input
rlabel metal3 s 13520 105408 14000 105528 6 right_width_0_height_0__pin_15_
port 20 nsew default tristate
rlabel metal3 s 13520 10208 14000 10328 6 right_width_0_height_0__pin_1_
port 21 nsew default tristate
rlabel metal3 s 13520 17008 14000 17128 6 right_width_0_height_0__pin_2_
port 22 nsew default input
rlabel metal3 s 13520 23808 14000 23928 6 right_width_0_height_0__pin_3_
port 23 nsew default tristate
rlabel metal3 s 13520 30608 14000 30728 6 right_width_0_height_0__pin_4_
port 24 nsew default input
rlabel metal3 s 13520 37408 14000 37528 6 right_width_0_height_0__pin_5_
port 25 nsew default tristate
rlabel metal3 s 13520 44208 14000 44328 6 right_width_0_height_0__pin_6_
port 26 nsew default input
rlabel metal3 s 13520 51008 14000 51128 6 right_width_0_height_0__pin_7_
port 27 nsew default tristate
rlabel metal3 s 13520 57808 14000 57928 6 right_width_0_height_0__pin_8_
port 28 nsew default input
rlabel metal3 s 13520 64608 14000 64728 6 right_width_0_height_0__pin_9_
port 29 nsew default tristate
rlabel metal4 s 3277 2128 3597 106672 6 vpwr
port 30 nsew default input
rlabel metal4 s 5611 2128 5931 106672 6 vgnd
port 31 nsew default input
<< end >>
