VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__1_
  CLASS BLOCK ;
  FOREIGN cbx_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 85.000 ;
  PIN REGIN_FEEDTHROUGH
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END REGIN_FEEDTHROUGH
  PIN REGOUT_FEEDTHROUGH
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END REGOUT_FEEDTHROUGH
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 81.000 10.030 85.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.530 81.000 29.810 85.000 ;
    END
  END SC_OUT_TOP
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END bottom_grid_pin_11_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END bottom_grid_pin_13_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END bottom_grid_pin_15_
  PIN bottom_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END bottom_grid_pin_1_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END bottom_grid_pin_3_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END bottom_grid_pin_5_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END bottom_grid_pin_7_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END bottom_grid_pin_8_
  PIN bottom_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END bottom_grid_pin_9_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.720 100.000 52.320 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.720 100.000 69.320 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.080 100.000 70.680 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 72.120 100.000 72.720 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 73.480 100.000 74.080 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 75.520 100.000 76.120 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 76.880 100.000 77.480 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 78.920 100.000 79.520 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 80.280 100.000 80.880 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 82.320 100.000 82.920 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 83.680 100.000 84.280 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 53.760 100.000 54.360 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.120 100.000 55.720 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 57.160 100.000 57.760 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 58.520 100.000 59.120 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 60.560 100.000 61.160 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 61.920 100.000 62.520 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 63.960 100.000 64.560 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 65.320 100.000 65.920 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 67.360 100.000 67.960 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 18.400 100.000 19.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 35.400 100.000 36.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 36.760 100.000 37.360 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 38.800 100.000 39.400 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 40.160 100.000 40.760 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 42.200 100.000 42.800 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.560 100.000 44.160 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 45.600 100.000 46.200 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 46.960 100.000 47.560 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 49.000 100.000 49.600 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 50.360 100.000 50.960 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 20.440 100.000 21.040 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 21.800 100.000 22.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 23.840 100.000 24.440 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 25.200 100.000 25.800 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 27.240 100.000 27.840 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 28.600 100.000 29.200 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 30.640 100.000 31.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 32.000 100.000 32.600 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 34.040 100.000 34.640 ;
    END
  END chanx_right_out[9]
  PIN clk_1_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 17.040 100.000 17.640 ;
    END
  END clk_1_E_in
  PIN clk_1_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.310 81.000 49.590 85.000 ;
    END
  END clk_1_N_out
  PIN clk_1_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END clk_1_S_out
  PIN clk_1_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END clk_1_W_in
  PIN clk_2_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 15.680 100.000 16.280 ;
    END
  END clk_2_E_in
  PIN clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END clk_2_E_out
  PIN clk_2_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END clk_2_W_in
  PIN clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END clk_2_W_out
  PIN clk_3_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 13.640 100.000 14.240 ;
    END
  END clk_3_E_in
  PIN clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 5.480 100.000 6.080 ;
    END
  END clk_3_E_out
  PIN clk_3_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END clk_3_W_in
  PIN clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END clk_3_W_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 81.000 69.830 85.000 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.330 81.000 89.610 85.000 ;
    END
  END prog_clk_0_W_out
  PIN prog_clk_1_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 12.280 100.000 12.880 ;
    END
  END prog_clk_1_E_in
  PIN prog_clk_1_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END prog_clk_1_N_out
  PIN prog_clk_1_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END prog_clk_1_S_out
  PIN prog_clk_1_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END prog_clk_1_W_in
  PIN prog_clk_2_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.240 100.000 10.840 ;
    END
  END prog_clk_2_E_in
  PIN prog_clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 2.080 100.000 2.680 ;
    END
  END prog_clk_2_E_out
  PIN prog_clk_2_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END prog_clk_2_W_in
  PIN prog_clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END prog_clk_2_W_out
  PIN prog_clk_3_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 96.000 8.880 100.000 9.480 ;
    END
  END prog_clk_3_E_in
  PIN prog_clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 96.000 0.720 100.000 1.320 ;
    END
  END prog_clk_3_E_out
  PIN prog_clk_3_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END prog_clk_3_W_in
  PIN prog_clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END prog_clk_3_W_out
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.375 10.640 35.975 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 73.525 ;
      LAYER met1 ;
        RECT 1.910 6.500 97.450 76.460 ;
      LAYER met2 ;
        RECT 1.940 80.720 9.470 84.165 ;
        RECT 10.310 80.720 29.250 84.165 ;
        RECT 30.090 80.720 49.030 84.165 ;
        RECT 49.870 80.720 69.270 84.165 ;
        RECT 70.110 80.720 89.050 84.165 ;
        RECT 89.890 80.720 97.420 84.165 ;
        RECT 1.940 4.280 97.420 80.720 ;
        RECT 2.490 0.835 5.790 4.280 ;
        RECT 6.630 0.835 10.390 4.280 ;
        RECT 11.230 0.835 14.990 4.280 ;
        RECT 15.830 0.835 19.590 4.280 ;
        RECT 20.430 0.835 24.190 4.280 ;
        RECT 25.030 0.835 28.790 4.280 ;
        RECT 29.630 0.835 33.390 4.280 ;
        RECT 34.230 0.835 37.530 4.280 ;
        RECT 38.370 0.835 42.130 4.280 ;
        RECT 42.970 0.835 46.730 4.280 ;
        RECT 47.570 0.835 51.330 4.280 ;
        RECT 52.170 0.835 55.930 4.280 ;
        RECT 56.770 0.835 60.530 4.280 ;
        RECT 61.370 0.835 65.130 4.280 ;
        RECT 65.970 0.835 69.270 4.280 ;
        RECT 70.110 0.835 73.870 4.280 ;
        RECT 74.710 0.835 78.470 4.280 ;
        RECT 79.310 0.835 83.070 4.280 ;
        RECT 83.910 0.835 87.670 4.280 ;
        RECT 88.510 0.835 92.270 4.280 ;
        RECT 93.110 0.835 96.870 4.280 ;
      LAYER met3 ;
        RECT 4.400 81.920 95.600 84.145 ;
        RECT 3.990 81.280 96.000 81.920 ;
        RECT 4.400 78.520 95.600 81.280 ;
        RECT 3.990 77.880 96.000 78.520 ;
        RECT 4.400 75.120 95.600 77.880 ;
        RECT 4.400 74.480 96.000 75.120 ;
        RECT 4.400 73.760 95.600 74.480 ;
        RECT 3.990 73.120 95.600 73.760 ;
        RECT 4.400 71.720 95.600 73.120 ;
        RECT 4.400 71.080 96.000 71.720 ;
        RECT 4.400 70.360 95.600 71.080 ;
        RECT 3.990 69.720 95.600 70.360 ;
        RECT 4.400 66.960 95.600 69.720 ;
        RECT 4.400 66.320 96.000 66.960 ;
        RECT 4.400 65.600 95.600 66.320 ;
        RECT 3.990 64.960 95.600 65.600 ;
        RECT 4.400 63.560 95.600 64.960 ;
        RECT 4.400 62.920 96.000 63.560 ;
        RECT 4.400 62.200 95.600 62.920 ;
        RECT 3.990 61.560 95.600 62.200 ;
        RECT 4.400 60.160 95.600 61.560 ;
        RECT 4.400 59.520 96.000 60.160 ;
        RECT 4.400 57.440 95.600 59.520 ;
        RECT 3.990 56.800 95.600 57.440 ;
        RECT 4.400 56.760 95.600 56.800 ;
        RECT 4.400 56.120 96.000 56.760 ;
        RECT 4.400 54.040 95.600 56.120 ;
        RECT 3.990 53.400 95.600 54.040 ;
        RECT 4.400 53.360 95.600 53.400 ;
        RECT 4.400 52.720 96.000 53.360 ;
        RECT 4.400 49.280 95.600 52.720 ;
        RECT 3.990 48.640 95.600 49.280 ;
        RECT 4.400 48.600 95.600 48.640 ;
        RECT 4.400 47.960 96.000 48.600 ;
        RECT 4.400 45.880 95.600 47.960 ;
        RECT 3.990 45.240 95.600 45.880 ;
        RECT 4.400 45.200 95.600 45.240 ;
        RECT 4.400 44.560 96.000 45.200 ;
        RECT 4.400 41.800 95.600 44.560 ;
        RECT 4.400 41.160 96.000 41.800 ;
        RECT 4.400 41.120 95.600 41.160 ;
        RECT 3.990 40.480 95.600 41.120 ;
        RECT 4.400 38.400 95.600 40.480 ;
        RECT 4.400 37.760 96.000 38.400 ;
        RECT 4.400 37.720 95.600 37.760 ;
        RECT 3.990 37.080 95.600 37.720 ;
        RECT 4.400 33.640 95.600 37.080 ;
        RECT 4.400 33.000 96.000 33.640 ;
        RECT 4.400 32.960 95.600 33.000 ;
        RECT 3.990 32.320 95.600 32.960 ;
        RECT 4.400 30.240 95.600 32.320 ;
        RECT 4.400 29.600 96.000 30.240 ;
        RECT 4.400 29.560 95.600 29.600 ;
        RECT 3.990 28.920 95.600 29.560 ;
        RECT 4.400 26.840 95.600 28.920 ;
        RECT 4.400 26.200 96.000 26.840 ;
        RECT 4.400 24.800 95.600 26.200 ;
        RECT 3.990 24.160 95.600 24.800 ;
        RECT 4.400 23.440 95.600 24.160 ;
        RECT 4.400 22.800 96.000 23.440 ;
        RECT 4.400 21.400 95.600 22.800 ;
        RECT 3.990 20.760 95.600 21.400 ;
        RECT 4.400 20.040 95.600 20.760 ;
        RECT 4.400 19.400 96.000 20.040 ;
        RECT 4.400 16.640 95.600 19.400 ;
        RECT 3.990 16.000 95.600 16.640 ;
        RECT 4.400 15.280 95.600 16.000 ;
        RECT 4.400 14.640 96.000 15.280 ;
        RECT 4.400 13.240 95.600 14.640 ;
        RECT 3.990 12.600 95.600 13.240 ;
        RECT 4.400 11.880 95.600 12.600 ;
        RECT 4.400 11.240 96.000 11.880 ;
        RECT 4.400 8.480 95.600 11.240 ;
        RECT 3.990 7.840 96.000 8.480 ;
        RECT 4.400 5.080 95.600 7.840 ;
        RECT 3.990 4.440 96.000 5.080 ;
        RECT 4.400 0.855 95.600 4.440 ;
      LAYER met4 ;
        RECT 22.375 74.080 86.185 84.145 ;
        RECT 22.375 10.640 33.975 74.080 ;
        RECT 36.375 10.640 86.185 74.080 ;
  END
END cbx_1__1_
END LIBRARY

