VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 115.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.400 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 112.600 1.290 115.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.400 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 112.600 113.990 115.000 ;
    END
  END SC_OUT_TOP
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 2.400 18.320 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 2.400 21.040 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 2.400 23.760 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.400 31.240 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 2.400 91.080 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 2.400 78.160 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 2.400 88.360 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 15.680 115.000 16.280 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 40.160 115.000 40.760 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 42.880 115.000 43.480 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 45.600 115.000 46.200 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 47.640 115.000 48.240 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 50.360 115.000 50.960 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 53.080 115.000 53.680 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 55.120 115.000 55.720 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 57.840 115.000 58.440 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 60.560 115.000 61.160 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 62.600 115.000 63.200 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 17.720 115.000 18.320 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 20.440 115.000 21.040 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 23.160 115.000 23.760 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 25.200 115.000 25.800 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 27.920 115.000 28.520 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 30.640 115.000 31.240 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 32.680 115.000 33.280 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 35.400 115.000 36.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 38.120 115.000 38.720 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 65.320 115.000 65.920 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 90.480 115.000 91.080 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 92.520 115.000 93.120 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 95.240 115.000 95.840 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 97.960 115.000 98.560 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 100.000 115.000 100.600 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 102.720 115.000 103.320 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 105.440 115.000 106.040 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 107.480 115.000 108.080 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 110.200 115.000 110.800 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 112.920 115.000 113.520 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 68.040 115.000 68.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 70.080 115.000 70.680 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 72.800 115.000 73.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 75.520 115.000 76.120 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 77.560 115.000 78.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 80.280 115.000 80.880 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 83.000 115.000 83.600 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 85.040 115.000 85.640 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 87.760 115.000 88.360 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 112.600 21.990 115.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 112.600 44.990 115.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 112.600 47.290 115.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 112.600 49.590 115.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 112.600 51.890 115.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 112.600 54.190 115.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 112.600 56.490 115.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 112.600 58.790 115.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 112.600 61.090 115.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 112.600 63.390 115.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 112.600 65.690 115.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 112.600 24.290 115.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 112.600 26.590 115.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 112.600 28.890 115.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 112.600 31.190 115.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 112.600 33.490 115.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 112.600 35.790 115.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 112.600 38.090 115.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 112.600 40.390 115.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 112.600 42.690 115.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 112.600 67.990 115.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.710 112.600 90.990 115.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 112.600 93.290 115.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 112.600 95.590 115.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 112.600 97.890 115.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.910 112.600 100.190 115.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 112.600 102.490 115.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 112.600 104.790 115.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 112.600 107.090 115.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.110 112.600 109.390 115.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.410 112.600 111.690 115.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 112.600 70.290 115.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 112.600 72.590 115.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 112.600 74.890 115.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 112.600 77.190 115.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 112.600 79.490 115.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.510 112.600 81.790 115.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 112.600 84.090 115.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.110 112.600 86.390 115.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 112.600 88.690 115.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 2.400 6.080 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END left_bottom_grid_pin_9_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 12.960 115.000 13.560 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 0.720 115.000 1.320 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 2.760 115.000 3.360 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 5.480 115.000 6.080 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 8.200 115.000 8.800 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 10.240 115.000 10.840 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 112.600 3.590 115.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 112.600 5.890 115.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 112.600 8.190 115.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 112.600 10.490 115.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 112.600 12.790 115.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 112.600 15.090 115.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 112.600 17.390 115.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 112.600 19.690 115.000 ;
    END
  END top_left_grid_pin_49_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.045 10.640 23.645 103.600 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.375 10.640 40.975 103.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 8.245 109.480 103.445 ;
      LAYER met1 ;
        RECT 0.070 6.160 114.010 108.420 ;
      LAYER met2 ;
        RECT 0.090 112.320 0.730 113.405 ;
        RECT 1.570 112.320 3.030 113.405 ;
        RECT 3.870 112.320 5.330 113.405 ;
        RECT 6.170 112.320 7.630 113.405 ;
        RECT 8.470 112.320 9.930 113.405 ;
        RECT 10.770 112.320 12.230 113.405 ;
        RECT 13.070 112.320 14.530 113.405 ;
        RECT 15.370 112.320 16.830 113.405 ;
        RECT 17.670 112.320 19.130 113.405 ;
        RECT 19.970 112.320 21.430 113.405 ;
        RECT 22.270 112.320 23.730 113.405 ;
        RECT 24.570 112.320 26.030 113.405 ;
        RECT 26.870 112.320 28.330 113.405 ;
        RECT 29.170 112.320 30.630 113.405 ;
        RECT 31.470 112.320 32.930 113.405 ;
        RECT 33.770 112.320 35.230 113.405 ;
        RECT 36.070 112.320 37.530 113.405 ;
        RECT 38.370 112.320 39.830 113.405 ;
        RECT 40.670 112.320 42.130 113.405 ;
        RECT 42.970 112.320 44.430 113.405 ;
        RECT 45.270 112.320 46.730 113.405 ;
        RECT 47.570 112.320 49.030 113.405 ;
        RECT 49.870 112.320 51.330 113.405 ;
        RECT 52.170 112.320 53.630 113.405 ;
        RECT 54.470 112.320 55.930 113.405 ;
        RECT 56.770 112.320 58.230 113.405 ;
        RECT 59.070 112.320 60.530 113.405 ;
        RECT 61.370 112.320 62.830 113.405 ;
        RECT 63.670 112.320 65.130 113.405 ;
        RECT 65.970 112.320 67.430 113.405 ;
        RECT 68.270 112.320 69.730 113.405 ;
        RECT 70.570 112.320 72.030 113.405 ;
        RECT 72.870 112.320 74.330 113.405 ;
        RECT 75.170 112.320 76.630 113.405 ;
        RECT 77.470 112.320 78.930 113.405 ;
        RECT 79.770 112.320 81.230 113.405 ;
        RECT 82.070 112.320 83.530 113.405 ;
        RECT 84.370 112.320 85.830 113.405 ;
        RECT 86.670 112.320 88.130 113.405 ;
        RECT 88.970 112.320 90.430 113.405 ;
        RECT 91.270 112.320 92.730 113.405 ;
        RECT 93.570 112.320 95.030 113.405 ;
        RECT 95.870 112.320 97.330 113.405 ;
        RECT 98.170 112.320 99.630 113.405 ;
        RECT 100.470 112.320 101.930 113.405 ;
        RECT 102.770 112.320 104.230 113.405 ;
        RECT 105.070 112.320 106.530 113.405 ;
        RECT 107.370 112.320 108.830 113.405 ;
        RECT 109.670 112.320 111.130 113.405 ;
        RECT 111.970 112.320 113.430 113.405 ;
        RECT 0.090 2.680 113.980 112.320 ;
        RECT 0.090 0.835 11.310 2.680 ;
        RECT 12.150 0.835 34.310 2.680 ;
        RECT 35.150 0.835 57.310 2.680 ;
        RECT 58.150 0.835 80.310 2.680 ;
        RECT 81.150 0.835 103.310 2.680 ;
        RECT 104.150 0.835 113.980 2.680 ;
      LAYER met3 ;
        RECT 2.800 112.520 112.200 113.385 ;
        RECT 0.065 111.200 112.600 112.520 ;
        RECT 2.800 109.800 112.200 111.200 ;
        RECT 0.065 108.480 112.600 109.800 ;
        RECT 2.800 107.080 112.200 108.480 ;
        RECT 0.065 106.440 112.600 107.080 ;
        RECT 2.800 105.040 112.200 106.440 ;
        RECT 0.065 103.720 112.600 105.040 ;
        RECT 2.800 102.320 112.200 103.720 ;
        RECT 0.065 101.000 112.600 102.320 ;
        RECT 2.800 99.600 112.200 101.000 ;
        RECT 0.065 98.960 112.600 99.600 ;
        RECT 2.800 97.560 112.200 98.960 ;
        RECT 0.065 96.240 112.600 97.560 ;
        RECT 2.800 94.840 112.200 96.240 ;
        RECT 0.065 93.520 112.600 94.840 ;
        RECT 2.800 92.120 112.200 93.520 ;
        RECT 0.065 91.480 112.600 92.120 ;
        RECT 2.800 90.080 112.200 91.480 ;
        RECT 0.065 88.760 112.600 90.080 ;
        RECT 2.800 87.360 112.200 88.760 ;
        RECT 0.065 86.040 112.600 87.360 ;
        RECT 2.800 84.640 112.200 86.040 ;
        RECT 0.065 84.000 112.600 84.640 ;
        RECT 2.800 82.600 112.200 84.000 ;
        RECT 0.065 81.280 112.600 82.600 ;
        RECT 2.800 79.880 112.200 81.280 ;
        RECT 0.065 78.560 112.600 79.880 ;
        RECT 2.800 77.160 112.200 78.560 ;
        RECT 0.065 76.520 112.600 77.160 ;
        RECT 2.800 75.120 112.200 76.520 ;
        RECT 0.065 73.800 112.600 75.120 ;
        RECT 2.800 72.400 112.200 73.800 ;
        RECT 0.065 71.080 112.600 72.400 ;
        RECT 2.800 69.680 112.200 71.080 ;
        RECT 0.065 69.040 112.600 69.680 ;
        RECT 2.800 67.640 112.200 69.040 ;
        RECT 0.065 66.320 112.600 67.640 ;
        RECT 2.800 64.920 112.200 66.320 ;
        RECT 0.065 63.600 112.600 64.920 ;
        RECT 2.800 62.200 112.200 63.600 ;
        RECT 0.065 61.560 112.600 62.200 ;
        RECT 2.800 60.160 112.200 61.560 ;
        RECT 0.065 58.840 112.600 60.160 ;
        RECT 2.800 57.440 112.200 58.840 ;
        RECT 0.065 56.120 112.600 57.440 ;
        RECT 2.800 54.720 112.200 56.120 ;
        RECT 0.065 54.080 112.600 54.720 ;
        RECT 2.800 52.680 112.200 54.080 ;
        RECT 0.065 51.360 112.600 52.680 ;
        RECT 2.800 49.960 112.200 51.360 ;
        RECT 0.065 48.640 112.600 49.960 ;
        RECT 2.800 47.240 112.200 48.640 ;
        RECT 0.065 46.600 112.600 47.240 ;
        RECT 2.800 45.200 112.200 46.600 ;
        RECT 0.065 43.880 112.600 45.200 ;
        RECT 2.800 42.480 112.200 43.880 ;
        RECT 0.065 41.160 112.600 42.480 ;
        RECT 2.800 39.760 112.200 41.160 ;
        RECT 0.065 39.120 112.600 39.760 ;
        RECT 2.800 37.720 112.200 39.120 ;
        RECT 0.065 36.400 112.600 37.720 ;
        RECT 2.800 35.000 112.200 36.400 ;
        RECT 0.065 33.680 112.600 35.000 ;
        RECT 2.800 32.280 112.200 33.680 ;
        RECT 0.065 31.640 112.600 32.280 ;
        RECT 2.800 30.240 112.200 31.640 ;
        RECT 0.065 28.920 112.600 30.240 ;
        RECT 2.800 27.520 112.200 28.920 ;
        RECT 0.065 26.200 112.600 27.520 ;
        RECT 2.800 24.800 112.200 26.200 ;
        RECT 0.065 24.160 112.600 24.800 ;
        RECT 2.800 22.760 112.200 24.160 ;
        RECT 0.065 21.440 112.600 22.760 ;
        RECT 2.800 20.040 112.200 21.440 ;
        RECT 0.065 18.720 112.600 20.040 ;
        RECT 2.800 17.320 112.200 18.720 ;
        RECT 0.065 16.680 112.600 17.320 ;
        RECT 2.800 15.280 112.200 16.680 ;
        RECT 0.065 13.960 112.600 15.280 ;
        RECT 2.800 12.560 112.200 13.960 ;
        RECT 0.065 11.240 112.600 12.560 ;
        RECT 2.800 9.840 112.200 11.240 ;
        RECT 0.065 9.200 112.600 9.840 ;
        RECT 2.800 7.800 112.200 9.200 ;
        RECT 0.065 6.480 112.600 7.800 ;
        RECT 2.800 5.080 112.200 6.480 ;
        RECT 0.065 3.760 112.600 5.080 ;
        RECT 2.800 2.360 112.200 3.760 ;
        RECT 0.065 1.720 112.600 2.360 ;
        RECT 2.800 0.855 112.200 1.720 ;
      LAYER met4 ;
        RECT 9.495 10.640 21.645 103.600 ;
        RECT 24.045 10.640 38.975 103.600 ;
        RECT 41.375 10.640 99.065 103.600 ;
  END
END sb_1__0_
END LIBRARY

