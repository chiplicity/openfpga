VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_0__1_
  CLASS BLOCK ;
  FOREIGN cby_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 197.600 41.310 200.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 197.600 61.090 200.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 197.600 62.930 200.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 197.600 65.230 200.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 197.600 67.070 200.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 197.600 68.910 200.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 197.600 71.210 200.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 197.600 73.050 200.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 197.600 74.890 200.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 197.600 77.190 200.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 197.600 79.030 200.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 197.600 43.150 200.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 197.600 44.990 200.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 197.600 47.290 200.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 197.600 49.130 200.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 197.600 50.970 200.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 197.600 53.270 200.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 197.600 55.110 200.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 197.600 56.950 200.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 197.600 59.250 200.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.010 197.600 1.290 200.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.790 197.600 21.070 200.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 197.600 22.910 200.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 197.600 25.210 200.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 197.600 27.050 200.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 197.600 28.890 200.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 197.600 31.190 200.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.750 197.600 33.030 200.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 197.600 34.870 200.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 197.600 37.170 200.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.730 197.600 39.010 200.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 197.600 3.130 200.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 197.600 4.970 200.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 197.600 7.270 200.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.830 197.600 9.110 200.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 197.600 10.950 200.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 197.600 13.250 200.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.810 197.600 15.090 200.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 197.600 16.930 200.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 197.600 19.230 200.000 ;
    END
  END chany_top_out[9]
  PIN left_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.400 167.240 ;
    END
  END left_grid_pin_0_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 49.680 80.000 50.280 ;
    END
  END prog_clk
  PIN right_grid_pin_52_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 149.640 80.000 150.240 ;
    END
  END right_grid_pin_52_
  PIN vpwr
    USE POWER ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 0.990 2.760 79.050 189.000 ;
      LAYER met2 ;
        RECT 1.570 197.320 2.570 197.610 ;
        RECT 3.410 197.320 4.410 197.610 ;
        RECT 5.250 197.320 6.710 197.610 ;
        RECT 7.550 197.320 8.550 197.610 ;
        RECT 9.390 197.320 10.390 197.610 ;
        RECT 11.230 197.320 12.690 197.610 ;
        RECT 13.530 197.320 14.530 197.610 ;
        RECT 15.370 197.320 16.370 197.610 ;
        RECT 17.210 197.320 18.670 197.610 ;
        RECT 19.510 197.320 20.510 197.610 ;
        RECT 21.350 197.320 22.350 197.610 ;
        RECT 23.190 197.320 24.650 197.610 ;
        RECT 25.490 197.320 26.490 197.610 ;
        RECT 27.330 197.320 28.330 197.610 ;
        RECT 29.170 197.320 30.630 197.610 ;
        RECT 31.470 197.320 32.470 197.610 ;
        RECT 33.310 197.320 34.310 197.610 ;
        RECT 35.150 197.320 36.610 197.610 ;
        RECT 37.450 197.320 38.450 197.610 ;
        RECT 39.290 197.320 40.750 197.610 ;
        RECT 41.590 197.320 42.590 197.610 ;
        RECT 43.430 197.320 44.430 197.610 ;
        RECT 45.270 197.320 46.730 197.610 ;
        RECT 47.570 197.320 48.570 197.610 ;
        RECT 49.410 197.320 50.410 197.610 ;
        RECT 51.250 197.320 52.710 197.610 ;
        RECT 53.550 197.320 54.550 197.610 ;
        RECT 55.390 197.320 56.390 197.610 ;
        RECT 57.230 197.320 58.690 197.610 ;
        RECT 59.530 197.320 60.530 197.610 ;
        RECT 61.370 197.320 62.370 197.610 ;
        RECT 63.210 197.320 64.670 197.610 ;
        RECT 65.510 197.320 66.510 197.610 ;
        RECT 67.350 197.320 68.350 197.610 ;
        RECT 69.190 197.320 70.650 197.610 ;
        RECT 71.490 197.320 72.490 197.610 ;
        RECT 73.330 197.320 74.330 197.610 ;
        RECT 75.170 197.320 76.630 197.610 ;
        RECT 77.470 197.320 78.470 197.610 ;
        RECT 1.010 2.680 79.030 197.320 ;
        RECT 1.570 2.400 2.570 2.680 ;
        RECT 3.410 2.400 4.410 2.680 ;
        RECT 5.250 2.400 6.710 2.680 ;
        RECT 7.550 2.400 8.550 2.680 ;
        RECT 9.390 2.400 10.390 2.680 ;
        RECT 11.230 2.400 12.690 2.680 ;
        RECT 13.530 2.400 14.530 2.680 ;
        RECT 15.370 2.400 16.370 2.680 ;
        RECT 17.210 2.400 18.670 2.680 ;
        RECT 19.510 2.400 20.510 2.680 ;
        RECT 21.350 2.400 22.350 2.680 ;
        RECT 23.190 2.400 24.650 2.680 ;
        RECT 25.490 2.400 26.490 2.680 ;
        RECT 27.330 2.400 28.330 2.680 ;
        RECT 29.170 2.400 30.630 2.680 ;
        RECT 31.470 2.400 32.470 2.680 ;
        RECT 33.310 2.400 34.310 2.680 ;
        RECT 35.150 2.400 36.610 2.680 ;
        RECT 37.450 2.400 38.450 2.680 ;
        RECT 39.290 2.400 40.750 2.680 ;
        RECT 41.590 2.400 42.590 2.680 ;
        RECT 43.430 2.400 44.430 2.680 ;
        RECT 45.270 2.400 46.730 2.680 ;
        RECT 47.570 2.400 48.570 2.680 ;
        RECT 49.410 2.400 50.410 2.680 ;
        RECT 51.250 2.400 52.710 2.680 ;
        RECT 53.550 2.400 54.550 2.680 ;
        RECT 55.390 2.400 56.390 2.680 ;
        RECT 57.230 2.400 58.690 2.680 ;
        RECT 59.530 2.400 60.530 2.680 ;
        RECT 61.370 2.400 62.370 2.680 ;
        RECT 63.210 2.400 64.670 2.680 ;
        RECT 65.510 2.400 66.510 2.680 ;
        RECT 67.350 2.400 68.350 2.680 ;
        RECT 69.190 2.400 70.650 2.680 ;
        RECT 71.490 2.400 72.490 2.680 ;
        RECT 73.330 2.400 74.330 2.680 ;
        RECT 75.170 2.400 76.630 2.680 ;
        RECT 77.470 2.400 78.470 2.680 ;
      LAYER met3 ;
        RECT 0.985 167.640 79.055 187.845 ;
        RECT 2.800 166.240 79.055 167.640 ;
        RECT 0.985 150.640 79.055 166.240 ;
        RECT 0.985 149.240 77.200 150.640 ;
        RECT 0.985 101.000 79.055 149.240 ;
        RECT 2.800 99.600 79.055 101.000 ;
        RECT 0.985 50.680 79.055 99.600 ;
        RECT 0.985 49.280 77.200 50.680 ;
        RECT 0.985 34.360 79.055 49.280 ;
        RECT 2.800 32.960 79.055 34.360 ;
        RECT 0.985 6.975 79.055 32.960 ;
      LAYER met4 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END cby_0__1_
END LIBRARY

