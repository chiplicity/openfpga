magic
tech sky130A
magscale 1 2
timestamp 1609024303
<< locali >>
rect 22017 18343 22051 19261
rect 12541 17663 12575 17765
rect 22017 16779 22051 17765
rect 9505 15555 9539 15657
rect 9229 14943 9263 15113
rect 17877 14943 17911 15113
rect 12725 12631 12759 12869
rect 14565 12767 14599 12869
rect 9873 12223 9907 12325
rect 13093 11679 13127 11849
rect 5365 9911 5399 10217
rect 9873 9367 9907 9469
rect 9505 7803 9539 8041
<< viali >>
rect 17693 20553 17727 20587
rect 19441 20553 19475 20587
rect 8769 20485 8803 20519
rect 17325 20485 17359 20519
rect 9413 20417 9447 20451
rect 2145 20349 2179 20383
rect 17141 20349 17175 20383
rect 17509 20349 17543 20383
rect 19165 20349 19199 20383
rect 19257 20349 19291 20383
rect 9137 20281 9171 20315
rect 1501 20213 1535 20247
rect 2329 20213 2363 20247
rect 9229 20213 9263 20247
rect 20361 20213 20395 20247
rect 20821 20213 20855 20247
rect 2053 20009 2087 20043
rect 8769 20009 8803 20043
rect 11529 20009 11563 20043
rect 13093 20009 13127 20043
rect 13461 20009 13495 20043
rect 14013 20009 14047 20043
rect 14565 20009 14599 20043
rect 15485 20009 15519 20043
rect 16865 20009 16899 20043
rect 17233 20009 17267 20043
rect 18429 20009 18463 20043
rect 21465 20009 21499 20043
rect 3249 19941 3283 19975
rect 10118 19941 10152 19975
rect 11897 19941 11931 19975
rect 13921 19941 13955 19975
rect 14749 19941 14783 19975
rect 16405 19941 16439 19975
rect 20085 19941 20119 19975
rect 1501 19873 1535 19907
rect 1869 19873 1903 19907
rect 2237 19873 2271 19907
rect 2593 19873 2627 19907
rect 9137 19873 9171 19907
rect 9689 19873 9723 19907
rect 12357 19873 12391 19907
rect 12633 19873 12667 19907
rect 12909 19873 12943 19907
rect 14381 19873 14415 19907
rect 15301 19873 15335 19907
rect 16129 19873 16163 19907
rect 16681 19873 16715 19907
rect 17049 19873 17083 19907
rect 17601 19873 17635 19907
rect 17877 19873 17911 19907
rect 18245 19873 18279 19907
rect 18613 19873 18647 19907
rect 19349 19873 19383 19907
rect 19441 19873 19475 19907
rect 19809 19873 19843 19907
rect 20453 19873 20487 19907
rect 20913 19873 20947 19907
rect 21281 19873 21315 19907
rect 3065 19805 3099 19839
rect 9229 19805 9263 19839
rect 9413 19805 9447 19839
rect 9873 19805 9907 19839
rect 11989 19805 12023 19839
rect 12081 19805 12115 19839
rect 14105 19805 14139 19839
rect 19533 19805 19567 19839
rect 13553 19737 13587 19771
rect 18797 19737 18831 19771
rect 18981 19737 19015 19771
rect 21097 19737 21131 19771
rect 1685 19669 1719 19703
rect 2421 19669 2455 19703
rect 2789 19669 2823 19703
rect 8585 19669 8619 19703
rect 11253 19669 11287 19703
rect 15025 19669 15059 19703
rect 20637 19669 20671 19703
rect 3157 19465 3191 19499
rect 3617 19465 3651 19499
rect 6377 19465 6411 19499
rect 9045 19465 9079 19499
rect 10517 19465 10551 19499
rect 15669 19465 15703 19499
rect 18061 19465 18095 19499
rect 20637 19465 20671 19499
rect 21005 19465 21039 19499
rect 21373 19465 21407 19499
rect 14013 19397 14047 19431
rect 14565 19329 14599 19363
rect 15393 19329 15427 19363
rect 16221 19329 16255 19363
rect 16773 19329 16807 19363
rect 18613 19329 18647 19363
rect 1501 19261 1535 19295
rect 1869 19261 1903 19295
rect 2237 19261 2271 19295
rect 2605 19261 2639 19295
rect 2973 19261 3007 19295
rect 3433 19261 3467 19295
rect 3985 19261 4019 19295
rect 4997 19261 5031 19295
rect 6193 19261 6227 19295
rect 7665 19261 7699 19295
rect 9137 19261 9171 19295
rect 9404 19261 9438 19295
rect 10885 19261 10919 19295
rect 12541 19261 12575 19295
rect 12797 19261 12831 19295
rect 16497 19261 16531 19295
rect 17049 19261 17083 19295
rect 17417 19261 17451 19295
rect 18981 19261 19015 19295
rect 20453 19261 20487 19295
rect 20821 19261 20855 19295
rect 21189 19261 21223 19295
rect 22017 19261 22051 19295
rect 4721 19193 4755 19227
rect 7932 19193 7966 19227
rect 11152 19193 11186 19227
rect 15301 19193 15335 19227
rect 18521 19193 18555 19227
rect 19248 19193 19282 19227
rect 1685 19125 1719 19159
rect 2053 19125 2087 19159
rect 2421 19125 2455 19159
rect 2789 19125 2823 19159
rect 10609 19125 10643 19159
rect 12265 19125 12299 19159
rect 13921 19125 13955 19159
rect 14381 19125 14415 19159
rect 14473 19125 14507 19159
rect 14841 19125 14875 19159
rect 15209 19125 15243 19159
rect 16037 19125 16071 19159
rect 16129 19125 16163 19159
rect 17233 19125 17267 19159
rect 17601 19125 17635 19159
rect 18429 19125 18463 19159
rect 20361 19125 20395 19159
rect 1593 18921 1627 18955
rect 1961 18921 1995 18955
rect 2329 18921 2363 18955
rect 3433 18921 3467 18955
rect 8769 18921 8803 18955
rect 9137 18921 9171 18955
rect 11161 18921 11195 18955
rect 11713 18921 11747 18955
rect 13369 18921 13403 18955
rect 15301 18921 15335 18955
rect 18245 18921 18279 18955
rect 19809 18921 19843 18955
rect 21097 18921 21131 18955
rect 21465 18921 21499 18955
rect 6837 18853 6871 18887
rect 11621 18853 11655 18887
rect 13912 18853 13946 18887
rect 15761 18853 15795 18887
rect 16405 18853 16439 18887
rect 18604 18853 18638 18887
rect 20269 18853 20303 18887
rect 1777 18785 1811 18819
rect 2145 18785 2179 18819
rect 2513 18785 2547 18819
rect 6009 18785 6043 18819
rect 6561 18785 6595 18819
rect 8401 18785 8435 18819
rect 9689 18785 9723 18819
rect 11069 18785 11103 18819
rect 12081 18785 12115 18819
rect 12909 18785 12943 18819
rect 13645 18785 13679 18819
rect 15669 18785 15703 18819
rect 16129 18785 16163 18819
rect 17132 18785 17166 18819
rect 20177 18785 20211 18819
rect 20913 18785 20947 18819
rect 21281 18785 21315 18819
rect 2973 18717 3007 18751
rect 9229 18717 9263 18751
rect 9413 18717 9447 18751
rect 9965 18717 9999 18751
rect 11345 18717 11379 18751
rect 12173 18717 12207 18751
rect 12357 18717 12391 18751
rect 13001 18717 13035 18751
rect 13093 18717 13127 18751
rect 15853 18717 15887 18751
rect 16865 18717 16899 18751
rect 18337 18717 18371 18751
rect 20361 18717 20395 18751
rect 2697 18649 2731 18683
rect 3065 18649 3099 18683
rect 3893 18649 3927 18683
rect 8309 18649 8343 18683
rect 10701 18649 10735 18683
rect 12541 18649 12575 18683
rect 15025 18649 15059 18683
rect 19717 18649 19751 18683
rect 1501 18581 1535 18615
rect 6193 18581 6227 18615
rect 8585 18581 8619 18615
rect 16773 18581 16807 18615
rect 20729 18581 20763 18615
rect 1961 18377 1995 18411
rect 13921 18377 13955 18411
rect 14473 18377 14507 18411
rect 16037 18377 16071 18411
rect 17509 18377 17543 18411
rect 18061 18377 18095 18411
rect 19257 18377 19291 18411
rect 19533 18377 19567 18411
rect 21005 18377 21039 18411
rect 12081 18309 12115 18343
rect 21189 18309 21223 18343
rect 22017 18309 22051 18343
rect 5457 18241 5491 18275
rect 7849 18241 7883 18275
rect 8401 18241 8435 18275
rect 12449 18241 12483 18275
rect 18613 18241 18647 18275
rect 20085 18241 20119 18275
rect 1777 18173 1811 18207
rect 5181 18173 5215 18207
rect 8125 18173 8159 18207
rect 10701 18173 10735 18207
rect 10968 18173 11002 18207
rect 14657 18173 14691 18207
rect 14924 18173 14958 18207
rect 16129 18173 16163 18207
rect 16385 18173 16419 18207
rect 20821 18173 20855 18207
rect 12173 18105 12207 18139
rect 17601 18105 17635 18139
rect 18429 18105 18463 18139
rect 19901 18105 19935 18139
rect 20361 18105 20395 18139
rect 21373 18105 21407 18139
rect 2237 18037 2271 18071
rect 2605 18037 2639 18071
rect 7297 18037 7331 18071
rect 7665 18037 7699 18071
rect 7757 18037 7791 18071
rect 18521 18037 18555 18071
rect 19441 18037 19475 18071
rect 19993 18037 20027 18071
rect 20729 18037 20763 18071
rect 4353 17833 4387 17867
rect 6745 17833 6779 17867
rect 7205 17833 7239 17867
rect 7573 17833 7607 17867
rect 8401 17833 8435 17867
rect 8677 17833 8711 17867
rect 9321 17833 9355 17867
rect 11253 17833 11287 17867
rect 13001 17833 13035 17867
rect 15301 17833 15335 17867
rect 15761 17833 15795 17867
rect 16957 17833 16991 17867
rect 21097 17833 21131 17867
rect 2605 17765 2639 17799
rect 4721 17765 4755 17799
rect 8033 17765 8067 17799
rect 8769 17765 8803 17799
rect 11713 17765 11747 17799
rect 12541 17765 12575 17799
rect 15117 17765 15151 17799
rect 17325 17765 17359 17799
rect 20085 17765 20119 17799
rect 22017 17765 22051 17799
rect 2329 17697 2363 17731
rect 5448 17697 5482 17731
rect 7113 17697 7147 17731
rect 7941 17697 7975 17731
rect 8953 17697 8987 17731
rect 10048 17697 10082 17731
rect 11621 17697 11655 17731
rect 12081 17697 12115 17731
rect 15669 17697 15703 17731
rect 16129 17697 16163 17731
rect 19625 17697 19659 17731
rect 20177 17697 20211 17731
rect 20913 17697 20947 17731
rect 21465 17697 21499 17731
rect 4813 17629 4847 17663
rect 4905 17629 4939 17663
rect 5181 17629 5215 17663
rect 7389 17629 7423 17663
rect 8125 17629 8159 17663
rect 9781 17629 9815 17663
rect 11805 17629 11839 17663
rect 12449 17629 12483 17663
rect 12541 17629 12575 17663
rect 15853 17629 15887 17663
rect 17417 17629 17451 17663
rect 17509 17629 17543 17663
rect 20361 17629 20395 17663
rect 11161 17561 11195 17595
rect 16773 17561 16807 17595
rect 18061 17561 18095 17595
rect 6561 17493 6595 17527
rect 9137 17493 9171 17527
rect 12817 17493 12851 17527
rect 17877 17493 17911 17527
rect 19717 17493 19751 17527
rect 20637 17493 20671 17527
rect 21281 17493 21315 17527
rect 1961 17289 1995 17323
rect 2329 17289 2363 17323
rect 6009 17289 6043 17323
rect 8309 17289 8343 17323
rect 8401 17289 8435 17323
rect 10333 17289 10367 17323
rect 12173 17289 12207 17323
rect 20545 17289 20579 17323
rect 21005 17289 21039 17323
rect 4537 17221 4571 17255
rect 2697 17153 2731 17187
rect 8953 17153 8987 17187
rect 10057 17153 10091 17187
rect 10885 17153 10919 17187
rect 11713 17153 11747 17187
rect 12817 17153 12851 17187
rect 13645 17153 13679 17187
rect 14565 17153 14599 17187
rect 14749 17153 14783 17187
rect 15209 17153 15243 17187
rect 17417 17153 17451 17187
rect 1777 17085 1811 17119
rect 2145 17085 2179 17119
rect 3157 17085 3191 17119
rect 4629 17085 4663 17119
rect 6929 17085 6963 17119
rect 9321 17085 9355 17119
rect 10793 17085 10827 17119
rect 12541 17085 12575 17119
rect 14933 17085 14967 17119
rect 17233 17085 17267 17119
rect 19165 17085 19199 17119
rect 20729 17085 20763 17119
rect 20821 17085 20855 17119
rect 3424 17017 3458 17051
rect 4874 17017 4908 17051
rect 7196 17017 7230 17051
rect 8861 17017 8895 17051
rect 11529 17017 11563 17051
rect 13461 17017 13495 17051
rect 19410 17017 19444 17051
rect 21373 17017 21407 17051
rect 2605 16949 2639 16983
rect 8769 16949 8803 16983
rect 9505 16949 9539 16983
rect 9873 16949 9907 16983
rect 9965 16949 9999 16983
rect 10701 16949 10735 16983
rect 11161 16949 11195 16983
rect 11621 16949 11655 16983
rect 12081 16949 12115 16983
rect 13093 16949 13127 16983
rect 13553 16949 13587 16983
rect 14105 16949 14139 16983
rect 14473 16949 14507 16983
rect 15577 16949 15611 16983
rect 21189 16949 21223 16983
rect 2789 16745 2823 16779
rect 3065 16745 3099 16779
rect 4537 16745 4571 16779
rect 5365 16745 5399 16779
rect 5917 16745 5951 16779
rect 7573 16745 7607 16779
rect 12909 16745 12943 16779
rect 14197 16745 14231 16779
rect 15761 16745 15795 16779
rect 18521 16745 18555 16779
rect 18889 16745 18923 16779
rect 21097 16745 21131 16779
rect 21281 16745 21315 16779
rect 22017 16745 22051 16779
rect 8370 16677 8404 16711
rect 9689 16677 9723 16711
rect 10425 16677 10459 16711
rect 13277 16677 13311 16711
rect 13369 16677 13403 16711
rect 16589 16677 16623 16711
rect 3433 16609 3467 16643
rect 4445 16609 4479 16643
rect 5273 16609 5307 16643
rect 5825 16609 5859 16643
rect 6193 16609 6227 16643
rect 6460 16609 6494 16643
rect 8125 16609 8159 16643
rect 11704 16609 11738 16643
rect 14105 16609 14139 16643
rect 14749 16609 14783 16643
rect 14933 16609 14967 16643
rect 15669 16609 15703 16643
rect 16313 16609 16347 16643
rect 17132 16609 17166 16643
rect 18981 16609 19015 16643
rect 19349 16609 19383 16643
rect 19616 16609 19650 16643
rect 20913 16609 20947 16643
rect 2881 16541 2915 16575
rect 3525 16541 3559 16575
rect 3709 16541 3743 16575
rect 4629 16541 4663 16575
rect 5457 16541 5491 16575
rect 9873 16541 9907 16575
rect 10517 16541 10551 16575
rect 10609 16541 10643 16575
rect 11437 16541 11471 16575
rect 13553 16541 13587 16575
rect 14289 16541 14323 16575
rect 15853 16541 15887 16575
rect 16865 16541 16899 16575
rect 19165 16541 19199 16575
rect 9505 16473 9539 16507
rect 12817 16473 12851 16507
rect 13737 16473 13771 16507
rect 2237 16405 2271 16439
rect 4077 16405 4111 16439
rect 4905 16405 4939 16439
rect 10057 16405 10091 16439
rect 14565 16405 14599 16439
rect 15301 16405 15335 16439
rect 18245 16405 18279 16439
rect 20729 16405 20763 16439
rect 1961 16201 1995 16235
rect 2329 16201 2363 16235
rect 3985 16201 4019 16235
rect 4261 16201 4295 16235
rect 5089 16201 5123 16235
rect 6837 16201 6871 16235
rect 9321 16201 9355 16235
rect 11529 16201 11563 16235
rect 12173 16201 12207 16235
rect 15301 16201 15335 16235
rect 16773 16201 16807 16235
rect 18337 16201 18371 16235
rect 20269 16201 20303 16235
rect 21281 16201 21315 16235
rect 4169 16133 4203 16167
rect 16865 16133 16899 16167
rect 20177 16133 20211 16167
rect 4721 16065 4755 16099
rect 4813 16065 4847 16099
rect 5641 16065 5675 16099
rect 7481 16065 7515 16099
rect 8309 16065 8343 16099
rect 9965 16065 9999 16099
rect 17417 16065 17451 16099
rect 20821 16065 20855 16099
rect 1777 15997 1811 16031
rect 2145 15997 2179 16031
rect 2605 15997 2639 16031
rect 4629 15997 4663 16031
rect 8769 15997 8803 16031
rect 9689 15997 9723 16031
rect 9781 15997 9815 16031
rect 10149 15997 10183 16031
rect 12449 15997 12483 16031
rect 12716 15997 12750 16031
rect 13921 15997 13955 16031
rect 15393 15997 15427 16031
rect 15649 15997 15683 16031
rect 17325 15997 17359 16031
rect 18797 15997 18831 16031
rect 21097 15997 21131 16031
rect 2872 15929 2906 15963
rect 5549 15929 5583 15963
rect 7205 15929 7239 15963
rect 8033 15929 8067 15963
rect 10416 15929 10450 15963
rect 14188 15929 14222 15963
rect 18061 15929 18095 15963
rect 19064 15929 19098 15963
rect 20729 15929 20763 15963
rect 5457 15861 5491 15895
rect 7297 15861 7331 15895
rect 7665 15861 7699 15895
rect 8125 15861 8159 15895
rect 8585 15861 8619 15895
rect 11621 15861 11655 15895
rect 13829 15861 13863 15895
rect 17233 15861 17267 15895
rect 17693 15861 17727 15895
rect 20637 15861 20671 15895
rect 21465 15861 21499 15895
rect 1961 15657 1995 15691
rect 2329 15657 2363 15691
rect 5181 15657 5215 15691
rect 6009 15657 6043 15691
rect 7941 15657 7975 15691
rect 8309 15657 8343 15691
rect 9229 15657 9263 15691
rect 9505 15657 9539 15691
rect 11161 15657 11195 15691
rect 12357 15657 12391 15691
rect 14197 15657 14231 15691
rect 14657 15657 14691 15691
rect 15301 15657 15335 15691
rect 17509 15657 17543 15691
rect 19165 15657 19199 15691
rect 19257 15657 19291 15691
rect 20637 15657 20671 15691
rect 21097 15657 21131 15691
rect 21465 15657 21499 15691
rect 2605 15589 2639 15623
rect 4077 15589 4111 15623
rect 5549 15589 5583 15623
rect 11529 15589 11563 15623
rect 12449 15589 12483 15623
rect 14565 15589 14599 15623
rect 15761 15589 15795 15623
rect 16396 15589 16430 15623
rect 18052 15589 18086 15623
rect 1777 15521 1811 15555
rect 2145 15521 2179 15555
rect 2697 15521 2731 15555
rect 4721 15521 4755 15555
rect 5641 15521 5675 15555
rect 6193 15521 6227 15555
rect 7573 15521 7607 15555
rect 9505 15521 9539 15555
rect 9956 15521 9990 15555
rect 15669 15521 15703 15555
rect 19625 15521 19659 15555
rect 20453 15521 20487 15555
rect 20913 15521 20947 15555
rect 21281 15521 21315 15555
rect 4813 15453 4847 15487
rect 4997 15453 5031 15487
rect 5825 15453 5859 15487
rect 6837 15453 6871 15487
rect 8401 15453 8435 15487
rect 8493 15453 8527 15487
rect 8769 15453 8803 15487
rect 9689 15453 9723 15487
rect 11621 15453 11655 15487
rect 11713 15453 11747 15487
rect 12541 15453 12575 15487
rect 14749 15453 14783 15487
rect 15853 15453 15887 15487
rect 16129 15453 16163 15487
rect 17785 15453 17819 15487
rect 19717 15453 19751 15487
rect 19809 15453 19843 15487
rect 7389 15385 7423 15419
rect 7757 15385 7791 15419
rect 11989 15385 12023 15419
rect 20085 15385 20119 15419
rect 4353 15317 4387 15351
rect 7021 15317 7055 15351
rect 9045 15317 9079 15351
rect 11069 15317 11103 15351
rect 12909 15317 12943 15351
rect 17693 15317 17727 15351
rect 20269 15317 20303 15351
rect 1961 15113 1995 15147
rect 3065 15113 3099 15147
rect 5641 15113 5675 15147
rect 7665 15113 7699 15147
rect 8677 15113 8711 15147
rect 9229 15113 9263 15147
rect 9413 15113 9447 15147
rect 10885 15113 10919 15147
rect 12265 15113 12299 15147
rect 15761 15113 15795 15147
rect 16221 15113 16255 15147
rect 17877 15113 17911 15147
rect 19073 15113 19107 15147
rect 21373 15113 21407 15147
rect 2329 14977 2363 15011
rect 3709 14977 3743 15011
rect 4261 14977 4295 15011
rect 6561 14977 6595 15011
rect 7389 14977 7423 15011
rect 8309 14977 8343 15011
rect 8585 14977 8619 15011
rect 9597 15045 9631 15079
rect 12449 15045 12483 15079
rect 11437 14977 11471 15011
rect 11713 14977 11747 15011
rect 12909 14977 12943 15011
rect 13093 14977 13127 15011
rect 16865 14977 16899 15011
rect 17509 14977 17543 15011
rect 17601 14977 17635 15011
rect 18613 14977 18647 15011
rect 20361 14977 20395 15011
rect 20913 14977 20947 15011
rect 1777 14909 1811 14943
rect 2145 14909 2179 14943
rect 4528 14909 4562 14943
rect 6285 14909 6319 14943
rect 9229 14909 9263 14943
rect 11253 14909 11287 14943
rect 12817 14909 12851 14943
rect 13277 14909 13311 14943
rect 13737 14909 13771 14943
rect 13829 14909 13863 14943
rect 16129 14909 16163 14943
rect 17417 14909 17451 14943
rect 17877 14909 17911 14943
rect 18429 14909 18463 14943
rect 18981 14909 19015 14943
rect 20085 14909 20119 14943
rect 20637 14909 20671 14943
rect 21189 14909 21223 14943
rect 2973 14841 3007 14875
rect 3433 14841 3467 14875
rect 5825 14841 5859 14875
rect 6377 14841 6411 14875
rect 7205 14841 7239 14875
rect 14096 14841 14130 14875
rect 16589 14841 16623 14875
rect 18521 14841 18555 14875
rect 2789 14773 2823 14807
rect 3525 14773 3559 14807
rect 3985 14773 4019 14807
rect 5917 14773 5951 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 8033 14773 8067 14807
rect 8125 14773 8159 14807
rect 11345 14773 11379 14807
rect 11989 14773 12023 14807
rect 13553 14773 13587 14807
rect 15209 14773 15243 14807
rect 15945 14773 15979 14807
rect 16681 14773 16715 14807
rect 17049 14773 17083 14807
rect 18061 14773 18095 14807
rect 1961 14569 1995 14603
rect 2329 14569 2363 14603
rect 8769 14569 8803 14603
rect 9229 14569 9263 14603
rect 9689 14569 9723 14603
rect 10149 14569 10183 14603
rect 12265 14569 12299 14603
rect 14197 14569 14231 14603
rect 14381 14569 14415 14603
rect 19809 14569 19843 14603
rect 19901 14569 19935 14603
rect 21097 14569 21131 14603
rect 5794 14501 5828 14535
rect 7564 14501 7598 14535
rect 16948 14501 16982 14535
rect 1777 14433 1811 14467
rect 2145 14433 2179 14467
rect 4077 14433 4111 14467
rect 4344 14433 4378 14467
rect 9137 14433 9171 14467
rect 10057 14433 10091 14467
rect 12992 14433 13026 14467
rect 14749 14433 14783 14467
rect 16037 14433 16071 14467
rect 16681 14433 16715 14467
rect 18429 14433 18463 14467
rect 18696 14433 18730 14467
rect 20269 14433 20303 14467
rect 20913 14433 20947 14467
rect 5549 14365 5583 14399
rect 7297 14365 7331 14399
rect 9321 14365 9355 14399
rect 10333 14365 10367 14399
rect 12357 14365 12391 14399
rect 12449 14365 12483 14399
rect 12725 14365 12759 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 16129 14365 16163 14399
rect 16313 14365 16347 14399
rect 18245 14365 18279 14399
rect 20361 14365 20395 14399
rect 20453 14365 20487 14399
rect 6929 14297 6963 14331
rect 8677 14297 8711 14331
rect 5457 14229 5491 14263
rect 11897 14229 11931 14263
rect 14105 14229 14139 14263
rect 15485 14229 15519 14263
rect 15669 14229 15703 14263
rect 18061 14229 18095 14263
rect 21281 14229 21315 14263
rect 3525 14025 3559 14059
rect 5181 14025 5215 14059
rect 8769 14025 8803 14059
rect 8953 14025 8987 14059
rect 9137 14025 9171 14059
rect 10057 14025 10091 14059
rect 14473 14025 14507 14059
rect 14933 14025 14967 14059
rect 19533 14025 19567 14059
rect 21097 14025 21131 14059
rect 12817 13957 12851 13991
rect 19441 13957 19475 13991
rect 1869 13889 1903 13923
rect 2329 13889 2363 13923
rect 4169 13889 4203 13923
rect 4997 13889 5031 13923
rect 5641 13889 5675 13923
rect 5733 13889 5767 13923
rect 9781 13889 9815 13923
rect 10517 13889 10551 13923
rect 10701 13889 10735 13923
rect 13277 13889 13311 13923
rect 13369 13889 13403 13923
rect 14289 13889 14323 13923
rect 15485 13889 15519 13923
rect 16313 13889 16347 13923
rect 19993 13889 20027 13923
rect 20085 13889 20119 13923
rect 1593 13821 1627 13855
rect 2145 13821 2179 13855
rect 3985 13821 4019 13855
rect 5549 13821 5583 13855
rect 7389 13821 7423 13855
rect 7656 13821 7690 13855
rect 9505 13821 9539 13855
rect 9597 13821 9631 13855
rect 10885 13821 10919 13855
rect 14841 13821 14875 13855
rect 15301 13821 15335 13855
rect 18061 13821 18095 13855
rect 20361 13821 20395 13855
rect 20637 13821 20671 13855
rect 20913 13821 20947 13855
rect 3893 13753 3927 13787
rect 4721 13753 4755 13787
rect 11152 13753 11186 13787
rect 13185 13753 13219 13787
rect 14013 13753 14047 13787
rect 14105 13753 14139 13787
rect 16129 13753 16163 13787
rect 16589 13753 16623 13787
rect 18328 13753 18362 13787
rect 4353 13685 4387 13719
rect 4813 13685 4847 13719
rect 6929 13685 6963 13719
rect 10425 13685 10459 13719
rect 12265 13685 12299 13719
rect 13645 13685 13679 13719
rect 15393 13685 15427 13719
rect 15761 13685 15795 13719
rect 16221 13685 16255 13719
rect 16957 13685 16991 13719
rect 19901 13685 19935 13719
rect 3709 13481 3743 13515
rect 4629 13481 4663 13515
rect 5457 13481 5491 13515
rect 6009 13481 6043 13515
rect 7205 13481 7239 13515
rect 7297 13481 7331 13515
rect 7665 13481 7699 13515
rect 8769 13481 8803 13515
rect 9781 13481 9815 13515
rect 10241 13481 10275 13515
rect 14197 13481 14231 13515
rect 19533 13481 19567 13515
rect 19993 13481 20027 13515
rect 20453 13481 20487 13515
rect 4261 13413 4295 13447
rect 5089 13413 5123 13447
rect 5733 13413 5767 13447
rect 8033 13413 8067 13447
rect 10057 13413 10091 13447
rect 10517 13413 10551 13447
rect 14657 13413 14691 13447
rect 15546 13413 15580 13447
rect 21189 13413 21223 13447
rect 2596 13345 2630 13379
rect 4997 13345 5031 13379
rect 6377 13345 6411 13379
rect 8677 13345 8711 13379
rect 12624 13345 12658 13379
rect 17132 13345 17166 13379
rect 20361 13345 20395 13379
rect 20913 13345 20947 13379
rect 2329 13277 2363 13311
rect 5273 13277 5307 13311
rect 6469 13277 6503 13311
rect 6653 13277 6687 13311
rect 7389 13277 7423 13311
rect 8125 13277 8159 13311
rect 8217 13277 8251 13311
rect 12357 13277 12391 13311
rect 14289 13277 14323 13311
rect 14381 13277 14415 13311
rect 15301 13277 15335 13311
rect 16865 13277 16899 13311
rect 18981 13277 19015 13311
rect 19625 13277 19659 13311
rect 19809 13277 19843 13311
rect 20545 13277 20579 13311
rect 6837 13209 6871 13243
rect 11805 13209 11839 13243
rect 19165 13209 19199 13243
rect 4445 13141 4479 13175
rect 8493 13141 8527 13175
rect 13737 13141 13771 13175
rect 13829 13141 13863 13175
rect 16681 13141 16715 13175
rect 18245 13141 18279 13175
rect 1409 12937 1443 12971
rect 3893 12937 3927 12971
rect 11345 12937 11379 12971
rect 12449 12937 12483 12971
rect 13461 12937 13495 12971
rect 19073 12937 19107 12971
rect 19257 12937 19291 12971
rect 20085 12937 20119 12971
rect 5917 12869 5951 12903
rect 9873 12869 9907 12903
rect 12725 12869 12759 12903
rect 12817 12869 12851 12903
rect 14565 12869 14599 12903
rect 18061 12869 18095 12903
rect 2053 12801 2087 12835
rect 2789 12801 2823 12835
rect 4077 12801 4111 12835
rect 5365 12801 5399 12835
rect 6469 12801 6503 12835
rect 8309 12801 8343 12835
rect 11897 12801 11931 12835
rect 12081 12801 12115 12835
rect 6837 12733 6871 12767
rect 8493 12733 8527 12767
rect 9965 12733 9999 12767
rect 2605 12665 2639 12699
rect 5273 12665 5307 12699
rect 7082 12665 7116 12699
rect 8760 12665 8794 12699
rect 10232 12665 10266 12699
rect 14013 12801 14047 12835
rect 15393 12801 15427 12835
rect 18613 12801 18647 12835
rect 19809 12801 19843 12835
rect 20637 12801 20671 12835
rect 20913 12801 20947 12835
rect 13001 12733 13035 12767
rect 13829 12733 13863 12767
rect 14473 12733 14507 12767
rect 14565 12733 14599 12767
rect 15301 12733 15335 12767
rect 19625 12733 19659 12767
rect 13921 12665 13955 12699
rect 14657 12665 14691 12699
rect 15209 12665 15243 12699
rect 15669 12665 15703 12699
rect 20453 12665 20487 12699
rect 21373 12665 21407 12699
rect 1777 12597 1811 12631
rect 1869 12597 1903 12631
rect 2237 12597 2271 12631
rect 2697 12597 2731 12631
rect 4813 12597 4847 12631
rect 5181 12597 5215 12631
rect 8217 12597 8251 12631
rect 11437 12597 11471 12631
rect 11805 12597 11839 12631
rect 12725 12597 12759 12631
rect 14289 12597 14323 12631
rect 14841 12597 14875 12631
rect 18429 12597 18463 12631
rect 18521 12597 18555 12631
rect 19717 12597 19751 12631
rect 20545 12597 20579 12631
rect 21189 12597 21223 12631
rect 2973 12393 3007 12427
rect 3065 12393 3099 12427
rect 3433 12393 3467 12427
rect 4537 12393 4571 12427
rect 7757 12393 7791 12427
rect 14013 12393 14047 12427
rect 14381 12393 14415 12427
rect 16589 12393 16623 12427
rect 18061 12393 18095 12427
rect 18521 12393 18555 12427
rect 19349 12393 19383 12427
rect 19717 12393 19751 12427
rect 20177 12393 20211 12427
rect 3525 12325 3559 12359
rect 5172 12325 5206 12359
rect 7665 12325 7699 12359
rect 8392 12325 8426 12359
rect 9873 12325 9907 12359
rect 10425 12325 10459 12359
rect 11253 12325 11287 12359
rect 11989 12325 12023 12359
rect 1860 12257 1894 12291
rect 4445 12257 4479 12291
rect 8125 12257 8159 12291
rect 10333 12257 10367 12291
rect 11161 12257 11195 12291
rect 12173 12257 12207 12291
rect 12808 12257 12842 12291
rect 14473 12257 14507 12291
rect 14841 12257 14875 12291
rect 15669 12257 15703 12291
rect 15761 12257 15795 12291
rect 16957 12257 16991 12291
rect 17969 12257 18003 12291
rect 18889 12257 18923 12291
rect 1593 12189 1627 12223
rect 3709 12189 3743 12223
rect 4721 12189 4755 12223
rect 4905 12189 4939 12223
rect 7941 12189 7975 12223
rect 9781 12189 9815 12223
rect 9873 12189 9907 12223
rect 10609 12189 10643 12223
rect 11437 12189 11471 12223
rect 12541 12189 12575 12223
rect 14657 12189 14691 12223
rect 15853 12189 15887 12223
rect 17049 12189 17083 12223
rect 17233 12189 17267 12223
rect 18153 12189 18187 12223
rect 18981 12189 19015 12223
rect 19165 12189 19199 12223
rect 19809 12189 19843 12223
rect 19901 12189 19935 12223
rect 4077 12121 4111 12155
rect 9505 12121 9539 12155
rect 10793 12121 10827 12155
rect 17601 12121 17635 12155
rect 6285 12053 6319 12087
rect 7297 12053 7331 12087
rect 9965 12053 9999 12087
rect 11621 12053 11655 12087
rect 11805 12053 11839 12087
rect 13921 12053 13955 12087
rect 15025 12053 15059 12087
rect 15301 12053 15335 12087
rect 16221 12053 16255 12087
rect 16405 12053 16439 12087
rect 1869 11849 1903 11883
rect 8309 11849 8343 11883
rect 9505 11849 9539 11883
rect 9689 11849 9723 11883
rect 13093 11849 13127 11883
rect 14657 11849 14691 11883
rect 17877 11849 17911 11883
rect 18521 11849 18555 11883
rect 5273 11781 5307 11815
rect 2421 11713 2455 11747
rect 6009 11713 6043 11747
rect 8033 11713 8067 11747
rect 8953 11713 8987 11747
rect 10149 11713 10183 11747
rect 10241 11713 10275 11747
rect 11161 11713 11195 11747
rect 12081 11713 12115 11747
rect 13185 11713 13219 11747
rect 15117 11713 15151 11747
rect 15209 11713 15243 11747
rect 19165 11713 19199 11747
rect 19901 11713 19935 11747
rect 20637 11713 20671 11747
rect 3893 11645 3927 11679
rect 5825 11645 5859 11679
rect 6285 11645 6319 11679
rect 7021 11645 7055 11679
rect 7849 11645 7883 11679
rect 8677 11645 8711 11679
rect 9137 11645 9171 11679
rect 10885 11645 10919 11679
rect 11897 11645 11931 11679
rect 12633 11645 12667 11679
rect 13093 11645 13127 11679
rect 13452 11645 13486 11679
rect 15025 11645 15059 11679
rect 15669 11645 15703 11679
rect 16497 11645 16531 11679
rect 16764 11645 16798 11679
rect 20361 11645 20395 11679
rect 21097 11645 21131 11679
rect 4160 11577 4194 11611
rect 5733 11577 5767 11611
rect 6469 11577 6503 11611
rect 8769 11577 8803 11611
rect 10977 11577 11011 11611
rect 19809 11577 19843 11611
rect 20177 11577 20211 11611
rect 2237 11509 2271 11543
rect 2329 11509 2363 11543
rect 5365 11509 5399 11543
rect 6837 11509 6871 11543
rect 7481 11509 7515 11543
rect 7941 11509 7975 11543
rect 9321 11509 9355 11543
rect 10057 11509 10091 11543
rect 10517 11509 10551 11543
rect 11345 11509 11379 11543
rect 11529 11509 11563 11543
rect 11989 11509 12023 11543
rect 12449 11509 12483 11543
rect 14565 11509 14599 11543
rect 15485 11509 15519 11543
rect 18889 11509 18923 11543
rect 18981 11509 19015 11543
rect 19349 11509 19383 11543
rect 19717 11509 19751 11543
rect 20913 11509 20947 11543
rect 21281 11509 21315 11543
rect 2973 11305 3007 11339
rect 3157 11305 3191 11339
rect 4537 11305 4571 11339
rect 4813 11305 4847 11339
rect 5181 11305 5215 11339
rect 5273 11305 5307 11339
rect 5641 11305 5675 11339
rect 7205 11305 7239 11339
rect 7665 11305 7699 11339
rect 8585 11305 8619 11339
rect 9045 11305 9079 11339
rect 9689 11305 9723 11339
rect 12173 11305 12207 11339
rect 12541 11305 12575 11339
rect 13093 11305 13127 11339
rect 13553 11305 13587 11339
rect 13921 11305 13955 11339
rect 16957 11305 16991 11339
rect 17785 11305 17819 11339
rect 17969 11305 18003 11339
rect 18245 11305 18279 11339
rect 19533 11305 19567 11339
rect 20269 11305 20303 11339
rect 21097 11305 21131 11339
rect 6101 11237 6135 11271
rect 6469 11237 6503 11271
rect 8401 11237 8435 11271
rect 10149 11237 10183 11271
rect 12633 11237 12667 11271
rect 15730 11237 15764 11271
rect 17417 11237 17451 11271
rect 20361 11237 20395 11271
rect 21281 11237 21315 11271
rect 1860 11169 1894 11203
rect 3525 11169 3559 11203
rect 4721 11169 4755 11203
rect 6009 11169 6043 11203
rect 7573 11169 7607 11203
rect 8953 11169 8987 11203
rect 10057 11169 10091 11203
rect 10968 11169 11002 11203
rect 13461 11169 13495 11203
rect 17325 11169 17359 11203
rect 18613 11169 18647 11203
rect 18705 11169 18739 11203
rect 19441 11169 19475 11203
rect 20913 11169 20947 11203
rect 1593 11101 1627 11135
rect 3617 11101 3651 11135
rect 3801 11101 3835 11135
rect 5457 11101 5491 11135
rect 6193 11101 6227 11135
rect 7757 11101 7791 11135
rect 9229 11101 9263 11135
rect 10241 11101 10275 11135
rect 10701 11101 10735 11135
rect 12817 11101 12851 11135
rect 13737 11101 13771 11135
rect 14197 11101 14231 11135
rect 15485 11101 15519 11135
rect 17601 11101 17635 11135
rect 18889 11101 18923 11135
rect 19625 11101 19659 11135
rect 20453 11101 20487 11135
rect 9413 11033 9447 11067
rect 16865 11033 16899 11067
rect 21465 11033 21499 11067
rect 4261 10965 4295 10999
rect 10609 10965 10643 10999
rect 12081 10965 12115 10999
rect 19073 10965 19107 10999
rect 19901 10965 19935 10999
rect 2053 10761 2087 10795
rect 3525 10761 3559 10795
rect 5181 10761 5215 10795
rect 6929 10761 6963 10795
rect 8677 10761 8711 10795
rect 9413 10761 9447 10795
rect 10517 10761 10551 10795
rect 12449 10761 12483 10795
rect 18613 10761 18647 10795
rect 20453 10761 20487 10795
rect 21465 10761 21499 10795
rect 9321 10693 9355 10727
rect 16773 10693 16807 10727
rect 2697 10625 2731 10659
rect 4077 10625 4111 10659
rect 4813 10625 4847 10659
rect 4997 10625 5031 10659
rect 5733 10625 5767 10659
rect 9873 10625 9907 10659
rect 10057 10625 10091 10659
rect 10885 10625 10919 10659
rect 13001 10625 13035 10659
rect 14105 10625 14139 10659
rect 15393 10625 15427 10659
rect 15577 10625 15611 10659
rect 16405 10625 16439 10659
rect 17877 10625 17911 10659
rect 19073 10625 19107 10659
rect 19257 10625 19291 10659
rect 20177 10625 20211 10659
rect 21005 10625 21039 10659
rect 1961 10557 1995 10591
rect 2513 10557 2547 10591
rect 7297 10557 7331 10591
rect 7564 10557 7598 10591
rect 11152 10557 11186 10591
rect 13921 10557 13955 10591
rect 16129 10557 16163 10591
rect 18061 10557 18095 10591
rect 18981 10557 19015 10591
rect 19993 10557 20027 10591
rect 21281 10557 21315 10591
rect 3893 10489 3927 10523
rect 12817 10489 12851 10523
rect 13277 10489 13311 10523
rect 16221 10489 16255 10523
rect 1777 10421 1811 10455
rect 2421 10421 2455 10455
rect 2881 10421 2915 10455
rect 3985 10421 4019 10455
rect 4353 10421 4387 10455
rect 4721 10421 4755 10455
rect 5549 10421 5583 10455
rect 5641 10421 5675 10455
rect 6009 10421 6043 10455
rect 9781 10421 9815 10455
rect 10241 10421 10275 10455
rect 12265 10421 12299 10455
rect 12909 10421 12943 10455
rect 13553 10421 13587 10455
rect 14013 10421 14047 10455
rect 14473 10421 14507 10455
rect 14933 10421 14967 10455
rect 15301 10421 15335 10455
rect 15761 10421 15795 10455
rect 19625 10421 19659 10455
rect 20085 10421 20119 10455
rect 20821 10421 20855 10455
rect 20913 10421 20947 10455
rect 2053 10217 2087 10251
rect 2421 10217 2455 10251
rect 3065 10217 3099 10251
rect 4537 10217 4571 10251
rect 4997 10217 5031 10251
rect 5365 10217 5399 10251
rect 6929 10217 6963 10251
rect 9229 10217 9263 10251
rect 10241 10217 10275 10251
rect 10517 10217 10551 10251
rect 13001 10217 13035 10251
rect 13369 10217 13403 10251
rect 14381 10217 14415 10251
rect 14749 10217 14783 10251
rect 16681 10217 16715 10251
rect 18153 10217 18187 10251
rect 18981 10217 19015 10251
rect 19349 10217 19383 10251
rect 3617 10149 3651 10183
rect 4169 10149 4203 10183
rect 4261 10149 4295 10183
rect 1685 10081 1719 10115
rect 2881 10081 2915 10115
rect 4905 10081 4939 10115
rect 1593 10013 1627 10047
rect 2513 10013 2547 10047
rect 2605 10013 2639 10047
rect 5089 10013 5123 10047
rect 15568 10149 15602 10183
rect 17018 10149 17052 10183
rect 18889 10149 18923 10183
rect 20545 10149 20579 10183
rect 5816 10081 5850 10115
rect 7389 10081 7423 10115
rect 8105 10081 8139 10115
rect 10425 10081 10459 10115
rect 10885 10081 10919 10115
rect 12909 10081 12943 10115
rect 15301 10081 15335 10115
rect 16773 10081 16807 10115
rect 19717 10081 19751 10115
rect 20269 10081 20303 10115
rect 5549 10013 5583 10047
rect 7481 10013 7515 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 10977 10013 11011 10047
rect 11161 10013 11195 10047
rect 13185 10013 13219 10047
rect 14841 10013 14875 10047
rect 15025 10013 15059 10047
rect 19073 10013 19107 10047
rect 19809 10013 19843 10047
rect 19993 10013 20027 10047
rect 12541 9945 12575 9979
rect 21281 9945 21315 9979
rect 1869 9877 1903 9911
rect 3801 9877 3835 9911
rect 5365 9877 5399 9911
rect 7021 9877 7055 9911
rect 18521 9877 18555 9911
rect 21557 9877 21591 9911
rect 6561 9673 6595 9707
rect 15485 9673 15519 9707
rect 20085 9673 20119 9707
rect 2053 9605 2087 9639
rect 4261 9605 4295 9639
rect 4629 9605 4663 9639
rect 7389 9605 7423 9639
rect 16313 9605 16347 9639
rect 19441 9605 19475 9639
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 5181 9537 5215 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 15945 9537 15979 9571
rect 16129 9537 16163 9571
rect 16865 9537 16899 9571
rect 19901 9537 19935 9571
rect 20637 9537 20671 9571
rect 21189 9537 21223 9571
rect 1501 9469 1535 9503
rect 8677 9469 8711 9503
rect 9873 9469 9907 9503
rect 9965 9469 9999 9503
rect 10232 9469 10266 9503
rect 12449 9469 12483 9503
rect 13921 9469 13955 9503
rect 14188 9469 14222 9503
rect 16773 9469 16807 9503
rect 18061 9469 18095 9503
rect 20913 9469 20947 9503
rect 1777 9401 1811 9435
rect 3148 9401 3182 9435
rect 4997 9401 5031 9435
rect 6929 9401 6963 9435
rect 7757 9401 7791 9435
rect 8217 9401 8251 9435
rect 12694 9401 12728 9435
rect 16681 9401 16715 9435
rect 18328 9401 18362 9435
rect 20453 9401 20487 9435
rect 2421 9333 2455 9367
rect 2513 9333 2547 9367
rect 4445 9333 4479 9367
rect 5089 9333 5123 9367
rect 8493 9333 8527 9367
rect 9873 9333 9907 9367
rect 11345 9333 11379 9367
rect 13829 9333 13863 9367
rect 15301 9333 15335 9367
rect 15853 9333 15887 9367
rect 17141 9333 17175 9367
rect 17325 9333 17359 9367
rect 20545 9333 20579 9367
rect 21557 9333 21591 9367
rect 3157 9129 3191 9163
rect 7113 9129 7147 9163
rect 7205 9129 7239 9163
rect 7665 9129 7699 9163
rect 8493 9129 8527 9163
rect 9045 9129 9079 9163
rect 9505 9129 9539 9163
rect 10241 9129 10275 9163
rect 10977 9129 11011 9163
rect 11069 9129 11103 9163
rect 13369 9129 13403 9163
rect 13737 9129 13771 9163
rect 14197 9129 14231 9163
rect 15301 9129 15335 9163
rect 15761 9129 15795 9163
rect 16129 9129 16163 9163
rect 18521 9129 18555 9163
rect 19993 9129 20027 9163
rect 21005 9129 21039 9163
rect 3525 9061 3559 9095
rect 12164 9061 12198 9095
rect 18880 9061 18914 9095
rect 1777 8993 1811 9027
rect 2044 8993 2078 9027
rect 3249 8993 3283 9027
rect 6193 8993 6227 9027
rect 8401 8993 8435 9027
rect 9321 8993 9355 9027
rect 10149 8993 10183 9027
rect 11437 8993 11471 9027
rect 11897 8993 11931 9027
rect 15669 8993 15703 9027
rect 16497 8993 16531 9027
rect 17408 8993 17442 9027
rect 6285 8925 6319 8959
rect 6377 8925 6411 8959
rect 7389 8925 7423 8959
rect 8585 8925 8619 8959
rect 8953 8925 8987 8959
rect 10425 8925 10459 8959
rect 11161 8925 11195 8959
rect 13829 8925 13863 8959
rect 13921 8925 13955 8959
rect 15853 8925 15887 8959
rect 17141 8925 17175 8959
rect 18613 8925 18647 8959
rect 20545 8925 20579 8959
rect 16681 8857 16715 8891
rect 21097 8857 21131 8891
rect 4261 8789 4295 8823
rect 5825 8789 5859 8823
rect 6745 8789 6779 8823
rect 8033 8789 8067 8823
rect 9781 8789 9815 8823
rect 10609 8789 10643 8823
rect 11713 8789 11747 8823
rect 13277 8789 13311 8823
rect 15025 8789 15059 8823
rect 21281 8789 21315 8823
rect 1961 8585 1995 8619
rect 2789 8585 2823 8619
rect 9873 8585 9907 8619
rect 13277 8585 13311 8619
rect 18889 8585 18923 8619
rect 19993 8585 20027 8619
rect 20821 8585 20855 8619
rect 4445 8517 4479 8551
rect 6837 8517 6871 8551
rect 7665 8517 7699 8551
rect 16681 8517 16715 8551
rect 2605 8449 2639 8483
rect 3433 8449 3467 8483
rect 4169 8449 4203 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 16313 8449 16347 8483
rect 17141 8449 17175 8483
rect 17325 8449 17359 8483
rect 18613 8449 18647 8483
rect 19349 8449 19383 8483
rect 19441 8449 19475 8483
rect 20545 8449 20579 8483
rect 21373 8449 21407 8483
rect 2329 8381 2363 8415
rect 5273 8381 5307 8415
rect 8401 8381 8435 8415
rect 8657 8381 8691 8415
rect 10241 8381 10275 8415
rect 16589 8381 16623 8415
rect 17049 8381 17083 8415
rect 18521 8381 18555 8415
rect 19717 8381 19751 8415
rect 20453 8381 20487 8415
rect 21189 8381 21223 8415
rect 2421 8313 2455 8347
rect 3157 8313 3191 8347
rect 4077 8313 4111 8347
rect 4813 8313 4847 8347
rect 5540 8313 5574 8347
rect 7205 8313 7239 8347
rect 19257 8313 19291 8347
rect 21281 8313 21315 8347
rect 3249 8245 3283 8279
rect 3617 8245 3651 8279
rect 3985 8245 4019 8279
rect 6653 8245 6687 8279
rect 9781 8245 9815 8279
rect 18061 8245 18095 8279
rect 18429 8245 18463 8279
rect 20361 8245 20395 8279
rect 3433 8041 3467 8075
rect 4537 8041 4571 8075
rect 6101 8041 6135 8075
rect 9505 8041 9539 8075
rect 18337 8041 18371 8075
rect 2320 7905 2354 7939
rect 4988 7905 5022 7939
rect 6817 7905 6851 7939
rect 8300 7905 8334 7939
rect 2053 7837 2087 7871
rect 3525 7837 3559 7871
rect 4721 7837 4755 7871
rect 6561 7837 6595 7871
rect 8033 7837 8067 7871
rect 17224 7973 17258 8007
rect 21189 7973 21223 8007
rect 19616 7905 19650 7939
rect 20913 7905 20947 7939
rect 16957 7837 16991 7871
rect 19349 7837 19383 7871
rect 7941 7769 7975 7803
rect 9505 7769 9539 7803
rect 3801 7701 3835 7735
rect 9413 7701 9447 7735
rect 19073 7701 19107 7735
rect 20729 7701 20763 7735
rect 2881 7497 2915 7531
rect 3709 7497 3743 7531
rect 5733 7497 5767 7531
rect 7297 7497 7331 7531
rect 8217 7497 8251 7531
rect 20637 7497 20671 7531
rect 20545 7429 20579 7463
rect 2605 7361 2639 7395
rect 3341 7361 3375 7395
rect 3525 7361 3559 7395
rect 4353 7361 4387 7395
rect 5365 7361 5399 7395
rect 5549 7361 5583 7395
rect 6377 7361 6411 7395
rect 7757 7361 7791 7395
rect 7941 7361 7975 7395
rect 19165 7361 19199 7395
rect 21189 7361 21223 7395
rect 4077 7293 4111 7327
rect 19432 7293 19466 7327
rect 6193 7225 6227 7259
rect 7665 7225 7699 7259
rect 21097 7225 21131 7259
rect 2697 7157 2731 7191
rect 3249 7157 3283 7191
rect 4169 7157 4203 7191
rect 4629 7157 4663 7191
rect 4905 7157 4939 7191
rect 5273 7157 5307 7191
rect 6101 7157 6135 7191
rect 21005 7157 21039 7191
rect 5181 6953 5215 6987
rect 4353 6885 4387 6919
rect 1961 6817 1995 6851
rect 2228 6817 2262 6851
rect 3433 6817 3467 6851
rect 20453 6817 20487 6851
rect 5273 6749 5307 6783
rect 5457 6749 5491 6783
rect 3341 6681 3375 6715
rect 4445 6681 4479 6715
rect 4813 6681 4847 6715
rect 3617 6613 3651 6647
rect 4629 6613 4663 6647
rect 20269 6409 20303 6443
rect 20821 6273 20855 6307
rect 20637 6137 20671 6171
rect 20085 6069 20119 6103
rect 20729 6069 20763 6103
rect 21097 6069 21131 6103
rect 5457 3009 5491 3043
rect 15669 3009 15703 3043
rect 4813 2941 4847 2975
rect 5089 2941 5123 2975
rect 5549 2941 5583 2975
rect 5825 2941 5859 2975
rect 15485 2941 15519 2975
rect 16037 2941 16071 2975
rect 6193 2805 6227 2839
<< metal1 >>
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 6362 21128 6368 21140
rect 4120 21100 6368 21128
rect 4120 21088 4126 21100
rect 6362 21088 6368 21100
rect 6420 21088 6426 21140
rect 2314 20884 2320 20936
rect 2372 20924 2378 20936
rect 3050 20924 3056 20936
rect 2372 20896 3056 20924
rect 2372 20884 2378 20896
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 17681 20587 17739 20593
rect 17681 20553 17693 20587
rect 17727 20584 17739 20587
rect 18598 20584 18604 20596
rect 17727 20556 18604 20584
rect 17727 20553 17739 20556
rect 17681 20547 17739 20553
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19702 20584 19708 20596
rect 19475 20556 19708 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19702 20544 19708 20556
rect 19760 20544 19766 20596
rect 8757 20519 8815 20525
rect 8757 20485 8769 20519
rect 8803 20516 8815 20519
rect 9674 20516 9680 20528
rect 8803 20488 9680 20516
rect 8803 20485 8815 20488
rect 8757 20479 8815 20485
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 17313 20519 17371 20525
rect 17313 20485 17325 20519
rect 17359 20516 17371 20519
rect 18046 20516 18052 20528
rect 17359 20488 18052 20516
rect 17359 20485 17371 20488
rect 17313 20479 17371 20485
rect 18046 20476 18052 20488
rect 18104 20476 18110 20528
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20448 9459 20451
rect 10042 20448 10048 20460
rect 9447 20420 10048 20448
rect 9447 20417 9459 20420
rect 9401 20411 9459 20417
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20380 2191 20383
rect 2222 20380 2228 20392
rect 2179 20352 2228 20380
rect 2179 20349 2191 20352
rect 2133 20343 2191 20349
rect 2222 20340 2228 20352
rect 2280 20340 2286 20392
rect 14090 20340 14096 20392
rect 14148 20380 14154 20392
rect 14642 20380 14648 20392
rect 14148 20352 14648 20380
rect 14148 20340 14154 20352
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 17126 20380 17132 20392
rect 17087 20352 17132 20380
rect 17126 20340 17132 20352
rect 17184 20340 17190 20392
rect 17494 20380 17500 20392
rect 17455 20352 17500 20380
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 19058 20340 19064 20392
rect 19116 20380 19122 20392
rect 19153 20383 19211 20389
rect 19153 20380 19165 20383
rect 19116 20352 19165 20380
rect 19116 20340 19122 20352
rect 19153 20349 19165 20352
rect 19199 20380 19211 20383
rect 19245 20383 19303 20389
rect 19245 20380 19257 20383
rect 19199 20352 19257 20380
rect 19199 20349 19211 20352
rect 19153 20343 19211 20349
rect 19245 20349 19257 20352
rect 19291 20349 19303 20383
rect 19245 20343 19303 20349
rect 8846 20272 8852 20324
rect 8904 20312 8910 20324
rect 9125 20315 9183 20321
rect 9125 20312 9137 20315
rect 8904 20284 9137 20312
rect 8904 20272 8910 20284
rect 9125 20281 9137 20284
rect 9171 20281 9183 20315
rect 9125 20275 9183 20281
rect 14550 20272 14556 20324
rect 14608 20312 14614 20324
rect 15102 20312 15108 20324
rect 14608 20284 15108 20312
rect 14608 20272 14614 20284
rect 15102 20272 15108 20284
rect 15160 20272 15166 20324
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 2130 20204 2136 20256
rect 2188 20244 2194 20256
rect 2317 20247 2375 20253
rect 2317 20244 2329 20247
rect 2188 20216 2329 20244
rect 2188 20204 2194 20216
rect 2317 20213 2329 20216
rect 2363 20244 2375 20247
rect 7282 20244 7288 20256
rect 2363 20216 7288 20244
rect 2363 20213 2375 20216
rect 2317 20207 2375 20213
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 9214 20244 9220 20256
rect 9175 20216 9220 20244
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 17218 20244 17224 20256
rect 13136 20216 17224 20244
rect 13136 20204 13142 20216
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 20346 20244 20352 20256
rect 20307 20216 20352 20244
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 20809 20247 20867 20253
rect 20809 20213 20821 20247
rect 20855 20244 20867 20247
rect 21174 20244 21180 20256
rect 20855 20216 21180 20244
rect 20855 20213 20867 20216
rect 20809 20207 20867 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 2041 20043 2099 20049
rect 2041 20009 2053 20043
rect 2087 20040 2099 20043
rect 2774 20040 2780 20052
rect 2087 20012 2780 20040
rect 2087 20009 2099 20012
rect 2041 20003 2099 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 8757 20043 8815 20049
rect 8757 20009 8769 20043
rect 8803 20040 8815 20043
rect 9214 20040 9220 20052
rect 8803 20012 9220 20040
rect 8803 20009 8815 20012
rect 8757 20003 8815 20009
rect 9214 20000 9220 20012
rect 9272 20000 9278 20052
rect 11517 20043 11575 20049
rect 11517 20009 11529 20043
rect 11563 20009 11575 20043
rect 13078 20040 13084 20052
rect 13039 20012 13084 20040
rect 11517 20003 11575 20009
rect 3237 19975 3295 19981
rect 2516 19944 3096 19972
rect 1486 19904 1492 19916
rect 1447 19876 1492 19904
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19904 1915 19907
rect 2130 19904 2136 19916
rect 1903 19876 2136 19904
rect 1903 19873 1915 19876
rect 1857 19867 1915 19873
rect 2130 19864 2136 19876
rect 2188 19864 2194 19916
rect 2222 19864 2228 19916
rect 2280 19904 2286 19916
rect 2516 19904 2544 19944
rect 2581 19907 2639 19913
rect 2581 19904 2593 19907
rect 2280 19876 2325 19904
rect 2516 19876 2593 19904
rect 2280 19864 2286 19876
rect 2581 19873 2593 19876
rect 2627 19873 2639 19907
rect 2581 19867 2639 19873
rect 3068 19845 3096 19944
rect 3237 19941 3249 19975
rect 3283 19972 3295 19975
rect 3418 19972 3424 19984
rect 3283 19944 3424 19972
rect 3283 19941 3295 19944
rect 3237 19935 3295 19941
rect 3418 19932 3424 19944
rect 3476 19972 3482 19984
rect 3476 19944 9812 19972
rect 3476 19932 3482 19944
rect 8478 19864 8484 19916
rect 8536 19904 8542 19916
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 8536 19876 9137 19904
rect 8536 19864 8542 19876
rect 9125 19873 9137 19876
rect 9171 19904 9183 19907
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9171 19876 9689 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9784 19904 9812 19944
rect 10042 19932 10048 19984
rect 10100 19981 10106 19984
rect 10100 19975 10164 19981
rect 10100 19941 10118 19975
rect 10152 19941 10164 19975
rect 10100 19935 10164 19941
rect 10100 19932 10106 19935
rect 10594 19904 10600 19916
rect 9784 19876 10600 19904
rect 9677 19867 9735 19873
rect 10594 19864 10600 19876
rect 10652 19864 10658 19916
rect 11532 19904 11560 20003
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13449 20043 13507 20049
rect 13449 20009 13461 20043
rect 13495 20040 13507 20043
rect 14001 20043 14059 20049
rect 14001 20040 14013 20043
rect 13495 20012 14013 20040
rect 13495 20009 13507 20012
rect 13449 20003 13507 20009
rect 14001 20009 14013 20012
rect 14047 20040 14059 20043
rect 14366 20040 14372 20052
rect 14047 20012 14372 20040
rect 14047 20009 14059 20012
rect 14001 20003 14059 20009
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 14550 20040 14556 20052
rect 14511 20012 14556 20040
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 15470 20040 15476 20052
rect 15431 20012 15476 20040
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 15930 20000 15936 20052
rect 15988 20040 15994 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 15988 20012 16865 20040
rect 15988 20000 15994 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 17221 20043 17279 20049
rect 17221 20009 17233 20043
rect 17267 20040 17279 20043
rect 17586 20040 17592 20052
rect 17267 20012 17592 20040
rect 17267 20009 17279 20012
rect 17221 20003 17279 20009
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 18417 20043 18475 20049
rect 18417 20009 18429 20043
rect 18463 20040 18475 20043
rect 18874 20040 18880 20052
rect 18463 20012 18880 20040
rect 18463 20009 18475 20012
rect 18417 20003 18475 20009
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 21453 20043 21511 20049
rect 21453 20040 21465 20043
rect 20680 20012 21465 20040
rect 20680 20000 20686 20012
rect 21453 20009 21465 20012
rect 21499 20009 21511 20043
rect 21453 20003 21511 20009
rect 11885 19975 11943 19981
rect 11885 19941 11897 19975
rect 11931 19972 11943 19975
rect 12526 19972 12532 19984
rect 11931 19944 12532 19972
rect 11931 19941 11943 19944
rect 11885 19935 11943 19941
rect 12526 19932 12532 19944
rect 12584 19932 12590 19984
rect 13909 19975 13967 19981
rect 13909 19941 13921 19975
rect 13955 19972 13967 19975
rect 14737 19975 14795 19981
rect 14737 19972 14749 19975
rect 13955 19944 14749 19972
rect 13955 19941 13967 19944
rect 13909 19935 13967 19941
rect 14737 19941 14749 19944
rect 14783 19941 14795 19975
rect 14737 19935 14795 19941
rect 16393 19975 16451 19981
rect 16393 19941 16405 19975
rect 16439 19972 16451 19975
rect 17494 19972 17500 19984
rect 16439 19944 17500 19972
rect 16439 19941 16451 19944
rect 16393 19935 16451 19941
rect 17494 19932 17500 19944
rect 17552 19932 17558 19984
rect 20073 19975 20131 19981
rect 20073 19972 20085 19975
rect 18616 19944 20085 19972
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 11532 19876 12357 19904
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 12345 19867 12403 19873
rect 12621 19907 12679 19913
rect 12621 19873 12633 19907
rect 12667 19904 12679 19907
rect 12897 19907 12955 19913
rect 12897 19904 12909 19907
rect 12667 19876 12909 19904
rect 12667 19873 12679 19876
rect 12621 19867 12679 19873
rect 12897 19873 12909 19876
rect 12943 19873 12955 19907
rect 14369 19907 14427 19913
rect 12897 19867 12955 19873
rect 13832 19876 14136 19904
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19836 3111 19839
rect 3234 19836 3240 19848
rect 3099 19808 3240 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9398 19836 9404 19848
rect 9359 19808 9404 19836
rect 9217 19799 9275 19805
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 2406 19700 2412 19712
rect 2367 19672 2412 19700
rect 2406 19660 2412 19672
rect 2464 19660 2470 19712
rect 2777 19703 2835 19709
rect 2777 19669 2789 19703
rect 2823 19700 2835 19703
rect 4062 19700 4068 19712
rect 2823 19672 4068 19700
rect 2823 19669 2835 19672
rect 2777 19663 2835 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 8573 19703 8631 19709
rect 8573 19700 8585 19703
rect 8352 19672 8585 19700
rect 8352 19660 8358 19672
rect 8573 19669 8585 19672
rect 8619 19700 8631 19703
rect 9232 19700 9260 19799
rect 9398 19796 9404 19808
rect 9456 19796 9462 19848
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 9861 19839 9919 19845
rect 9861 19836 9873 19839
rect 9824 19808 9873 19836
rect 9824 19796 9830 19808
rect 9861 19805 9873 19808
rect 9907 19805 9919 19839
rect 11974 19836 11980 19848
rect 11935 19808 11980 19836
rect 9861 19799 9919 19805
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 13832 19836 13860 19876
rect 14108 19845 14136 19876
rect 14369 19873 14381 19907
rect 14415 19873 14427 19907
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 14369 19867 14427 19873
rect 12124 19808 12169 19836
rect 12636 19808 13860 19836
rect 14093 19839 14151 19845
rect 12124 19796 12130 19808
rect 11698 19728 11704 19780
rect 11756 19768 11762 19780
rect 12158 19768 12164 19780
rect 11756 19740 12164 19768
rect 11756 19728 11762 19740
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 12636 19712 12664 19808
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 13538 19768 13544 19780
rect 13499 19740 13544 19768
rect 13538 19728 13544 19740
rect 13596 19728 13602 19780
rect 9306 19700 9312 19712
rect 8619 19672 9312 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 11241 19703 11299 19709
rect 11241 19669 11253 19703
rect 11287 19700 11299 19703
rect 12618 19700 12624 19712
rect 11287 19672 12624 19700
rect 11287 19669 11299 19672
rect 11241 19663 11299 19669
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 13170 19660 13176 19712
rect 13228 19700 13234 19712
rect 14384 19700 14412 19867
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 16114 19904 16120 19916
rect 16075 19876 16120 19904
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 18616 19913 18644 19944
rect 20073 19941 20085 19944
rect 20119 19941 20131 19975
rect 20073 19935 20131 19941
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 16632 19876 16681 19904
rect 16632 19864 16638 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 17037 19907 17095 19913
rect 17037 19873 17049 19907
rect 17083 19873 17095 19907
rect 17037 19867 17095 19873
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19873 17647 19907
rect 17589 19867 17647 19873
rect 17865 19907 17923 19913
rect 17865 19873 17877 19907
rect 17911 19904 17923 19907
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 17911 19876 18245 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 18233 19867 18291 19873
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19873 18659 19907
rect 19334 19904 19340 19916
rect 19295 19876 19340 19904
rect 18601 19867 18659 19873
rect 15562 19796 15568 19848
rect 15620 19836 15626 19848
rect 17052 19836 17080 19867
rect 15620 19808 17080 19836
rect 17604 19836 17632 19867
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19797 19907 19855 19913
rect 19797 19904 19809 19907
rect 19484 19876 19529 19904
rect 19628 19876 19809 19904
rect 19484 19864 19490 19876
rect 18046 19836 18052 19848
rect 17604 19808 18052 19836
rect 15620 19796 15626 19808
rect 18046 19796 18052 19808
rect 18104 19796 18110 19848
rect 19242 19836 19248 19848
rect 18800 19808 19248 19836
rect 14550 19728 14556 19780
rect 14608 19768 14614 19780
rect 18800 19777 18828 19808
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 19518 19836 19524 19848
rect 19479 19808 19524 19836
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 18785 19771 18843 19777
rect 14608 19740 18736 19768
rect 14608 19728 14614 19740
rect 13228 19672 14412 19700
rect 13228 19660 13234 19672
rect 14458 19660 14464 19712
rect 14516 19700 14522 19712
rect 15013 19703 15071 19709
rect 15013 19700 15025 19703
rect 14516 19672 15025 19700
rect 14516 19660 14522 19672
rect 15013 19669 15025 19672
rect 15059 19669 15071 19703
rect 18708 19700 18736 19740
rect 18785 19737 18797 19771
rect 18831 19737 18843 19771
rect 18785 19731 18843 19737
rect 18969 19771 19027 19777
rect 18969 19737 18981 19771
rect 19015 19768 19027 19771
rect 19628 19768 19656 19876
rect 19797 19873 19809 19876
rect 19843 19873 19855 19907
rect 19797 19867 19855 19873
rect 20441 19907 20499 19913
rect 20441 19873 20453 19907
rect 20487 19904 20499 19907
rect 20806 19904 20812 19916
rect 20487 19876 20812 19904
rect 20487 19873 20499 19876
rect 20441 19867 20499 19873
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19904 20959 19907
rect 21174 19904 21180 19916
rect 20947 19876 21180 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 20916 19836 20944 19867
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19904 21327 19907
rect 21450 19904 21456 19916
rect 21315 19876 21456 19904
rect 21315 19873 21327 19876
rect 21269 19867 21327 19873
rect 21450 19864 21456 19876
rect 21508 19864 21514 19916
rect 19015 19740 19656 19768
rect 20456 19808 20944 19836
rect 19015 19737 19027 19740
rect 18969 19731 19027 19737
rect 20456 19700 20484 19808
rect 20530 19728 20536 19780
rect 20588 19768 20594 19780
rect 21085 19771 21143 19777
rect 21085 19768 21097 19771
rect 20588 19740 21097 19768
rect 20588 19728 20594 19740
rect 21085 19737 21097 19740
rect 21131 19737 21143 19771
rect 21085 19731 21143 19737
rect 18708 19672 20484 19700
rect 20625 19703 20683 19709
rect 15013 19663 15071 19669
rect 20625 19669 20637 19703
rect 20671 19700 20683 19703
rect 22278 19700 22284 19712
rect 20671 19672 22284 19700
rect 20671 19669 20683 19672
rect 20625 19663 20683 19669
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 3142 19496 3148 19508
rect 3103 19468 3148 19496
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 3602 19496 3608 19508
rect 3563 19468 3608 19496
rect 3602 19456 3608 19468
rect 3660 19456 3666 19508
rect 6362 19496 6368 19508
rect 6323 19468 6368 19496
rect 6362 19456 6368 19468
rect 6420 19456 6426 19508
rect 9033 19499 9091 19505
rect 9033 19465 9045 19499
rect 9079 19496 9091 19499
rect 9398 19496 9404 19508
rect 9079 19468 9404 19496
rect 9079 19465 9091 19468
rect 9033 19459 9091 19465
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10505 19499 10563 19505
rect 10505 19496 10517 19499
rect 10100 19468 10517 19496
rect 10100 19456 10106 19468
rect 10505 19465 10517 19468
rect 10551 19465 10563 19499
rect 10505 19459 10563 19465
rect 10594 19456 10600 19508
rect 10652 19496 10658 19508
rect 14366 19496 14372 19508
rect 10652 19468 14372 19496
rect 10652 19456 10658 19468
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 15657 19499 15715 19505
rect 15657 19465 15669 19499
rect 15703 19496 15715 19499
rect 16114 19496 16120 19508
rect 15703 19468 16120 19496
rect 15703 19465 15715 19468
rect 15657 19459 15715 19465
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 18046 19496 18052 19508
rect 18007 19468 18052 19496
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 20625 19499 20683 19505
rect 20625 19465 20637 19499
rect 20671 19496 20683 19499
rect 20714 19496 20720 19508
rect 20671 19468 20720 19496
rect 20671 19465 20683 19468
rect 20625 19459 20683 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 20990 19496 20996 19508
rect 20951 19468 20996 19496
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21358 19496 21364 19508
rect 21319 19468 21364 19496
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 2590 19388 2596 19440
rect 2648 19428 2654 19440
rect 14001 19431 14059 19437
rect 2648 19400 2728 19428
rect 2648 19388 2654 19400
rect 1489 19295 1547 19301
rect 1489 19261 1501 19295
rect 1535 19292 1547 19295
rect 1578 19292 1584 19304
rect 1535 19264 1584 19292
rect 1535 19261 1547 19264
rect 1489 19255 1547 19261
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 2225 19295 2283 19301
rect 2225 19261 2237 19295
rect 2271 19292 2283 19295
rect 2314 19292 2320 19304
rect 2271 19264 2320 19292
rect 2271 19261 2283 19264
rect 2225 19255 2283 19261
rect 198 19184 204 19236
rect 256 19224 262 19236
rect 1302 19224 1308 19236
rect 256 19196 1308 19224
rect 256 19184 262 19196
rect 1302 19184 1308 19196
rect 1360 19224 1366 19236
rect 1872 19224 1900 19255
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 2700 19292 2728 19400
rect 14001 19397 14013 19431
rect 14047 19428 14059 19431
rect 14918 19428 14924 19440
rect 14047 19400 14924 19428
rect 14047 19397 14059 19400
rect 14001 19391 14059 19397
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 13556 19332 14565 19360
rect 2639 19264 2728 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 2774 19252 2780 19304
rect 2832 19252 2838 19304
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 3142 19292 3148 19304
rect 3007 19264 3148 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 3421 19295 3479 19301
rect 3421 19261 3433 19295
rect 3467 19292 3479 19295
rect 3510 19292 3516 19304
rect 3467 19264 3516 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 3510 19252 3516 19264
rect 3568 19252 3574 19304
rect 3970 19292 3976 19304
rect 3931 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19292 4034 19304
rect 4985 19295 5043 19301
rect 4985 19292 4997 19295
rect 4028 19264 4997 19292
rect 4028 19252 4034 19264
rect 4985 19261 4997 19264
rect 5031 19261 5043 19295
rect 4985 19255 5043 19261
rect 6181 19295 6239 19301
rect 6181 19261 6193 19295
rect 6227 19292 6239 19295
rect 6822 19292 6828 19304
rect 6227 19264 6828 19292
rect 6227 19261 6239 19264
rect 6181 19255 6239 19261
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 7006 19252 7012 19304
rect 7064 19292 7070 19304
rect 9398 19301 9404 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 7064 19264 7665 19292
rect 7064 19252 7070 19264
rect 7653 19261 7665 19264
rect 7699 19292 7711 19295
rect 9125 19295 9183 19301
rect 9125 19292 9137 19295
rect 7699 19264 9137 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 9125 19261 9137 19264
rect 9171 19261 9183 19295
rect 9392 19292 9404 19301
rect 9359 19264 9404 19292
rect 9125 19255 9183 19261
rect 9392 19255 9404 19264
rect 9398 19252 9404 19255
rect 9456 19252 9462 19304
rect 10870 19292 10876 19304
rect 10831 19264 10876 19292
rect 10870 19252 10876 19264
rect 10928 19292 10934 19304
rect 12529 19295 12587 19301
rect 12529 19292 12541 19295
rect 10928 19264 12541 19292
rect 10928 19252 10934 19264
rect 12529 19261 12541 19264
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 12785 19295 12843 19301
rect 12785 19292 12797 19295
rect 12676 19264 12797 19292
rect 12676 19252 12682 19264
rect 12785 19261 12797 19264
rect 12831 19292 12843 19295
rect 13556 19292 13584 19332
rect 14553 19329 14565 19332
rect 14599 19329 14611 19363
rect 15381 19363 15439 19369
rect 15381 19360 15393 19363
rect 14553 19323 14611 19329
rect 14752 19332 15393 19360
rect 14752 19292 14780 19332
rect 15381 19329 15393 19332
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 16022 19320 16028 19372
rect 16080 19360 16086 19372
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 16080 19332 16221 19360
rect 16080 19320 16086 19332
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 16761 19363 16819 19369
rect 16761 19329 16773 19363
rect 16807 19360 16819 19363
rect 17126 19360 17132 19372
rect 16807 19332 17132 19360
rect 16807 19329 16819 19332
rect 16761 19323 16819 19329
rect 17126 19320 17132 19332
rect 17184 19320 17190 19372
rect 18598 19360 18604 19372
rect 18559 19332 18604 19360
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 16485 19295 16543 19301
rect 16485 19292 16497 19295
rect 12831 19264 13584 19292
rect 13924 19264 14780 19292
rect 14844 19264 16497 19292
rect 12831 19261 12843 19264
rect 12785 19255 12843 19261
rect 2792 19224 2820 19252
rect 1360 19196 1900 19224
rect 2424 19196 2820 19224
rect 1360 19184 1366 19196
rect 1673 19159 1731 19165
rect 1673 19125 1685 19159
rect 1719 19156 1731 19159
rect 1854 19156 1860 19168
rect 1719 19128 1860 19156
rect 1719 19125 1731 19128
rect 1673 19119 1731 19125
rect 1854 19116 1860 19128
rect 1912 19116 1918 19168
rect 2038 19156 2044 19168
rect 1999 19128 2044 19156
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 2424 19165 2452 19196
rect 3050 19184 3056 19236
rect 3108 19224 3114 19236
rect 4338 19224 4344 19236
rect 3108 19196 4344 19224
rect 3108 19184 3114 19196
rect 4338 19184 4344 19196
rect 4396 19184 4402 19236
rect 4709 19227 4767 19233
rect 4709 19193 4721 19227
rect 4755 19224 4767 19227
rect 7558 19224 7564 19236
rect 4755 19196 7564 19224
rect 4755 19193 4767 19196
rect 4709 19187 4767 19193
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 7920 19227 7978 19233
rect 7920 19193 7932 19227
rect 7966 19224 7978 19227
rect 11140 19227 11198 19233
rect 7966 19196 10824 19224
rect 7966 19193 7978 19196
rect 7920 19187 7978 19193
rect 2409 19159 2467 19165
rect 2409 19125 2421 19159
rect 2455 19125 2467 19159
rect 2409 19119 2467 19125
rect 2777 19159 2835 19165
rect 2777 19125 2789 19159
rect 2823 19156 2835 19159
rect 2866 19156 2872 19168
rect 2823 19128 2872 19156
rect 2823 19125 2835 19128
rect 2777 19119 2835 19125
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 4356 19156 4384 19184
rect 8294 19156 8300 19168
rect 4356 19128 8300 19156
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 10594 19116 10600 19168
rect 10652 19156 10658 19168
rect 10796 19156 10824 19196
rect 11140 19193 11152 19227
rect 11186 19224 11198 19227
rect 12342 19224 12348 19236
rect 11186 19196 12348 19224
rect 11186 19193 11198 19196
rect 11140 19187 11198 19193
rect 12342 19184 12348 19196
rect 12400 19224 12406 19236
rect 13078 19224 13084 19236
rect 12400 19196 13084 19224
rect 12400 19184 12406 19196
rect 13078 19184 13084 19196
rect 13136 19184 13142 19236
rect 13924 19168 13952 19264
rect 12066 19156 12072 19168
rect 10652 19128 10697 19156
rect 10796 19128 12072 19156
rect 10652 19116 10658 19128
rect 12066 19116 12072 19128
rect 12124 19156 12130 19168
rect 12253 19159 12311 19165
rect 12253 19156 12265 19159
rect 12124 19128 12265 19156
rect 12124 19116 12130 19128
rect 12253 19125 12265 19128
rect 12299 19125 12311 19159
rect 13906 19156 13912 19168
rect 13819 19128 13912 19156
rect 12253 19119 12311 19125
rect 13906 19116 13912 19128
rect 13964 19116 13970 19168
rect 14366 19156 14372 19168
rect 14327 19128 14372 19156
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 14844 19165 14872 19264
rect 16485 19261 16497 19264
rect 16531 19261 16543 19295
rect 17034 19292 17040 19304
rect 16995 19264 17040 19292
rect 16485 19255 16543 19261
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 17402 19292 17408 19304
rect 17363 19264 17408 19292
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18969 19295 19027 19301
rect 18969 19292 18981 19295
rect 17920 19264 18981 19292
rect 17920 19252 17926 19264
rect 18969 19261 18981 19264
rect 19015 19261 19027 19295
rect 18969 19255 19027 19261
rect 19978 19252 19984 19304
rect 20036 19292 20042 19304
rect 20346 19292 20352 19304
rect 20036 19264 20352 19292
rect 20036 19252 20042 19264
rect 20346 19252 20352 19264
rect 20404 19292 20410 19304
rect 20441 19295 20499 19301
rect 20441 19292 20453 19295
rect 20404 19264 20453 19292
rect 20404 19252 20410 19264
rect 20441 19261 20453 19264
rect 20487 19261 20499 19295
rect 20441 19255 20499 19261
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20772 19264 20821 19292
rect 20772 19252 20778 19264
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 21177 19295 21235 19301
rect 21177 19261 21189 19295
rect 21223 19292 21235 19295
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21223 19264 22017 19292
rect 21223 19261 21235 19264
rect 21177 19255 21235 19261
rect 22005 19261 22017 19264
rect 22051 19261 22063 19295
rect 22005 19255 22063 19261
rect 14918 19184 14924 19236
rect 14976 19224 14982 19236
rect 15289 19227 15347 19233
rect 15289 19224 15301 19227
rect 14976 19196 15301 19224
rect 14976 19184 14982 19196
rect 15289 19193 15301 19196
rect 15335 19193 15347 19227
rect 15289 19187 15347 19193
rect 16758 19184 16764 19236
rect 16816 19224 16822 19236
rect 16816 19196 17632 19224
rect 16816 19184 16822 19196
rect 14829 19159 14887 19165
rect 14516 19128 14561 19156
rect 14516 19116 14522 19128
rect 14829 19125 14841 19159
rect 14875 19125 14887 19159
rect 15194 19156 15200 19168
rect 15155 19128 15200 19156
rect 14829 19119 14887 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15436 19128 16037 19156
rect 15436 19116 15442 19128
rect 16025 19125 16037 19128
rect 16071 19125 16083 19159
rect 16025 19119 16083 19125
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16172 19128 16217 19156
rect 16172 19116 16178 19128
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 17604 19165 17632 19196
rect 17954 19184 17960 19236
rect 18012 19224 18018 19236
rect 18509 19227 18567 19233
rect 18509 19224 18521 19227
rect 18012 19196 18521 19224
rect 18012 19184 18018 19196
rect 18509 19193 18521 19196
rect 18555 19193 18567 19227
rect 18509 19187 18567 19193
rect 19236 19227 19294 19233
rect 19236 19193 19248 19227
rect 19282 19224 19294 19227
rect 19702 19224 19708 19236
rect 19282 19196 19708 19224
rect 19282 19193 19294 19196
rect 19236 19187 19294 19193
rect 19702 19184 19708 19196
rect 19760 19184 19766 19236
rect 17221 19159 17279 19165
rect 17221 19156 17233 19159
rect 16356 19128 17233 19156
rect 16356 19116 16362 19128
rect 17221 19125 17233 19128
rect 17267 19125 17279 19159
rect 17221 19119 17279 19125
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19125 17647 19159
rect 17589 19119 17647 19125
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18417 19159 18475 19165
rect 18417 19156 18429 19159
rect 18104 19128 18429 19156
rect 18104 19116 18110 19128
rect 18417 19125 18429 19128
rect 18463 19125 18475 19159
rect 18417 19119 18475 19125
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 20349 19159 20407 19165
rect 20349 19156 20361 19159
rect 19576 19128 20361 19156
rect 19576 19116 19582 19128
rect 20349 19125 20361 19128
rect 20395 19125 20407 19159
rect 20349 19119 20407 19125
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1302 18912 1308 18964
rect 1360 18952 1366 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1360 18924 1593 18952
rect 1360 18912 1366 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 1762 18912 1768 18964
rect 1820 18912 1826 18964
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 2317 18955 2375 18961
rect 2317 18921 2329 18955
rect 2363 18952 2375 18955
rect 2958 18952 2964 18964
rect 2363 18924 2964 18952
rect 2363 18921 2375 18924
rect 2317 18915 2375 18921
rect 2958 18912 2964 18924
rect 3016 18912 3022 18964
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3421 18955 3479 18961
rect 3421 18952 3433 18955
rect 3200 18924 3433 18952
rect 3200 18912 3206 18924
rect 3421 18921 3433 18924
rect 3467 18952 3479 18955
rect 3786 18952 3792 18964
rect 3467 18924 3792 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 3786 18912 3792 18924
rect 3844 18952 3850 18964
rect 8294 18952 8300 18964
rect 3844 18924 6132 18952
rect 3844 18912 3850 18924
rect 1780 18884 1808 18912
rect 6104 18884 6132 18924
rect 6463 18924 8300 18952
rect 6463 18884 6491 18924
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 8757 18955 8815 18961
rect 8757 18921 8769 18955
rect 8803 18952 8815 18955
rect 8846 18952 8852 18964
rect 8803 18924 8852 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 8846 18912 8852 18924
rect 8904 18912 8910 18964
rect 9125 18955 9183 18961
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 10594 18952 10600 18964
rect 9171 18924 10600 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 10594 18912 10600 18924
rect 10652 18912 10658 18964
rect 11149 18955 11207 18961
rect 11149 18921 11161 18955
rect 11195 18952 11207 18955
rect 11330 18952 11336 18964
rect 11195 18924 11336 18952
rect 11195 18921 11207 18924
rect 11149 18915 11207 18921
rect 11330 18912 11336 18924
rect 11388 18912 11394 18964
rect 11701 18955 11759 18961
rect 11701 18921 11713 18955
rect 11747 18952 11759 18955
rect 11974 18952 11980 18964
rect 11747 18924 11980 18952
rect 11747 18921 11759 18924
rect 11701 18915 11759 18921
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 12066 18912 12072 18964
rect 12124 18952 12130 18964
rect 13357 18955 13415 18961
rect 13357 18952 13369 18955
rect 12124 18924 13369 18952
rect 12124 18912 12130 18924
rect 13357 18921 13369 18924
rect 13403 18921 13415 18955
rect 13357 18915 13415 18921
rect 15289 18955 15347 18961
rect 15289 18921 15301 18955
rect 15335 18952 15347 18955
rect 16114 18952 16120 18964
rect 15335 18924 16120 18952
rect 15335 18921 15347 18924
rect 15289 18915 15347 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 18233 18955 18291 18961
rect 18233 18921 18245 18955
rect 18279 18921 18291 18955
rect 18233 18915 18291 18921
rect 6822 18884 6828 18896
rect 1780 18856 5396 18884
rect 6104 18856 6491 18884
rect 6783 18856 6828 18884
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18785 2191 18819
rect 2133 18779 2191 18785
rect 2501 18819 2559 18825
rect 2501 18785 2513 18819
rect 2547 18816 2559 18819
rect 2547 18788 3004 18816
rect 2547 18785 2559 18788
rect 2501 18779 2559 18785
rect 2148 18680 2176 18779
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 2976 18757 3004 18788
rect 2961 18751 3019 18757
rect 2372 18720 2912 18748
rect 2372 18708 2378 18720
rect 2498 18680 2504 18692
rect 2148 18652 2504 18680
rect 2498 18640 2504 18652
rect 2556 18640 2562 18692
rect 2682 18680 2688 18692
rect 2643 18652 2688 18680
rect 2682 18640 2688 18652
rect 2740 18640 2746 18692
rect 2884 18680 2912 18720
rect 2961 18717 2973 18751
rect 3007 18748 3019 18751
rect 3602 18748 3608 18760
rect 3007 18720 3608 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 5368 18748 5396 18856
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 7558 18844 7564 18896
rect 7616 18884 7622 18896
rect 13906 18893 13912 18896
rect 11609 18887 11667 18893
rect 7616 18856 10364 18884
rect 7616 18844 7622 18856
rect 5442 18776 5448 18828
rect 5500 18816 5506 18828
rect 5997 18819 6055 18825
rect 5997 18816 6009 18819
rect 5500 18788 6009 18816
rect 5500 18776 5506 18788
rect 5997 18785 6009 18788
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 6454 18776 6460 18828
rect 6512 18816 6518 18828
rect 6549 18819 6607 18825
rect 6549 18816 6561 18819
rect 6512 18788 6561 18816
rect 6512 18776 6518 18788
rect 6549 18785 6561 18788
rect 6595 18785 6607 18819
rect 6549 18779 6607 18785
rect 6638 18776 6644 18828
rect 6696 18816 6702 18828
rect 8294 18816 8300 18828
rect 6696 18788 8300 18816
rect 6696 18776 6702 18788
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 9674 18816 9680 18828
rect 8444 18788 8489 18816
rect 9635 18788 9680 18816
rect 8444 18776 8450 18788
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10336 18816 10364 18856
rect 11609 18853 11621 18887
rect 11655 18884 11667 18887
rect 13900 18884 13912 18893
rect 11655 18856 12388 18884
rect 13867 18856 13912 18884
rect 11655 18853 11667 18856
rect 11609 18847 11667 18853
rect 10594 18816 10600 18828
rect 10336 18788 10600 18816
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 11054 18816 11060 18828
rect 11015 18788 11060 18816
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 12066 18816 12072 18828
rect 11256 18788 12072 18816
rect 8846 18748 8852 18760
rect 5368 18720 8852 18748
rect 8846 18708 8852 18720
rect 8904 18708 8910 18760
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9398 18748 9404 18760
rect 9359 18720 9404 18748
rect 9217 18711 9275 18717
rect 3053 18683 3111 18689
rect 3053 18680 3065 18683
rect 2884 18652 3065 18680
rect 3053 18649 3065 18652
rect 3099 18649 3111 18683
rect 3053 18643 3111 18649
rect 1489 18615 1547 18621
rect 1489 18581 1501 18615
rect 1535 18612 1547 18615
rect 1578 18612 1584 18624
rect 1535 18584 1584 18612
rect 1535 18581 1547 18584
rect 1489 18575 1547 18581
rect 1578 18572 1584 18584
rect 1636 18612 1642 18624
rect 2774 18612 2780 18624
rect 1636 18584 2780 18612
rect 1636 18572 1642 18584
rect 2774 18572 2780 18584
rect 2832 18572 2838 18624
rect 3068 18612 3096 18643
rect 3510 18640 3516 18692
rect 3568 18680 3574 18692
rect 3881 18683 3939 18689
rect 3881 18680 3893 18683
rect 3568 18652 3893 18680
rect 3568 18640 3574 18652
rect 3881 18649 3893 18652
rect 3927 18680 3939 18683
rect 6638 18680 6644 18692
rect 3927 18652 6644 18680
rect 3927 18649 3939 18652
rect 3881 18643 3939 18649
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 8297 18683 8355 18689
rect 8297 18649 8309 18683
rect 8343 18680 8355 18683
rect 8754 18680 8760 18692
rect 8343 18652 8760 18680
rect 8343 18649 8355 18652
rect 8297 18643 8355 18649
rect 8754 18640 8760 18652
rect 8812 18680 8818 18692
rect 9232 18680 9260 18711
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 9950 18748 9956 18760
rect 9911 18720 9956 18748
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 11256 18748 11284 18788
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 12360 18816 12388 18856
rect 13900 18847 13912 18856
rect 13906 18844 13912 18847
rect 13964 18844 13970 18896
rect 14458 18844 14464 18896
rect 14516 18884 14522 18896
rect 15749 18887 15807 18893
rect 15749 18884 15761 18887
rect 14516 18856 15761 18884
rect 14516 18844 14522 18856
rect 15749 18853 15761 18856
rect 15795 18853 15807 18887
rect 16393 18887 16451 18893
rect 15749 18847 15807 18853
rect 15856 18856 16252 18884
rect 12894 18816 12900 18828
rect 12360 18788 12756 18816
rect 12855 18788 12900 18816
rect 10612 18720 11284 18748
rect 8812 18652 9260 18680
rect 8812 18640 8818 18652
rect 9582 18640 9588 18692
rect 9640 18680 9646 18692
rect 10612 18680 10640 18720
rect 11330 18708 11336 18760
rect 11388 18748 11394 18760
rect 11388 18720 11433 18748
rect 11388 18708 11394 18720
rect 11974 18708 11980 18760
rect 12032 18748 12038 18760
rect 12161 18751 12219 18757
rect 12161 18748 12173 18751
rect 12032 18720 12173 18748
rect 12032 18708 12038 18720
rect 12161 18717 12173 18720
rect 12207 18717 12219 18751
rect 12342 18748 12348 18760
rect 12303 18720 12348 18748
rect 12161 18711 12219 18717
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 12728 18748 12756 18788
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 14182 18816 14188 18828
rect 13679 18788 14188 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 14642 18776 14648 18828
rect 14700 18816 14706 18828
rect 15657 18819 15715 18825
rect 15657 18816 15669 18819
rect 14700 18788 15669 18816
rect 14700 18776 14706 18788
rect 15657 18785 15669 18788
rect 15703 18816 15715 18819
rect 15856 18816 15884 18856
rect 15703 18788 15884 18816
rect 16117 18819 16175 18825
rect 15703 18785 15715 18788
rect 15657 18779 15715 18785
rect 16117 18785 16129 18819
rect 16163 18785 16175 18819
rect 16224 18816 16252 18856
rect 16393 18853 16405 18887
rect 16439 18884 16451 18887
rect 17402 18884 17408 18896
rect 16439 18856 17408 18884
rect 16439 18853 16451 18856
rect 16393 18847 16451 18853
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 18248 18884 18276 18915
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19484 18924 19809 18952
rect 19484 18912 19490 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 21082 18952 21088 18964
rect 21043 18924 21088 18952
rect 19797 18915 19855 18921
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 21453 18955 21511 18961
rect 21453 18921 21465 18955
rect 21499 18952 21511 18955
rect 21542 18952 21548 18964
rect 21499 18924 21548 18952
rect 21499 18921 21511 18924
rect 21453 18915 21511 18921
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 18598 18893 18604 18896
rect 18592 18884 18604 18893
rect 18248 18856 18604 18884
rect 18592 18847 18604 18856
rect 18598 18844 18604 18847
rect 18656 18844 18662 18896
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 20257 18887 20315 18893
rect 20257 18884 20269 18887
rect 19300 18856 20269 18884
rect 19300 18844 19306 18856
rect 20257 18853 20269 18856
rect 20303 18853 20315 18887
rect 20257 18847 20315 18853
rect 16758 18816 16764 18828
rect 16224 18788 16764 18816
rect 16117 18779 16175 18785
rect 12986 18748 12992 18760
rect 12728 18720 12992 18748
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 13078 18708 13084 18760
rect 13136 18748 13142 18760
rect 15838 18748 15844 18760
rect 13136 18720 13181 18748
rect 15799 18720 15844 18748
rect 13136 18708 13142 18720
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 9640 18652 10640 18680
rect 10689 18683 10747 18689
rect 9640 18640 9646 18652
rect 10689 18649 10701 18683
rect 10735 18680 10747 18683
rect 12526 18680 12532 18692
rect 10735 18652 12388 18680
rect 12487 18652 12532 18680
rect 10735 18649 10747 18652
rect 10689 18643 10747 18649
rect 5994 18612 6000 18624
rect 3068 18584 6000 18612
rect 5994 18572 6000 18584
rect 6052 18572 6058 18624
rect 6178 18612 6184 18624
rect 6139 18584 6184 18612
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 6656 18612 6684 18640
rect 8478 18612 8484 18624
rect 6656 18584 8484 18612
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 8573 18615 8631 18621
rect 8573 18581 8585 18615
rect 8619 18612 8631 18615
rect 11698 18612 11704 18624
rect 8619 18584 11704 18612
rect 8619 18581 8631 18584
rect 8573 18575 8631 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12360 18612 12388 18652
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 15013 18683 15071 18689
rect 15013 18649 15025 18683
rect 15059 18680 15071 18683
rect 15856 18680 15884 18708
rect 15059 18652 15884 18680
rect 15059 18649 15071 18652
rect 15013 18643 15071 18649
rect 16132 18612 16160 18779
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 17120 18819 17178 18825
rect 17120 18785 17132 18819
rect 17166 18816 17178 18819
rect 17494 18816 17500 18828
rect 17166 18788 17500 18816
rect 17166 18785 17178 18788
rect 17120 18779 17178 18785
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 20162 18816 20168 18828
rect 20123 18788 20168 18816
rect 20162 18776 20168 18788
rect 20220 18776 20226 18828
rect 20438 18816 20444 18828
rect 20272 18788 20444 18816
rect 16666 18708 16672 18760
rect 16724 18748 16730 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16724 18720 16865 18748
rect 16724 18708 16730 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 16758 18612 16764 18624
rect 12360 18584 16160 18612
rect 16719 18584 16764 18612
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 16868 18612 16896 18711
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 17920 18720 18337 18748
rect 17920 18708 17926 18720
rect 18325 18717 18337 18720
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 20272 18748 20300 18788
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 20898 18816 20904 18828
rect 20859 18788 20904 18816
rect 20898 18776 20904 18788
rect 20956 18776 20962 18828
rect 21269 18819 21327 18825
rect 21269 18785 21281 18819
rect 21315 18816 21327 18819
rect 21358 18816 21364 18828
rect 21315 18788 21364 18816
rect 21315 18785 21327 18788
rect 21269 18779 21327 18785
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 19484 18720 20300 18748
rect 20349 18751 20407 18757
rect 19484 18708 19490 18720
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 17880 18612 17908 18708
rect 19702 18680 19708 18692
rect 19663 18652 19708 18680
rect 19702 18640 19708 18652
rect 19760 18680 19766 18692
rect 20364 18680 20392 18711
rect 19760 18652 20392 18680
rect 19760 18640 19766 18652
rect 16868 18584 17908 18612
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 20714 18612 20720 18624
rect 18196 18584 20720 18612
rect 18196 18572 18202 18584
rect 20714 18572 20720 18584
rect 20772 18612 20778 18624
rect 21726 18612 21732 18624
rect 20772 18584 21732 18612
rect 20772 18572 20778 18584
rect 21726 18572 21732 18584
rect 21784 18572 21790 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2866 18368 2872 18420
rect 2924 18408 2930 18420
rect 3418 18408 3424 18420
rect 2924 18380 3424 18408
rect 2924 18368 2930 18380
rect 3418 18368 3424 18380
rect 3476 18368 3482 18420
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 10410 18408 10416 18420
rect 5776 18380 10416 18408
rect 5776 18368 5782 18380
rect 10410 18368 10416 18380
rect 10468 18368 10474 18420
rect 13906 18408 13912 18420
rect 10520 18380 12388 18408
rect 13819 18380 13912 18408
rect 1026 18300 1032 18352
rect 1084 18340 1090 18352
rect 8110 18340 8116 18352
rect 1084 18312 8116 18340
rect 1084 18300 1090 18312
rect 8110 18300 8116 18312
rect 8168 18300 8174 18352
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 9582 18340 9588 18352
rect 8352 18312 9588 18340
rect 8352 18300 8358 18312
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 9950 18300 9956 18352
rect 10008 18340 10014 18352
rect 10520 18340 10548 18380
rect 10008 18312 10548 18340
rect 12069 18343 12127 18349
rect 10008 18300 10014 18312
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 12250 18340 12256 18352
rect 12115 18312 12256 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 12360 18340 12388 18380
rect 13906 18368 13912 18380
rect 13964 18408 13970 18420
rect 14366 18408 14372 18420
rect 13964 18380 14372 18408
rect 13964 18368 13970 18380
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 15562 18408 15568 18420
rect 14516 18380 14561 18408
rect 14660 18380 15568 18408
rect 14516 18368 14522 18380
rect 14660 18340 14688 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 16022 18408 16028 18420
rect 15983 18380 16028 18408
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 17494 18408 17500 18420
rect 17455 18380 17500 18408
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 18046 18408 18052 18420
rect 18007 18380 18052 18408
rect 18046 18368 18052 18380
rect 18104 18368 18110 18420
rect 18690 18368 18696 18420
rect 18748 18408 18754 18420
rect 19242 18408 19248 18420
rect 18748 18380 19248 18408
rect 18748 18368 18754 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19521 18411 19579 18417
rect 19521 18408 19533 18411
rect 19392 18380 19533 18408
rect 19392 18368 19398 18380
rect 19521 18377 19533 18380
rect 19567 18377 19579 18411
rect 20990 18408 20996 18420
rect 20951 18380 20996 18408
rect 19521 18371 19579 18377
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 12360 18312 14688 18340
rect 17126 18300 17132 18352
rect 17184 18340 17190 18352
rect 21177 18343 21235 18349
rect 21177 18340 21189 18343
rect 17184 18312 21189 18340
rect 17184 18300 17190 18312
rect 21177 18309 21189 18312
rect 21223 18340 21235 18343
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21223 18312 22017 18340
rect 21223 18309 21235 18312
rect 21177 18303 21235 18309
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22005 18303 22063 18309
rect 1394 18232 1400 18284
rect 1452 18272 1458 18284
rect 1452 18244 2544 18272
rect 1452 18232 1458 18244
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18204 1823 18207
rect 2516 18204 2544 18244
rect 2590 18232 2596 18284
rect 2648 18272 2654 18284
rect 5442 18272 5448 18284
rect 2648 18244 5304 18272
rect 5403 18244 5448 18272
rect 2648 18232 2654 18244
rect 2958 18204 2964 18216
rect 1811 18176 2268 18204
rect 2516 18176 2964 18204
rect 1811 18173 1823 18176
rect 1765 18167 1823 18173
rect 2240 18077 2268 18176
rect 2958 18164 2964 18176
rect 3016 18164 3022 18216
rect 4154 18204 4160 18216
rect 3252 18176 4160 18204
rect 2225 18071 2283 18077
rect 2225 18037 2237 18071
rect 2271 18068 2283 18071
rect 2314 18068 2320 18080
rect 2271 18040 2320 18068
rect 2271 18037 2283 18040
rect 2225 18031 2283 18037
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 2498 18028 2504 18080
rect 2556 18068 2562 18080
rect 2593 18071 2651 18077
rect 2593 18068 2605 18071
rect 2556 18040 2605 18068
rect 2556 18028 2562 18040
rect 2593 18037 2605 18040
rect 2639 18068 2651 18071
rect 3252 18068 3280 18176
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 5166 18204 5172 18216
rect 5127 18176 5172 18204
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 5276 18204 5304 18244
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 7466 18272 7472 18284
rect 6604 18244 7472 18272
rect 6604 18232 6610 18244
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 7558 18232 7564 18284
rect 7616 18272 7622 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7616 18244 7849 18272
rect 7616 18232 7622 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 8386 18272 8392 18284
rect 8347 18244 8392 18272
rect 7837 18235 7895 18241
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 10134 18272 10140 18284
rect 8536 18244 10140 18272
rect 8536 18232 8542 18244
rect 10134 18232 10140 18244
rect 10192 18232 10198 18284
rect 11698 18232 11704 18284
rect 11756 18232 11762 18284
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18272 12495 18275
rect 12894 18272 12900 18284
rect 12483 18244 12900 18272
rect 12483 18241 12495 18244
rect 12437 18235 12495 18241
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 16022 18232 16028 18284
rect 16080 18272 16086 18284
rect 16080 18244 16252 18272
rect 16080 18232 16086 18244
rect 6822 18204 6828 18216
rect 5276 18176 6828 18204
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 8113 18207 8171 18213
rect 8113 18204 8125 18207
rect 6972 18176 8125 18204
rect 6972 18164 6978 18176
rect 8113 18173 8125 18176
rect 8159 18173 8171 18207
rect 8113 18167 8171 18173
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 10956 18207 11014 18213
rect 10956 18173 10968 18207
rect 11002 18204 11014 18207
rect 11238 18204 11244 18216
rect 11002 18176 11244 18204
rect 11002 18173 11014 18176
rect 10956 18167 11014 18173
rect 3326 18096 3332 18148
rect 3384 18136 3390 18148
rect 4890 18136 4896 18148
rect 3384 18108 4896 18136
rect 3384 18096 3390 18108
rect 4890 18096 4896 18108
rect 4948 18096 4954 18148
rect 2639 18040 3280 18068
rect 2639 18037 2651 18040
rect 2593 18031 2651 18037
rect 3694 18028 3700 18080
rect 3752 18068 3758 18080
rect 6730 18068 6736 18080
rect 3752 18040 6736 18068
rect 3752 18028 3758 18040
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 7282 18068 7288 18080
rect 7243 18040 7288 18068
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7650 18068 7656 18080
rect 7611 18040 7656 18068
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 7745 18071 7803 18077
rect 7745 18037 7757 18071
rect 7791 18068 7803 18071
rect 8386 18068 8392 18080
rect 7791 18040 8392 18068
rect 7791 18037 7803 18040
rect 7745 18031 7803 18037
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 8662 18028 8668 18080
rect 8720 18068 8726 18080
rect 10134 18068 10140 18080
rect 8720 18040 10140 18068
rect 8720 18028 8726 18040
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10704 18068 10732 18167
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 11716 18204 11744 18232
rect 14090 18204 14096 18216
rect 11716 18176 14096 18204
rect 14090 18164 14096 18176
rect 14148 18164 14154 18216
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14645 18207 14703 18213
rect 14645 18204 14657 18207
rect 14240 18176 14657 18204
rect 14240 18164 14246 18176
rect 14645 18173 14657 18176
rect 14691 18204 14703 18207
rect 14734 18204 14740 18216
rect 14691 18176 14740 18204
rect 14691 18173 14703 18176
rect 14645 18167 14703 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 14912 18207 14970 18213
rect 14912 18173 14924 18207
rect 14958 18204 14970 18207
rect 15838 18204 15844 18216
rect 14958 18176 15844 18204
rect 14958 18173 14970 18176
rect 14912 18167 14970 18173
rect 15838 18164 15844 18176
rect 15896 18164 15902 18216
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18173 16175 18207
rect 16224 18204 16252 18244
rect 17494 18232 17500 18284
rect 17552 18272 17558 18284
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 17552 18244 18613 18272
rect 17552 18232 17558 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 20073 18275 20131 18281
rect 20073 18272 20085 18275
rect 19760 18244 20085 18272
rect 19760 18232 19766 18244
rect 20073 18241 20085 18244
rect 20119 18241 20131 18275
rect 20073 18235 20131 18241
rect 16373 18207 16431 18213
rect 16373 18204 16385 18207
rect 16224 18176 16385 18204
rect 16117 18167 16175 18173
rect 16373 18173 16385 18176
rect 16419 18173 16431 18207
rect 16373 18167 16431 18173
rect 18524 18176 20484 18204
rect 11698 18096 11704 18148
rect 11756 18136 11762 18148
rect 11974 18136 11980 18148
rect 11756 18108 11980 18136
rect 11756 18096 11762 18108
rect 11974 18096 11980 18108
rect 12032 18136 12038 18148
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 12032 18108 12173 18136
rect 12032 18096 12038 18108
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 16132 18136 16160 18167
rect 16666 18136 16672 18148
rect 16132 18108 16672 18136
rect 12161 18099 12219 18105
rect 16666 18096 16672 18108
rect 16724 18096 16730 18148
rect 17589 18139 17647 18145
rect 17589 18105 17601 18139
rect 17635 18136 17647 18139
rect 18417 18139 18475 18145
rect 18417 18136 18429 18139
rect 17635 18108 18429 18136
rect 17635 18105 17647 18108
rect 17589 18099 17647 18105
rect 18417 18105 18429 18108
rect 18463 18105 18475 18139
rect 18417 18099 18475 18105
rect 10870 18068 10876 18080
rect 10704 18040 10876 18068
rect 10870 18028 10876 18040
rect 10928 18068 10934 18080
rect 11790 18068 11796 18080
rect 10928 18040 11796 18068
rect 10928 18028 10934 18040
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 15746 18028 15752 18080
rect 15804 18068 15810 18080
rect 17678 18068 17684 18080
rect 15804 18040 17684 18068
rect 15804 18028 15810 18040
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 18524 18077 18552 18176
rect 19889 18139 19947 18145
rect 19889 18105 19901 18139
rect 19935 18136 19947 18139
rect 20349 18139 20407 18145
rect 20349 18136 20361 18139
rect 19935 18108 20361 18136
rect 19935 18105 19947 18108
rect 19889 18099 19947 18105
rect 20349 18105 20361 18108
rect 20395 18105 20407 18139
rect 20456 18136 20484 18176
rect 20714 18164 20720 18216
rect 20772 18204 20778 18216
rect 20809 18207 20867 18213
rect 20809 18204 20821 18207
rect 20772 18176 20821 18204
rect 20772 18164 20778 18176
rect 20809 18173 20821 18176
rect 20855 18173 20867 18207
rect 20809 18167 20867 18173
rect 20898 18136 20904 18148
rect 20456 18108 20904 18136
rect 20349 18099 20407 18105
rect 20898 18096 20904 18108
rect 20956 18136 20962 18148
rect 21361 18139 21419 18145
rect 21361 18136 21373 18139
rect 20956 18108 21373 18136
rect 20956 18096 20962 18108
rect 21361 18105 21373 18108
rect 21407 18105 21419 18139
rect 21361 18099 21419 18105
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 18104 18040 18521 18068
rect 18104 18028 18110 18040
rect 18509 18037 18521 18040
rect 18555 18037 18567 18071
rect 18509 18031 18567 18037
rect 19429 18071 19487 18077
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19475 18040 19993 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 19981 18037 19993 18040
rect 20027 18068 20039 18071
rect 20530 18068 20536 18080
rect 20027 18040 20536 18068
rect 20027 18037 20039 18040
rect 19981 18031 20039 18037
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 20714 18068 20720 18080
rect 20675 18040 20720 18068
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 4341 17867 4399 17873
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 5166 17864 5172 17876
rect 4387 17836 5172 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 6733 17867 6791 17873
rect 6733 17833 6745 17867
rect 6779 17864 6791 17867
rect 6914 17864 6920 17876
rect 6779 17836 6920 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7193 17867 7251 17873
rect 7193 17833 7205 17867
rect 7239 17864 7251 17867
rect 7282 17864 7288 17876
rect 7239 17836 7288 17864
rect 7239 17833 7251 17836
rect 7193 17827 7251 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 7561 17867 7619 17873
rect 7561 17833 7573 17867
rect 7607 17864 7619 17867
rect 7650 17864 7656 17876
rect 7607 17836 7656 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 8202 17824 8208 17876
rect 8260 17864 8266 17876
rect 8389 17867 8447 17873
rect 8389 17864 8401 17867
rect 8260 17836 8401 17864
rect 8260 17824 8266 17836
rect 8389 17833 8401 17836
rect 8435 17833 8447 17867
rect 8389 17827 8447 17833
rect 8665 17867 8723 17873
rect 8665 17833 8677 17867
rect 8711 17864 8723 17867
rect 8846 17864 8852 17876
rect 8711 17836 8852 17864
rect 8711 17833 8723 17836
rect 8665 17827 8723 17833
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 9306 17864 9312 17876
rect 9267 17836 9312 17864
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11241 17867 11299 17873
rect 11241 17864 11253 17867
rect 11112 17836 11253 17864
rect 11112 17824 11118 17836
rect 11241 17833 11253 17836
rect 11287 17833 11299 17867
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 11241 17827 11299 17833
rect 11348 17836 13001 17864
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2593 17799 2651 17805
rect 2593 17796 2605 17799
rect 1820 17768 2605 17796
rect 1820 17756 1826 17768
rect 2593 17765 2605 17768
rect 2639 17765 2651 17799
rect 2593 17759 2651 17765
rect 4709 17799 4767 17805
rect 4709 17765 4721 17799
rect 4755 17796 4767 17799
rect 5534 17796 5540 17808
rect 4755 17768 5540 17796
rect 4755 17765 4767 17768
rect 4709 17759 4767 17765
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 8021 17799 8079 17805
rect 8021 17796 8033 17799
rect 6880 17768 8033 17796
rect 6880 17756 6886 17768
rect 8021 17765 8033 17768
rect 8067 17796 8079 17799
rect 8757 17799 8815 17805
rect 8757 17796 8769 17799
rect 8067 17768 8769 17796
rect 8067 17765 8079 17768
rect 8021 17759 8079 17765
rect 8757 17765 8769 17768
rect 8803 17796 8815 17799
rect 11348 17796 11376 17836
rect 12989 17833 13001 17836
rect 13035 17864 13047 17867
rect 13906 17864 13912 17876
rect 13035 17836 13912 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 15289 17867 15347 17873
rect 15289 17833 15301 17867
rect 15335 17864 15347 17867
rect 15378 17864 15384 17876
rect 15335 17836 15384 17864
rect 15335 17833 15347 17836
rect 15289 17827 15347 17833
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 15746 17864 15752 17876
rect 15707 17836 15752 17864
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 16945 17867 17003 17873
rect 16945 17833 16957 17867
rect 16991 17864 17003 17867
rect 17954 17864 17960 17876
rect 16991 17836 17960 17864
rect 16991 17833 17003 17836
rect 16945 17827 17003 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 21082 17864 21088 17876
rect 21043 17836 21088 17864
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 8803 17768 11376 17796
rect 11701 17799 11759 17805
rect 8803 17765 8815 17768
rect 8757 17759 8815 17765
rect 11701 17765 11713 17799
rect 11747 17796 11759 17799
rect 12529 17799 12587 17805
rect 12529 17796 12541 17799
rect 11747 17768 12541 17796
rect 11747 17765 11759 17768
rect 11701 17759 11759 17765
rect 12529 17765 12541 17768
rect 12575 17765 12587 17799
rect 12529 17759 12587 17765
rect 15105 17799 15163 17805
rect 15105 17765 15117 17799
rect 15151 17796 15163 17799
rect 15764 17796 15792 17824
rect 15151 17768 15792 17796
rect 17313 17799 17371 17805
rect 15151 17765 15163 17768
rect 15105 17759 15163 17765
rect 17313 17765 17325 17799
rect 17359 17796 17371 17799
rect 17402 17796 17408 17808
rect 17359 17768 17408 17796
rect 17359 17765 17371 17768
rect 17313 17759 17371 17765
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 17678 17756 17684 17808
rect 17736 17796 17742 17808
rect 18782 17796 18788 17808
rect 17736 17768 18788 17796
rect 17736 17756 17742 17768
rect 18782 17756 18788 17768
rect 18840 17796 18846 17808
rect 19978 17796 19984 17808
rect 18840 17768 19984 17796
rect 18840 17756 18846 17768
rect 19978 17756 19984 17768
rect 20036 17756 20042 17808
rect 20073 17799 20131 17805
rect 20073 17765 20085 17799
rect 20119 17796 20131 17799
rect 22005 17799 22063 17805
rect 22005 17796 22017 17799
rect 20119 17768 22017 17796
rect 20119 17765 20131 17768
rect 20073 17759 20131 17765
rect 22005 17765 22017 17768
rect 22051 17765 22063 17799
rect 22005 17759 22063 17765
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17697 2375 17731
rect 5436 17731 5494 17737
rect 5436 17728 5448 17731
rect 2317 17691 2375 17697
rect 4908 17700 5448 17728
rect 2332 17592 2360 17691
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4908 17669 4936 17700
rect 5436 17697 5448 17700
rect 5482 17728 5494 17731
rect 5994 17728 6000 17740
rect 5482 17700 6000 17728
rect 5482 17697 5494 17700
rect 5436 17691 5494 17697
rect 5994 17688 6000 17700
rect 6052 17688 6058 17740
rect 6730 17688 6736 17740
rect 6788 17728 6794 17740
rect 7098 17728 7104 17740
rect 6788 17700 6960 17728
rect 7059 17700 7104 17728
rect 6788 17688 6794 17700
rect 4801 17663 4859 17669
rect 4801 17660 4813 17663
rect 4304 17632 4813 17660
rect 4304 17620 4310 17632
rect 4801 17629 4813 17632
rect 4847 17629 4859 17663
rect 4801 17623 4859 17629
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17629 4951 17663
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 4893 17623 4951 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6932 17660 6960 17700
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7300 17700 7941 17728
rect 7300 17660 7328 17700
rect 7929 17697 7941 17700
rect 7975 17728 7987 17731
rect 8941 17731 8999 17737
rect 8941 17728 8953 17731
rect 7975 17700 8953 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 8941 17697 8953 17700
rect 8987 17697 8999 17731
rect 8941 17691 8999 17697
rect 10036 17731 10094 17737
rect 10036 17697 10048 17731
rect 10082 17728 10094 17731
rect 10870 17728 10876 17740
rect 10082 17700 10876 17728
rect 10082 17697 10094 17700
rect 10036 17691 10094 17697
rect 6932 17632 7328 17660
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17660 7435 17663
rect 7834 17660 7840 17672
rect 7423 17632 7840 17660
rect 7423 17629 7435 17632
rect 7377 17623 7435 17629
rect 7834 17620 7840 17632
rect 7892 17620 7898 17672
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 8128 17592 8156 17623
rect 8478 17592 8484 17604
rect 2332 17564 4936 17592
rect 2314 17484 2320 17536
rect 2372 17524 2378 17536
rect 4798 17524 4804 17536
rect 2372 17496 4804 17524
rect 2372 17484 2378 17496
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 4908 17524 4936 17564
rect 6564 17564 8484 17592
rect 6362 17524 6368 17536
rect 4908 17496 6368 17524
rect 6362 17484 6368 17496
rect 6420 17484 6426 17536
rect 6454 17484 6460 17536
rect 6512 17524 6518 17536
rect 6564 17533 6592 17564
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 8956 17592 8984 17691
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 11609 17731 11667 17737
rect 11609 17697 11621 17731
rect 11655 17728 11667 17731
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11655 17700 12081 17728
rect 11655 17697 11667 17700
rect 11609 17691 11667 17697
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 14458 17728 14464 17740
rect 12069 17691 12127 17697
rect 12176 17700 14464 17728
rect 9766 17660 9772 17672
rect 9727 17632 9772 17660
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 10888 17660 10916 17688
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 10888 17632 11805 17660
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11149 17595 11207 17601
rect 8956 17564 9812 17592
rect 6549 17527 6607 17533
rect 6549 17524 6561 17527
rect 6512 17496 6561 17524
rect 6512 17484 6518 17496
rect 6549 17493 6561 17496
rect 6595 17493 6607 17527
rect 6549 17487 6607 17493
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 7432 17496 9137 17524
rect 7432 17484 7438 17496
rect 9125 17493 9137 17496
rect 9171 17524 9183 17527
rect 9674 17524 9680 17536
rect 9171 17496 9680 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 9784 17524 9812 17564
rect 11149 17561 11161 17595
rect 11195 17592 11207 17595
rect 11238 17592 11244 17604
rect 11195 17564 11244 17592
rect 11195 17561 11207 17564
rect 11149 17555 11207 17561
rect 11238 17552 11244 17564
rect 11296 17552 11302 17604
rect 11808 17592 11836 17623
rect 11974 17620 11980 17672
rect 12032 17660 12038 17672
rect 12176 17660 12204 17700
rect 14458 17688 14464 17700
rect 14516 17688 14522 17740
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 16117 17731 16175 17737
rect 16117 17728 16129 17731
rect 15703 17700 16129 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 16117 17697 16129 17700
rect 16163 17697 16175 17731
rect 16117 17691 16175 17697
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17728 19671 17731
rect 20165 17731 20223 17737
rect 20165 17728 20177 17731
rect 19659 17700 20177 17728
rect 19659 17697 19671 17700
rect 19613 17691 19671 17697
rect 20165 17697 20177 17700
rect 20211 17728 20223 17731
rect 20254 17728 20260 17740
rect 20211 17700 20260 17728
rect 20211 17697 20223 17700
rect 20165 17691 20223 17697
rect 20254 17688 20260 17700
rect 20312 17728 20318 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20312 17700 20913 17728
rect 20312 17688 20318 17700
rect 20901 17697 20913 17700
rect 20947 17728 20959 17731
rect 21453 17731 21511 17737
rect 21453 17728 21465 17731
rect 20947 17700 21465 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21453 17697 21465 17700
rect 21499 17697 21511 17731
rect 21453 17691 21511 17697
rect 12032 17632 12204 17660
rect 12437 17663 12495 17669
rect 12032 17620 12038 17632
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 12483 17632 12541 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 12529 17629 12541 17632
rect 12575 17660 12587 17663
rect 12986 17660 12992 17672
rect 12575 17632 12992 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 12986 17620 12992 17632
rect 13044 17660 13050 17672
rect 15470 17660 15476 17672
rect 13044 17632 15476 17660
rect 13044 17620 13050 17632
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 13538 17592 13544 17604
rect 11808 17564 13544 17592
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 13630 17552 13636 17604
rect 13688 17592 13694 17604
rect 16761 17595 16819 17601
rect 16761 17592 16773 17595
rect 13688 17564 16773 17592
rect 13688 17552 13694 17564
rect 16761 17561 16773 17564
rect 16807 17592 16819 17595
rect 17420 17592 17448 17623
rect 17494 17620 17500 17672
rect 17552 17660 17558 17672
rect 20346 17660 20352 17672
rect 17552 17632 17597 17660
rect 20307 17632 20352 17660
rect 17552 17620 17558 17632
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 18049 17595 18107 17601
rect 18049 17592 18061 17595
rect 16807 17564 17448 17592
rect 17512 17564 18061 17592
rect 16807 17561 16819 17564
rect 16761 17555 16819 17561
rect 11974 17524 11980 17536
rect 9784 17496 11980 17524
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12768 17496 12817 17524
rect 12768 17484 12774 17496
rect 12805 17493 12817 17496
rect 12851 17524 12863 17527
rect 13446 17524 13452 17536
rect 12851 17496 13452 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 17512 17524 17540 17564
rect 18049 17561 18061 17564
rect 18095 17561 18107 17595
rect 18049 17555 18107 17561
rect 20530 17552 20536 17604
rect 20588 17592 20594 17604
rect 20588 17564 21128 17592
rect 20588 17552 20594 17564
rect 21100 17536 21128 17564
rect 17862 17524 17868 17536
rect 17460 17496 17540 17524
rect 17823 17496 17868 17524
rect 17460 17484 17466 17496
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 19702 17524 19708 17536
rect 19663 17496 19708 17524
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 20162 17484 20168 17536
rect 20220 17524 20226 17536
rect 20625 17527 20683 17533
rect 20625 17524 20637 17527
rect 20220 17496 20637 17524
rect 20220 17484 20226 17496
rect 20625 17493 20637 17496
rect 20671 17493 20683 17527
rect 20625 17487 20683 17493
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 21269 17527 21327 17533
rect 21269 17524 21281 17527
rect 21140 17496 21281 17524
rect 21140 17484 21146 17496
rect 21269 17493 21281 17496
rect 21315 17524 21327 17527
rect 21358 17524 21364 17536
rect 21315 17496 21364 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 21358 17484 21364 17496
rect 21416 17484 21422 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2317 17323 2375 17329
rect 2317 17289 2329 17323
rect 2363 17320 2375 17323
rect 2682 17320 2688 17332
rect 2363 17292 2688 17320
rect 2363 17289 2375 17292
rect 2317 17283 2375 17289
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 2958 17280 2964 17332
rect 3016 17320 3022 17332
rect 5994 17320 6000 17332
rect 3016 17292 5856 17320
rect 5955 17292 6000 17320
rect 3016 17280 3022 17292
rect 4522 17252 4528 17264
rect 4483 17224 4528 17252
rect 4522 17212 4528 17224
rect 4580 17212 4586 17264
rect 2682 17184 2688 17196
rect 2148 17156 2688 17184
rect 2148 17125 2176 17156
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 2774 17144 2780 17196
rect 2832 17184 2838 17196
rect 2958 17184 2964 17196
rect 2832 17156 2964 17184
rect 2832 17144 2838 17156
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 5828 17184 5856 17292
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 8294 17320 8300 17332
rect 7892 17292 8300 17320
rect 7892 17280 7898 17292
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 8444 17292 8489 17320
rect 8444 17280 8450 17292
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 10042 17320 10048 17332
rect 9364 17292 10048 17320
rect 9364 17280 9370 17292
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 10321 17323 10379 17329
rect 10321 17289 10333 17323
rect 10367 17320 10379 17323
rect 11054 17320 11060 17332
rect 10367 17292 11060 17320
rect 10367 17289 10379 17292
rect 10321 17283 10379 17289
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11698 17320 11704 17332
rect 11256 17292 11704 17320
rect 8846 17212 8852 17264
rect 8904 17252 8910 17264
rect 11256 17252 11284 17292
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 12032 17292 12173 17320
rect 12032 17280 12038 17292
rect 12161 17289 12173 17292
rect 12207 17320 12219 17323
rect 12250 17320 12256 17332
rect 12207 17292 12256 17320
rect 12207 17289 12219 17292
rect 12161 17283 12219 17289
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 13538 17280 13544 17332
rect 13596 17320 13602 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 13596 17292 20545 17320
rect 13596 17280 13602 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 20990 17320 20996 17332
rect 20951 17292 20996 17320
rect 20533 17283 20591 17289
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 12710 17252 12716 17264
rect 8904 17224 11284 17252
rect 11348 17224 12716 17252
rect 8904 17212 8910 17224
rect 5828 17156 7052 17184
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 3142 17116 3148 17128
rect 3055 17088 3148 17116
rect 2133 17079 2191 17085
rect 1780 17048 1808 17079
rect 3142 17076 3148 17088
rect 3200 17116 3206 17128
rect 4617 17119 4675 17125
rect 4617 17116 4629 17119
rect 3200 17088 4629 17116
rect 3200 17076 3206 17088
rect 4617 17085 4629 17088
rect 4663 17116 4675 17119
rect 5166 17116 5172 17128
rect 4663 17088 5172 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 5166 17076 5172 17088
rect 5224 17116 5230 17128
rect 6178 17116 6184 17128
rect 5224 17088 6184 17116
rect 5224 17076 5230 17088
rect 6178 17076 6184 17088
rect 6236 17076 6242 17128
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17085 6975 17119
rect 7024 17116 7052 17156
rect 8478 17144 8484 17196
rect 8536 17184 8542 17196
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8536 17156 8953 17184
rect 8536 17144 8542 17156
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9858 17184 9864 17196
rect 9732 17156 9864 17184
rect 9732 17144 9738 17156
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 10008 17156 10057 17184
rect 10008 17144 10014 17156
rect 10045 17153 10057 17156
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 10410 17144 10416 17196
rect 10468 17184 10474 17196
rect 10686 17184 10692 17196
rect 10468 17156 10692 17184
rect 10468 17144 10474 17156
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 10870 17184 10876 17196
rect 10831 17156 10876 17184
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 9306 17116 9312 17128
rect 7024 17088 9312 17116
rect 6917 17079 6975 17085
rect 3412 17051 3470 17057
rect 1780 17020 2636 17048
rect 2608 16989 2636 17020
rect 3412 17017 3424 17051
rect 3458 17048 3470 17051
rect 3970 17048 3976 17060
rect 3458 17020 3976 17048
rect 3458 17017 3470 17020
rect 3412 17011 3470 17017
rect 3970 17008 3976 17020
rect 4028 17008 4034 17060
rect 4522 17008 4528 17060
rect 4580 17048 4586 17060
rect 4798 17048 4804 17060
rect 4580 17020 4804 17048
rect 4580 17008 4586 17020
rect 4798 17008 4804 17020
rect 4856 17057 4862 17060
rect 4856 17051 4920 17057
rect 4856 17017 4874 17051
rect 4908 17017 4920 17051
rect 6932 17048 6960 17079
rect 9306 17076 9312 17088
rect 9364 17116 9370 17128
rect 10781 17119 10839 17125
rect 10781 17116 10793 17119
rect 9364 17088 10793 17116
rect 9364 17076 9370 17088
rect 10781 17085 10793 17088
rect 10827 17085 10839 17119
rect 11348 17116 11376 17224
rect 12710 17212 12716 17224
rect 12768 17212 12774 17264
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 17862 17252 17868 17264
rect 16540 17224 17868 17252
rect 16540 17212 16546 17224
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 20714 17252 20720 17264
rect 20364 17224 20720 17252
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 12805 17187 12863 17193
rect 12805 17153 12817 17187
rect 12851 17184 12863 17187
rect 13170 17184 13176 17196
rect 12851 17156 13176 17184
rect 12851 17153 12863 17156
rect 12805 17147 12863 17153
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13596 17156 13645 17184
rect 13596 17144 13602 17156
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 14553 17187 14611 17193
rect 14553 17184 14565 17187
rect 13780 17156 14565 17184
rect 13780 17144 13786 17156
rect 14553 17153 14565 17156
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17184 14795 17187
rect 15197 17187 15255 17193
rect 14783 17156 15148 17184
rect 14783 17153 14795 17156
rect 14737 17147 14795 17153
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 10781 17079 10839 17085
rect 11256 17088 11376 17116
rect 11440 17088 12541 17116
rect 7006 17048 7012 17060
rect 6932 17020 7012 17048
rect 4856 17011 4920 17017
rect 4856 17008 4862 17011
rect 7006 17008 7012 17020
rect 7064 17008 7070 17060
rect 7184 17051 7242 17057
rect 7184 17017 7196 17051
rect 7230 17048 7242 17051
rect 7558 17048 7564 17060
rect 7230 17020 7564 17048
rect 7230 17017 7242 17020
rect 7184 17011 7242 17017
rect 7558 17008 7564 17020
rect 7616 17008 7622 17060
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 8849 17051 8907 17057
rect 8849 17048 8861 17051
rect 8260 17020 8861 17048
rect 8260 17008 8266 17020
rect 8849 17017 8861 17020
rect 8895 17048 8907 17051
rect 11256 17048 11284 17088
rect 11440 17048 11468 17088
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 12529 17079 12587 17085
rect 14108 17088 14933 17116
rect 8895 17020 11284 17048
rect 11348 17020 11468 17048
rect 11517 17051 11575 17057
rect 8895 17017 8907 17020
rect 8849 17011 8907 17017
rect 2593 16983 2651 16989
rect 2593 16949 2605 16983
rect 2639 16980 2651 16983
rect 6270 16980 6276 16992
rect 2639 16952 6276 16980
rect 2639 16949 2651 16952
rect 2593 16943 2651 16949
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 8754 16980 8760 16992
rect 8715 16952 8760 16980
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 9674 16980 9680 16992
rect 9539 16952 9680 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 9858 16980 9864 16992
rect 9819 16952 9864 16980
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 9953 16983 10011 16989
rect 9953 16949 9965 16983
rect 9999 16980 10011 16983
rect 10042 16980 10048 16992
rect 9999 16952 10048 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10376 16952 10701 16980
rect 10376 16940 10382 16952
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10689 16943 10747 16949
rect 11149 16983 11207 16989
rect 11149 16949 11161 16983
rect 11195 16980 11207 16983
rect 11348 16980 11376 17020
rect 11517 17017 11529 17051
rect 11563 17048 11575 17051
rect 11882 17048 11888 17060
rect 11563 17020 11888 17048
rect 11563 17017 11575 17020
rect 11517 17011 11575 17017
rect 11882 17008 11888 17020
rect 11940 17008 11946 17060
rect 12250 17008 12256 17060
rect 12308 17048 12314 17060
rect 13449 17051 13507 17057
rect 13449 17048 13461 17051
rect 12308 17020 13461 17048
rect 12308 17008 12314 17020
rect 13449 17017 13461 17020
rect 13495 17048 13507 17051
rect 13630 17048 13636 17060
rect 13495 17020 13636 17048
rect 13495 17017 13507 17020
rect 13449 17011 13507 17017
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 11195 16952 11376 16980
rect 11195 16949 11207 16952
rect 11149 16943 11207 16949
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11609 16983 11667 16989
rect 11609 16980 11621 16983
rect 11480 16952 11621 16980
rect 11480 16940 11486 16952
rect 11609 16949 11621 16952
rect 11655 16949 11667 16983
rect 11609 16943 11667 16949
rect 12069 16983 12127 16989
rect 12069 16949 12081 16983
rect 12115 16980 12127 16983
rect 12342 16980 12348 16992
rect 12115 16952 12348 16980
rect 12115 16949 12127 16952
rect 12069 16943 12127 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 13078 16980 13084 16992
rect 13039 16952 13084 16980
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 13541 16983 13599 16989
rect 13541 16949 13553 16983
rect 13587 16980 13599 16983
rect 13906 16980 13912 16992
rect 13587 16952 13912 16980
rect 13587 16949 13599 16952
rect 13541 16943 13599 16949
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14108 16989 14136 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 15120 17048 15148 17156
rect 15197 17153 15209 17187
rect 15243 17184 15255 17187
rect 15286 17184 15292 17196
rect 15243 17156 15292 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 17034 17144 17040 17196
rect 17092 17184 17098 17196
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 17092 17156 17417 17184
rect 17092 17144 17098 17156
rect 17405 17153 17417 17156
rect 17451 17153 17463 17187
rect 17405 17147 17463 17153
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17116 17279 17119
rect 18506 17116 18512 17128
rect 17267 17088 18512 17116
rect 17267 17085 17279 17088
rect 17221 17079 17279 17085
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 19150 17116 19156 17128
rect 19111 17088 19156 17116
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 20364 17116 20392 17224
rect 20714 17212 20720 17224
rect 20772 17212 20778 17264
rect 20714 17116 20720 17128
rect 19260 17088 20392 17116
rect 20627 17088 20720 17116
rect 15286 17048 15292 17060
rect 15120 17020 15292 17048
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 15470 17008 15476 17060
rect 15528 17048 15534 17060
rect 19260 17048 19288 17088
rect 20714 17076 20720 17088
rect 20772 17116 20778 17128
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 20772 17088 20821 17116
rect 20772 17076 20778 17088
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 15528 17020 19288 17048
rect 15528 17008 15534 17020
rect 19334 17008 19340 17060
rect 19392 17057 19398 17060
rect 19392 17051 19456 17057
rect 19392 17017 19410 17051
rect 19444 17017 19456 17051
rect 19392 17011 19456 17017
rect 19392 17008 19398 17011
rect 20530 17008 20536 17060
rect 20588 17048 20594 17060
rect 21361 17051 21419 17057
rect 21361 17048 21373 17051
rect 20588 17020 21373 17048
rect 20588 17008 20594 17020
rect 21361 17017 21373 17020
rect 21407 17017 21419 17051
rect 21361 17011 21419 17017
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16949 14151 16983
rect 14458 16980 14464 16992
rect 14419 16952 14464 16980
rect 14093 16943 14151 16949
rect 14458 16940 14464 16952
rect 14516 16940 14522 16992
rect 15562 16980 15568 16992
rect 15523 16952 15568 16980
rect 15562 16940 15568 16952
rect 15620 16980 15626 16992
rect 18966 16980 18972 16992
rect 15620 16952 18972 16980
rect 15620 16940 15626 16952
rect 18966 16940 18972 16952
rect 19024 16980 19030 16992
rect 20898 16980 20904 16992
rect 19024 16952 20904 16980
rect 19024 16940 19030 16952
rect 20898 16940 20904 16952
rect 20956 16980 20962 16992
rect 21177 16983 21235 16989
rect 21177 16980 21189 16983
rect 20956 16952 21189 16980
rect 20956 16940 20962 16952
rect 21177 16949 21189 16952
rect 21223 16949 21235 16983
rect 21177 16943 21235 16949
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 3053 16779 3111 16785
rect 2832 16748 2877 16776
rect 2832 16736 2838 16748
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 3099 16748 4537 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 5353 16779 5411 16785
rect 5353 16776 5365 16779
rect 4948 16748 5365 16776
rect 4948 16736 4954 16748
rect 5353 16745 5365 16748
rect 5399 16776 5411 16779
rect 5905 16779 5963 16785
rect 5905 16776 5917 16779
rect 5399 16748 5917 16776
rect 5399 16745 5411 16748
rect 5353 16739 5411 16745
rect 5905 16745 5917 16748
rect 5951 16776 5963 16779
rect 7374 16776 7380 16788
rect 5951 16748 7380 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 7558 16776 7564 16788
rect 7519 16748 7564 16776
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 9858 16776 9864 16788
rect 7659 16748 9864 16776
rect 7659 16708 7687 16748
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 12897 16779 12955 16785
rect 12124 16748 12388 16776
rect 12124 16736 12130 16748
rect 4080 16680 7687 16708
rect 3050 16600 3056 16652
rect 3108 16640 3114 16652
rect 3421 16643 3479 16649
rect 3421 16640 3433 16643
rect 3108 16612 3433 16640
rect 3108 16600 3114 16612
rect 3421 16609 3433 16612
rect 3467 16609 3479 16643
rect 4080 16640 4108 16680
rect 8294 16668 8300 16720
rect 8352 16717 8358 16720
rect 8352 16711 8416 16717
rect 8352 16677 8370 16711
rect 8404 16677 8416 16711
rect 8352 16671 8416 16677
rect 8352 16668 8358 16671
rect 9306 16668 9312 16720
rect 9364 16708 9370 16720
rect 9677 16711 9735 16717
rect 9677 16708 9689 16711
rect 9364 16680 9689 16708
rect 9364 16668 9370 16680
rect 9677 16677 9689 16680
rect 9723 16708 9735 16711
rect 10413 16711 10471 16717
rect 10413 16708 10425 16711
rect 9723 16680 10425 16708
rect 9723 16677 9735 16680
rect 9677 16671 9735 16677
rect 10413 16677 10425 16680
rect 10459 16677 10471 16711
rect 12360 16708 12388 16748
rect 12897 16745 12909 16779
rect 12943 16776 12955 16779
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 12943 16748 14197 16776
rect 12943 16745 12955 16748
rect 12897 16739 12955 16745
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 14185 16739 14243 16745
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 15749 16779 15807 16785
rect 15749 16776 15761 16779
rect 15620 16748 15761 16776
rect 15620 16736 15626 16748
rect 15749 16745 15761 16748
rect 15795 16745 15807 16779
rect 18506 16776 18512 16788
rect 15749 16739 15807 16745
rect 15856 16748 17632 16776
rect 18467 16748 18512 16776
rect 13265 16711 13323 16717
rect 13265 16708 13277 16711
rect 12360 16680 13277 16708
rect 10413 16671 10471 16677
rect 13265 16677 13277 16680
rect 13311 16677 13323 16711
rect 13265 16671 13323 16677
rect 13357 16711 13415 16717
rect 13357 16677 13369 16711
rect 13403 16708 13415 16711
rect 13446 16708 13452 16720
rect 13403 16680 13452 16708
rect 13403 16677 13415 16680
rect 13357 16671 13415 16677
rect 13446 16668 13452 16680
rect 13504 16708 13510 16720
rect 15856 16708 15884 16748
rect 16574 16708 16580 16720
rect 13504 16680 15884 16708
rect 16535 16680 16580 16708
rect 13504 16668 13510 16680
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 3421 16603 3479 16609
rect 3528 16612 4108 16640
rect 566 16532 572 16584
rect 624 16572 630 16584
rect 3528 16581 3556 16612
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4338 16640 4344 16652
rect 4212 16612 4344 16640
rect 4212 16600 4218 16612
rect 4338 16600 4344 16612
rect 4396 16640 4402 16652
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 4396 16612 4445 16640
rect 4396 16600 4402 16612
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 5810 16640 5816 16652
rect 5307 16612 5816 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 6178 16640 6184 16652
rect 6139 16612 6184 16640
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 6454 16649 6460 16652
rect 6448 16640 6460 16649
rect 6415 16612 6460 16640
rect 6448 16603 6460 16612
rect 6454 16600 6460 16603
rect 6512 16600 6518 16652
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 7064 16612 8125 16640
rect 7064 16600 7070 16612
rect 8113 16609 8125 16612
rect 8159 16640 8171 16643
rect 9766 16640 9772 16652
rect 8159 16612 9772 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 11698 16649 11704 16652
rect 11692 16640 11704 16649
rect 11659 16612 11704 16640
rect 11692 16603 11704 16612
rect 11698 16600 11704 16603
rect 11756 16600 11762 16652
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13136 16612 14105 16640
rect 13136 16600 13142 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 14642 16600 14648 16652
rect 14700 16640 14706 16652
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14700 16612 14749 16640
rect 14700 16600 14706 16612
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 14967 16612 15669 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 16298 16640 16304 16652
rect 16259 16612 16304 16640
rect 15657 16603 15715 16609
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 17120 16643 17178 16649
rect 17120 16609 17132 16643
rect 17166 16640 17178 16643
rect 17494 16640 17500 16652
rect 17166 16612 17500 16640
rect 17166 16609 17178 16612
rect 17120 16603 17178 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 17604 16640 17632 16748
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 18877 16779 18935 16785
rect 18877 16745 18889 16779
rect 18923 16776 18935 16779
rect 19702 16776 19708 16788
rect 18923 16748 19708 16776
rect 18923 16745 18935 16748
rect 18877 16739 18935 16745
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 21082 16776 21088 16788
rect 21043 16748 21088 16776
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 21269 16779 21327 16785
rect 21269 16745 21281 16779
rect 21315 16776 21327 16779
rect 22005 16779 22063 16785
rect 22005 16776 22017 16779
rect 21315 16748 22017 16776
rect 21315 16745 21327 16748
rect 21269 16739 21327 16745
rect 22005 16745 22017 16748
rect 22051 16745 22063 16779
rect 22005 16739 22063 16745
rect 17770 16668 17776 16720
rect 17828 16708 17834 16720
rect 19150 16708 19156 16720
rect 17828 16680 19156 16708
rect 17828 16668 17834 16680
rect 19150 16668 19156 16680
rect 19208 16708 19214 16720
rect 19208 16680 19380 16708
rect 19208 16668 19214 16680
rect 18969 16643 19027 16649
rect 17604 16612 17908 16640
rect 2869 16575 2927 16581
rect 2869 16572 2881 16575
rect 624 16544 2881 16572
rect 624 16532 630 16544
rect 2869 16541 2881 16544
rect 2915 16572 2927 16575
rect 3513 16575 3571 16581
rect 3513 16572 3525 16575
rect 2915 16544 3525 16572
rect 2915 16541 2927 16544
rect 2869 16535 2927 16541
rect 3513 16541 3525 16544
rect 3559 16541 3571 16575
rect 3513 16535 3571 16541
rect 3697 16575 3755 16581
rect 3697 16541 3709 16575
rect 3743 16572 3755 16575
rect 3878 16572 3884 16584
rect 3743 16544 3884 16572
rect 3743 16541 3755 16544
rect 3697 16535 3755 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 3970 16532 3976 16584
rect 4028 16572 4034 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4028 16544 4629 16572
rect 4028 16532 4034 16544
rect 4617 16541 4629 16544
rect 4663 16572 4675 16575
rect 5445 16575 5503 16581
rect 5445 16572 5457 16575
rect 4663 16544 5457 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 5445 16541 5457 16544
rect 5491 16572 5503 16575
rect 5902 16572 5908 16584
rect 5491 16544 5908 16572
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 5902 16532 5908 16544
rect 5960 16532 5966 16584
rect 9858 16572 9864 16584
rect 9771 16544 9864 16572
rect 9858 16532 9864 16544
rect 9916 16572 9922 16584
rect 10410 16572 10416 16584
rect 9916 16544 10416 16572
rect 9916 16532 9922 16544
rect 10410 16532 10416 16544
rect 10468 16572 10474 16584
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 10468 16544 10517 16572
rect 10468 16532 10474 16544
rect 10505 16541 10517 16544
rect 10551 16541 10563 16575
rect 10505 16535 10563 16541
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16572 10655 16575
rect 11146 16572 11152 16584
rect 10643 16544 11152 16572
rect 10643 16541 10655 16544
rect 10597 16535 10655 16541
rect 2682 16464 2688 16516
rect 2740 16504 2746 16516
rect 9493 16507 9551 16513
rect 2740 16476 5672 16504
rect 2740 16464 2746 16476
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 2225 16439 2283 16445
rect 2225 16436 2237 16439
rect 1820 16408 2237 16436
rect 1820 16396 1826 16408
rect 2225 16405 2237 16408
rect 2271 16436 2283 16439
rect 3326 16436 3332 16448
rect 2271 16408 3332 16436
rect 2271 16405 2283 16408
rect 2225 16399 2283 16405
rect 3326 16396 3332 16408
rect 3384 16396 3390 16448
rect 4065 16439 4123 16445
rect 4065 16405 4077 16439
rect 4111 16436 4123 16439
rect 4338 16436 4344 16448
rect 4111 16408 4344 16436
rect 4111 16405 4123 16408
rect 4065 16399 4123 16405
rect 4338 16396 4344 16408
rect 4396 16396 4402 16448
rect 4890 16436 4896 16448
rect 4851 16408 4896 16436
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 5644 16436 5672 16476
rect 9493 16473 9505 16507
rect 9539 16504 9551 16507
rect 9950 16504 9956 16516
rect 9539 16476 9956 16504
rect 9539 16473 9551 16476
rect 9493 16467 9551 16473
rect 9950 16464 9956 16476
rect 10008 16504 10014 16516
rect 10612 16504 10640 16535
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 11425 16575 11483 16581
rect 11425 16541 11437 16575
rect 11471 16541 11483 16575
rect 13538 16572 13544 16584
rect 11425 16535 11483 16541
rect 12820 16544 13544 16572
rect 10008 16476 10640 16504
rect 10008 16464 10014 16476
rect 8754 16436 8760 16448
rect 5644 16408 8760 16436
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 11440 16436 11468 16535
rect 12710 16464 12716 16516
rect 12768 16504 12774 16516
rect 12820 16513 12848 16544
rect 13538 16532 13544 16544
rect 13596 16572 13602 16584
rect 14274 16572 14280 16584
rect 13596 16544 14044 16572
rect 14235 16544 14280 16572
rect 13596 16532 13602 16544
rect 12805 16507 12863 16513
rect 12805 16504 12817 16507
rect 12768 16476 12817 16504
rect 12768 16464 12774 16476
rect 12805 16473 12817 16476
rect 12851 16473 12863 16507
rect 13722 16504 13728 16516
rect 13683 16476 13728 16504
rect 12805 16467 12863 16473
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 14016 16504 14044 16544
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 16724 16544 16865 16572
rect 16724 16532 16730 16544
rect 16853 16541 16865 16544
rect 16899 16541 16911 16575
rect 17880 16572 17908 16612
rect 18969 16609 18981 16643
rect 19015 16640 19027 16643
rect 19242 16640 19248 16652
rect 19015 16612 19248 16640
rect 19015 16609 19027 16612
rect 18969 16603 19027 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19352 16649 19380 16680
rect 19337 16643 19395 16649
rect 19337 16609 19349 16643
rect 19383 16609 19395 16643
rect 19337 16603 19395 16609
rect 19604 16643 19662 16649
rect 19604 16609 19616 16643
rect 19650 16640 19662 16643
rect 20346 16640 20352 16652
rect 19650 16612 20352 16640
rect 19650 16609 19662 16612
rect 19604 16603 19662 16609
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 20898 16640 20904 16652
rect 20859 16612 20904 16640
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 19058 16572 19064 16584
rect 17880 16544 19064 16572
rect 16853 16535 16911 16541
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 19153 16575 19211 16581
rect 19153 16541 19165 16575
rect 19199 16572 19211 16575
rect 19199 16544 19288 16572
rect 19199 16541 19211 16544
rect 19153 16535 19211 16541
rect 15856 16504 15884 16532
rect 14016 16476 15884 16504
rect 11790 16436 11796 16448
rect 11440 16408 11796 16436
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 13262 16396 13268 16448
rect 13320 16436 13326 16448
rect 13814 16436 13820 16448
rect 13320 16408 13820 16436
rect 13320 16396 13326 16408
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 13906 16396 13912 16448
rect 13964 16436 13970 16448
rect 14553 16439 14611 16445
rect 14553 16436 14565 16439
rect 13964 16408 14565 16436
rect 13964 16396 13970 16408
rect 14553 16405 14565 16408
rect 14599 16436 14611 16439
rect 14734 16436 14740 16448
rect 14599 16408 14740 16436
rect 14599 16405 14611 16408
rect 14553 16399 14611 16405
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 15289 16439 15347 16445
rect 15289 16436 15301 16439
rect 15252 16408 15301 16436
rect 15252 16396 15258 16408
rect 15289 16405 15301 16408
rect 15335 16405 15347 16439
rect 15289 16399 15347 16405
rect 18046 16396 18052 16448
rect 18104 16436 18110 16448
rect 18233 16439 18291 16445
rect 18233 16436 18245 16439
rect 18104 16408 18245 16436
rect 18104 16396 18110 16408
rect 18233 16405 18245 16408
rect 18279 16405 18291 16439
rect 19260 16436 19288 16544
rect 19334 16436 19340 16448
rect 19247 16408 19340 16436
rect 18233 16399 18291 16405
rect 19334 16396 19340 16408
rect 19392 16436 19398 16448
rect 20717 16439 20775 16445
rect 20717 16436 20729 16439
rect 19392 16408 20729 16436
rect 19392 16396 19398 16408
rect 20717 16405 20729 16408
rect 20763 16405 20775 16439
rect 20717 16399 20775 16405
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2317 16235 2375 16241
rect 2317 16201 2329 16235
rect 2363 16232 2375 16235
rect 2866 16232 2872 16244
rect 2363 16204 2872 16232
rect 2363 16201 2375 16204
rect 2317 16195 2375 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3970 16232 3976 16244
rect 3931 16204 3976 16232
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4246 16232 4252 16244
rect 4207 16204 4252 16232
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 5077 16235 5135 16241
rect 5077 16201 5089 16235
rect 5123 16232 5135 16235
rect 5534 16232 5540 16244
rect 5123 16204 5540 16232
rect 5123 16201 5135 16204
rect 5077 16195 5135 16201
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 6825 16235 6883 16241
rect 6825 16201 6837 16235
rect 6871 16232 6883 16235
rect 7098 16232 7104 16244
rect 6871 16204 7104 16232
rect 6871 16201 6883 16204
rect 6825 16195 6883 16201
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 11238 16232 11244 16244
rect 9355 16204 11244 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 11517 16235 11575 16241
rect 11517 16201 11529 16235
rect 11563 16232 11575 16235
rect 11698 16232 11704 16244
rect 11563 16204 11704 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 12124 16204 12173 16232
rect 12124 16192 12130 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 12161 16195 12219 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16684 16204 16773 16232
rect 4154 16164 4160 16176
rect 4115 16136 4160 16164
rect 4154 16124 4160 16136
rect 4212 16124 4218 16176
rect 9858 16164 9864 16176
rect 4264 16136 9864 16164
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 2314 16028 2320 16040
rect 2179 16000 2320 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2593 16031 2651 16037
rect 2593 15997 2605 16031
rect 2639 16028 2651 16031
rect 3142 16028 3148 16040
rect 2639 16000 3148 16028
rect 2639 15997 2651 16000
rect 2593 15991 2651 15997
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3786 16028 3792 16040
rect 3384 16000 3792 16028
rect 3384 15988 3390 16000
rect 3786 15988 3792 16000
rect 3844 16028 3850 16040
rect 4264 16028 4292 16136
rect 9858 16124 9864 16136
rect 9916 16124 9922 16176
rect 4338 16056 4344 16108
rect 4396 16096 4402 16108
rect 4709 16099 4767 16105
rect 4709 16096 4721 16099
rect 4396 16068 4721 16096
rect 4396 16056 4402 16068
rect 4709 16065 4721 16068
rect 4755 16065 4767 16099
rect 4709 16059 4767 16065
rect 4798 16056 4804 16108
rect 4856 16096 4862 16108
rect 5629 16099 5687 16105
rect 5629 16096 5641 16099
rect 4856 16068 5641 16096
rect 4856 16056 4862 16068
rect 5629 16065 5641 16068
rect 5675 16065 5687 16099
rect 5629 16059 5687 16065
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 7558 16096 7564 16108
rect 7515 16068 7564 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 8478 16096 8484 16108
rect 8343 16068 8484 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16096 10011 16099
rect 15304 16096 15332 16192
rect 9999 16068 10272 16096
rect 15304 16068 15516 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 3844 16000 4292 16028
rect 4617 16031 4675 16037
rect 3844 15988 3850 16000
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 4890 16028 4896 16040
rect 4663 16000 4896 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 7374 15988 7380 16040
rect 7432 16028 7438 16040
rect 8757 16031 8815 16037
rect 8757 16028 8769 16031
rect 7432 16000 8769 16028
rect 7432 15988 7438 16000
rect 8757 15997 8769 16000
rect 8803 15997 8815 16031
rect 9674 16028 9680 16040
rect 9635 16000 9680 16028
rect 8757 15991 8815 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 16028 9827 16031
rect 10042 16028 10048 16040
rect 9815 16000 10048 16028
rect 9815 15997 9827 16000
rect 9769 15991 9827 15997
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 2860 15963 2918 15969
rect 2860 15929 2872 15963
rect 2906 15960 2918 15963
rect 3878 15960 3884 15972
rect 2906 15932 3884 15960
rect 2906 15929 2918 15932
rect 2860 15923 2918 15929
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 4982 15920 4988 15972
rect 5040 15960 5046 15972
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 5040 15932 5549 15960
rect 5040 15920 5046 15932
rect 5537 15929 5549 15932
rect 5583 15929 5595 15963
rect 5537 15923 5595 15929
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 8021 15963 8079 15969
rect 7239 15932 7696 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5445 15895 5503 15901
rect 5445 15892 5457 15895
rect 5224 15864 5457 15892
rect 5224 15852 5230 15864
rect 5445 15861 5457 15864
rect 5491 15861 5503 15895
rect 5445 15855 5503 15861
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7558 15892 7564 15904
rect 7331 15864 7564 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7558 15852 7564 15864
rect 7616 15852 7622 15904
rect 7668 15901 7696 15932
rect 8021 15929 8033 15963
rect 8067 15960 8079 15963
rect 8846 15960 8852 15972
rect 8067 15932 8852 15960
rect 8067 15929 8079 15932
rect 8021 15923 8079 15929
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 10152 15960 10180 15991
rect 9692 15932 10180 15960
rect 10244 15960 10272 16068
rect 11790 15988 11796 16040
rect 11848 16028 11854 16040
rect 12066 16028 12072 16040
rect 11848 16000 12072 16028
rect 11848 15988 11854 16000
rect 12066 15988 12072 16000
rect 12124 16028 12130 16040
rect 12710 16037 12716 16040
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 12124 16000 12449 16028
rect 12124 15988 12130 16000
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12704 16028 12716 16037
rect 12671 16000 12716 16028
rect 12437 15991 12495 15997
rect 12704 15991 12716 16000
rect 10410 15969 10416 15972
rect 10404 15960 10416 15969
rect 10244 15932 10416 15960
rect 9692 15904 9720 15932
rect 10404 15923 10416 15932
rect 10410 15920 10416 15923
rect 10468 15920 10474 15972
rect 12452 15960 12480 15991
rect 12710 15988 12716 15991
rect 12768 15988 12774 16040
rect 13906 16028 13912 16040
rect 12811 16000 13912 16028
rect 12811 15960 12839 16000
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 15381 16031 15439 16037
rect 15381 15997 15393 16031
rect 15427 15997 15439 16031
rect 15488 16028 15516 16068
rect 16390 16056 16396 16108
rect 16448 16096 16454 16108
rect 16684 16096 16712 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 16761 16195 16819 16201
rect 18325 16235 18383 16241
rect 18325 16201 18337 16235
rect 18371 16232 18383 16235
rect 18690 16232 18696 16244
rect 18371 16204 18696 16232
rect 18371 16201 18383 16204
rect 18325 16195 18383 16201
rect 16853 16167 16911 16173
rect 16853 16133 16865 16167
rect 16899 16164 16911 16167
rect 17218 16164 17224 16176
rect 16899 16136 17224 16164
rect 16899 16133 16911 16136
rect 16853 16127 16911 16133
rect 17218 16124 17224 16136
rect 17276 16124 17282 16176
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 16448 16068 17417 16096
rect 16448 16056 16454 16068
rect 17405 16065 17417 16068
rect 17451 16065 17463 16099
rect 18340 16096 18368 16195
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 20257 16235 20315 16241
rect 20257 16232 20269 16235
rect 19484 16204 20269 16232
rect 19484 16192 19490 16204
rect 20257 16201 20269 16204
rect 20303 16201 20315 16235
rect 21266 16232 21272 16244
rect 21227 16204 21272 16232
rect 20257 16195 20315 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 20165 16167 20223 16173
rect 20165 16133 20177 16167
rect 20211 16164 20223 16167
rect 20346 16164 20352 16176
rect 20211 16136 20352 16164
rect 20211 16133 20223 16136
rect 20165 16127 20223 16133
rect 20346 16124 20352 16136
rect 20404 16124 20410 16176
rect 17405 16059 17463 16065
rect 17512 16068 18368 16096
rect 20364 16096 20392 16124
rect 20809 16099 20867 16105
rect 20809 16096 20821 16099
rect 20364 16068 20821 16096
rect 15637 16031 15695 16037
rect 15637 16028 15649 16031
rect 15488 16000 15649 16028
rect 15381 15991 15439 15997
rect 15637 15997 15649 16000
rect 15683 15997 15695 16031
rect 17310 16028 17316 16040
rect 17223 16000 17316 16028
rect 15637 15991 15695 15997
rect 14176 15963 14234 15969
rect 14176 15960 14188 15963
rect 10520 15932 11744 15960
rect 12452 15932 12839 15960
rect 13832 15932 14188 15960
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15861 7711 15895
rect 7653 15855 7711 15861
rect 8113 15895 8171 15901
rect 8113 15861 8125 15895
rect 8159 15892 8171 15895
rect 8202 15892 8208 15904
rect 8159 15864 8208 15892
rect 8159 15861 8171 15864
rect 8113 15855 8171 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8573 15895 8631 15901
rect 8573 15861 8585 15895
rect 8619 15892 8631 15895
rect 9674 15892 9680 15904
rect 8619 15864 9680 15892
rect 8619 15861 8631 15864
rect 8573 15855 8631 15861
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10520 15892 10548 15932
rect 11606 15892 11612 15904
rect 9916 15864 10548 15892
rect 11567 15864 11612 15892
rect 9916 15852 9922 15864
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 11716 15892 11744 15932
rect 13722 15892 13728 15904
rect 11716 15864 13728 15892
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 13832 15901 13860 15932
rect 14176 15929 14188 15932
rect 14222 15960 14234 15963
rect 14274 15960 14280 15972
rect 14222 15932 14280 15960
rect 14222 15929 14234 15932
rect 14176 15923 14234 15929
rect 14274 15920 14280 15932
rect 14332 15960 14338 15972
rect 14734 15960 14740 15972
rect 14332 15932 14740 15960
rect 14332 15920 14338 15932
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 15396 15960 15424 15991
rect 17310 15988 17316 16000
rect 17368 16028 17374 16040
rect 17512 16028 17540 16068
rect 20809 16065 20821 16068
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 17368 16000 17540 16028
rect 17368 15988 17374 16000
rect 17770 15988 17776 16040
rect 17828 16028 17834 16040
rect 18785 16031 18843 16037
rect 18785 16028 18797 16031
rect 17828 16000 18797 16028
rect 17828 15988 17834 16000
rect 18785 15997 18797 16000
rect 18831 15997 18843 16031
rect 18785 15991 18843 15997
rect 19518 15988 19524 16040
rect 19576 16028 19582 16040
rect 19978 16028 19984 16040
rect 19576 16000 19984 16028
rect 19576 15988 19582 16000
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 21085 16031 21143 16037
rect 21085 15997 21097 16031
rect 21131 16028 21143 16031
rect 21131 16000 21312 16028
rect 21131 15997 21143 16000
rect 21085 15991 21143 15997
rect 16666 15960 16672 15972
rect 15396 15932 16672 15960
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 18049 15963 18107 15969
rect 18049 15960 18061 15963
rect 17236 15932 18061 15960
rect 13817 15895 13875 15901
rect 13817 15861 13829 15895
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 14090 15852 14096 15904
rect 14148 15892 14154 15904
rect 17236 15901 17264 15932
rect 18049 15929 18061 15932
rect 18095 15960 18107 15963
rect 18874 15960 18880 15972
rect 18095 15932 18880 15960
rect 18095 15929 18107 15932
rect 18049 15923 18107 15929
rect 18874 15920 18880 15932
rect 18932 15920 18938 15972
rect 19052 15963 19110 15969
rect 19052 15929 19064 15963
rect 19098 15960 19110 15963
rect 19150 15960 19156 15972
rect 19098 15932 19156 15960
rect 19098 15929 19110 15932
rect 19052 15923 19110 15929
rect 19150 15920 19156 15932
rect 19208 15920 19214 15972
rect 19242 15920 19248 15972
rect 19300 15960 19306 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 19300 15932 20729 15960
rect 19300 15920 19306 15932
rect 20717 15929 20729 15932
rect 20763 15929 20775 15963
rect 20717 15923 20775 15929
rect 21284 15904 21312 16000
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 14148 15864 17233 15892
rect 14148 15852 14154 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 17681 15895 17739 15901
rect 17681 15861 17693 15895
rect 17727 15892 17739 15895
rect 17954 15892 17960 15904
rect 17727 15864 17960 15892
rect 17727 15861 17739 15864
rect 17681 15855 17739 15861
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 20530 15852 20536 15904
rect 20588 15892 20594 15904
rect 20625 15895 20683 15901
rect 20625 15892 20637 15895
rect 20588 15864 20637 15892
rect 20588 15852 20594 15864
rect 20625 15861 20637 15864
rect 20671 15861 20683 15895
rect 20625 15855 20683 15861
rect 21266 15852 21272 15904
rect 21324 15892 21330 15904
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 21324 15864 21465 15892
rect 21324 15852 21330 15864
rect 21453 15861 21465 15864
rect 21499 15861 21511 15895
rect 21453 15855 21511 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2317 15691 2375 15697
rect 2317 15657 2329 15691
rect 2363 15688 2375 15691
rect 2774 15688 2780 15700
rect 2363 15660 2780 15688
rect 2363 15657 2375 15660
rect 2317 15651 2375 15657
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5997 15691 6055 15697
rect 5997 15657 6009 15691
rect 6043 15688 6055 15691
rect 6178 15688 6184 15700
rect 6043 15660 6184 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7616 15660 7941 15688
rect 7616 15648 7622 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 7929 15651 7987 15657
rect 8036 15660 8309 15688
rect 2593 15623 2651 15629
rect 2593 15620 2605 15623
rect 1780 15592 2605 15620
rect 1780 15561 1808 15592
rect 2593 15589 2605 15592
rect 2639 15620 2651 15623
rect 4065 15623 4123 15629
rect 2639 15592 4016 15620
rect 2639 15589 2651 15592
rect 2593 15583 2651 15589
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 2685 15555 2743 15561
rect 2685 15552 2697 15555
rect 2179 15524 2697 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 2685 15521 2697 15524
rect 2731 15521 2743 15555
rect 2685 15515 2743 15521
rect 2700 15484 2728 15515
rect 3988 15484 4016 15592
rect 4065 15589 4077 15623
rect 4111 15620 4123 15623
rect 5537 15623 5595 15629
rect 5537 15620 5549 15623
rect 4111 15592 5549 15620
rect 4111 15589 4123 15592
rect 4065 15583 4123 15589
rect 5537 15589 5549 15592
rect 5583 15589 5595 15623
rect 8036 15620 8064 15660
rect 8297 15657 8309 15660
rect 8343 15688 8355 15691
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 8343 15660 9229 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 9217 15657 9229 15660
rect 9263 15688 9275 15691
rect 9398 15688 9404 15700
rect 9263 15660 9404 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 10870 15688 10876 15700
rect 9539 15660 10876 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11149 15691 11207 15697
rect 11149 15657 11161 15691
rect 11195 15688 11207 15691
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11195 15660 12357 15688
rect 11195 15657 11207 15660
rect 11149 15651 11207 15657
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 14185 15691 14243 15697
rect 14185 15657 14197 15691
rect 14231 15688 14243 15691
rect 14458 15688 14464 15700
rect 14231 15660 14464 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14645 15691 14703 15697
rect 14645 15657 14657 15691
rect 14691 15688 14703 15691
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 14691 15660 15301 15688
rect 14691 15657 14703 15660
rect 14645 15651 14703 15657
rect 15289 15657 15301 15660
rect 15335 15657 15347 15691
rect 15289 15651 15347 15657
rect 15930 15648 15936 15700
rect 15988 15688 15994 15700
rect 17494 15688 17500 15700
rect 15988 15660 17356 15688
rect 17455 15660 17500 15688
rect 15988 15648 15994 15660
rect 5537 15583 5595 15589
rect 6104 15592 8064 15620
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 4304 15524 4721 15552
rect 4304 15512 4310 15524
rect 4709 15521 4721 15524
rect 4755 15521 4767 15555
rect 4709 15515 4767 15521
rect 5350 15512 5356 15564
rect 5408 15552 5414 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5408 15524 5641 15552
rect 5408 15512 5414 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 4798 15484 4804 15496
rect 2700 15456 3924 15484
rect 3988 15456 4660 15484
rect 4759 15456 4804 15484
rect 3896 15416 3924 15456
rect 4632 15416 4660 15456
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15484 5043 15487
rect 5534 15484 5540 15496
rect 5031 15456 5540 15484
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 5902 15484 5908 15496
rect 5859 15456 5908 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 6104 15416 6132 15592
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 11517 15623 11575 15629
rect 8260 15592 10088 15620
rect 8260 15580 8266 15592
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 7374 15552 7380 15564
rect 6227 15524 7380 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 7374 15512 7380 15524
rect 7432 15512 7438 15564
rect 7558 15552 7564 15564
rect 7519 15524 7564 15552
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 9950 15561 9956 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 7668 15524 9505 15552
rect 6270 15444 6276 15496
rect 6328 15484 6334 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6328 15456 6837 15484
rect 6328 15444 6334 15456
rect 6825 15453 6837 15456
rect 6871 15484 6883 15487
rect 7668 15484 7696 15524
rect 9493 15521 9505 15524
rect 9539 15521 9551 15555
rect 9944 15552 9956 15561
rect 9911 15524 9956 15552
rect 9493 15515 9551 15521
rect 9944 15515 9956 15524
rect 9950 15512 9956 15515
rect 10008 15512 10014 15564
rect 10060 15552 10088 15592
rect 11517 15589 11529 15623
rect 11563 15620 11575 15623
rect 11698 15620 11704 15632
rect 11563 15592 11704 15620
rect 11563 15589 11575 15592
rect 11517 15583 11575 15589
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 12437 15623 12495 15629
rect 12437 15620 12449 15623
rect 11848 15592 12449 15620
rect 11848 15580 11854 15592
rect 12437 15589 12449 15592
rect 12483 15589 12495 15623
rect 12437 15583 12495 15589
rect 14553 15623 14611 15629
rect 14553 15589 14565 15623
rect 14599 15620 14611 15623
rect 15194 15620 15200 15632
rect 14599 15592 15200 15620
rect 14599 15589 14611 15592
rect 14553 15583 14611 15589
rect 15194 15580 15200 15592
rect 15252 15580 15258 15632
rect 15746 15620 15752 15632
rect 15304 15592 15752 15620
rect 10060 15524 13676 15552
rect 6871 15456 7696 15484
rect 8389 15487 8447 15493
rect 6871 15453 6883 15456
rect 6825 15447 6883 15453
rect 8389 15453 8401 15487
rect 8435 15453 8447 15487
rect 8389 15447 8447 15453
rect 7374 15416 7380 15428
rect 3896 15388 4568 15416
rect 4632 15388 6132 15416
rect 7335 15388 7380 15416
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 4341 15351 4399 15357
rect 4341 15348 4353 15351
rect 2188 15320 4353 15348
rect 2188 15308 2194 15320
rect 4341 15317 4353 15320
rect 4387 15317 4399 15351
rect 4540 15348 4568 15388
rect 7374 15376 7380 15388
rect 7432 15376 7438 15428
rect 7745 15419 7803 15425
rect 7745 15385 7757 15419
rect 7791 15416 7803 15419
rect 8202 15416 8208 15428
rect 7791 15388 8208 15416
rect 7791 15385 7803 15388
rect 7745 15379 7803 15385
rect 8202 15376 8208 15388
rect 8260 15376 8266 15428
rect 8404 15416 8432 15447
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 8757 15487 8815 15493
rect 8536 15456 8581 15484
rect 8536 15444 8542 15456
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 8846 15484 8852 15496
rect 8803 15456 8852 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11606 15484 11612 15496
rect 11296 15456 11612 15484
rect 11296 15444 11302 15456
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15453 11759 15487
rect 11701 15447 11759 15453
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 8404 15388 9076 15416
rect 9048 15360 9076 15388
rect 11146 15376 11152 15428
rect 11204 15416 11210 15428
rect 11716 15416 11744 15447
rect 11204 15388 11744 15416
rect 11204 15376 11210 15388
rect 11882 15376 11888 15428
rect 11940 15416 11946 15428
rect 11977 15419 12035 15425
rect 11977 15416 11989 15419
rect 11940 15388 11989 15416
rect 11940 15376 11946 15388
rect 11977 15385 11989 15388
rect 12023 15385 12035 15419
rect 11977 15379 12035 15385
rect 6730 15348 6736 15360
rect 4540 15320 6736 15348
rect 4341 15311 4399 15317
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 7006 15348 7012 15360
rect 6967 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 9030 15348 9036 15360
rect 8991 15320 9036 15348
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 9858 15308 9864 15360
rect 9916 15348 9922 15360
rect 10318 15348 10324 15360
rect 9916 15320 10324 15348
rect 9916 15308 9922 15320
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 10410 15308 10416 15360
rect 10468 15348 10474 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 10468 15320 11069 15348
rect 10468 15308 10474 15320
rect 11057 15317 11069 15320
rect 11103 15348 11115 15351
rect 12544 15348 12572 15447
rect 13648 15416 13676 15524
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 15304 15552 15332 15592
rect 15746 15580 15752 15592
rect 15804 15580 15810 15632
rect 16390 15629 16396 15632
rect 16384 15620 16396 15629
rect 16351 15592 16396 15620
rect 16384 15583 16396 15592
rect 16390 15580 16396 15583
rect 16448 15580 16454 15632
rect 17328 15620 17356 15660
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 19150 15688 19156 15700
rect 19111 15660 19156 15688
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 19242 15648 19248 15700
rect 19300 15688 19306 15700
rect 20622 15688 20628 15700
rect 19300 15660 19345 15688
rect 20583 15660 20628 15688
rect 19300 15648 19306 15660
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 21082 15688 21088 15700
rect 21043 15660 21088 15688
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 21450 15688 21456 15700
rect 21411 15660 21456 15688
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 18046 15629 18052 15632
rect 18040 15620 18052 15629
rect 17328 15592 17816 15620
rect 18007 15592 18052 15620
rect 13780 15524 15332 15552
rect 15657 15555 15715 15561
rect 13780 15512 13786 15524
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 17678 15552 17684 15564
rect 15703 15524 17684 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 17788 15552 17816 15592
rect 18040 15583 18052 15592
rect 18046 15580 18052 15583
rect 18104 15580 18110 15632
rect 19168 15620 19196 15648
rect 19168 15592 19840 15620
rect 17788 15524 18828 15552
rect 14734 15484 14740 15496
rect 14695 15456 14740 15484
rect 14734 15444 14740 15456
rect 14792 15444 14798 15496
rect 15838 15484 15844 15496
rect 15799 15456 15844 15484
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15453 16175 15487
rect 17770 15484 17776 15496
rect 16117 15447 16175 15453
rect 17420 15456 17776 15484
rect 15930 15416 15936 15428
rect 13648 15388 15936 15416
rect 15930 15376 15936 15388
rect 15988 15376 15994 15428
rect 12894 15348 12900 15360
rect 11103 15320 12572 15348
rect 12855 15320 12900 15348
rect 11103 15317 11115 15320
rect 11057 15311 11115 15317
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 16132 15348 16160 15447
rect 16758 15348 16764 15360
rect 16132 15320 16764 15348
rect 16758 15308 16764 15320
rect 16816 15348 16822 15360
rect 17420 15348 17448 15456
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 17678 15348 17684 15360
rect 16816 15320 17448 15348
rect 17639 15320 17684 15348
rect 16816 15308 16822 15320
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18690 15348 18696 15360
rect 18012 15320 18696 15348
rect 18012 15308 18018 15320
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 18800 15348 18828 15524
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 19392 15524 19625 15552
rect 19392 15512 19398 15524
rect 19613 15521 19625 15524
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 19058 15444 19064 15496
rect 19116 15484 19122 15496
rect 19812 15493 19840 15592
rect 20438 15552 20444 15564
rect 20399 15524 20444 15552
rect 20438 15512 20444 15524
rect 20496 15512 20502 15564
rect 20898 15552 20904 15564
rect 20859 15524 20904 15552
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15521 21327 15555
rect 21269 15515 21327 15521
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19116 15456 19717 15484
rect 19116 15444 19122 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15453 19855 15487
rect 21284 15484 21312 15515
rect 19797 15447 19855 15453
rect 20272 15456 21312 15484
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 20073 15419 20131 15425
rect 20073 15416 20085 15419
rect 19392 15388 20085 15416
rect 19392 15376 19398 15388
rect 20073 15385 20085 15388
rect 20119 15385 20131 15419
rect 20073 15379 20131 15385
rect 20272 15357 20300 15456
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 18800 15320 20269 15348
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1946 15144 1952 15156
rect 1907 15116 1952 15144
rect 1946 15104 1952 15116
rect 2004 15104 2010 15156
rect 3053 15147 3111 15153
rect 3053 15113 3065 15147
rect 3099 15144 3111 15147
rect 4982 15144 4988 15156
rect 3099 15116 4988 15144
rect 3099 15113 3111 15116
rect 3053 15107 3111 15113
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 5592 15116 5641 15144
rect 5592 15104 5598 15116
rect 5629 15113 5641 15116
rect 5675 15113 5687 15147
rect 5629 15107 5687 15113
rect 6362 15104 6368 15156
rect 6420 15144 6426 15156
rect 7653 15147 7711 15153
rect 7653 15144 7665 15147
rect 6420 15116 7665 15144
rect 6420 15104 6426 15116
rect 7653 15113 7665 15116
rect 7699 15113 7711 15147
rect 7653 15107 7711 15113
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8260 15116 8677 15144
rect 8260 15104 8266 15116
rect 8665 15113 8677 15116
rect 8711 15144 8723 15147
rect 9217 15147 9275 15153
rect 9217 15144 9229 15147
rect 8711 15116 9229 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 9217 15113 9229 15116
rect 9263 15113 9275 15147
rect 9217 15107 9275 15113
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 9490 15144 9496 15156
rect 9447 15116 9496 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 11790 15144 11796 15156
rect 10919 15116 11796 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12253 15147 12311 15153
rect 12253 15144 12265 15147
rect 11940 15116 12265 15144
rect 11940 15104 11946 15116
rect 12253 15113 12265 15116
rect 12299 15144 12311 15147
rect 15746 15144 15752 15156
rect 12299 15116 14780 15144
rect 15707 15116 15752 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 4062 15076 4068 15088
rect 3200 15048 4068 15076
rect 3200 15036 3206 15048
rect 4062 15036 4068 15048
rect 4120 15076 4126 15088
rect 4120 15048 4292 15076
rect 4120 15036 4126 15048
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 15008 3755 15011
rect 3970 15008 3976 15020
rect 3743 14980 3976 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4264 15017 4292 15048
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 8938 15076 8944 15088
rect 7524 15048 8944 15076
rect 7524 15036 7530 15048
rect 8938 15036 8944 15048
rect 8996 15076 9002 15088
rect 9585 15079 9643 15085
rect 9585 15076 9597 15079
rect 8996 15048 9597 15076
rect 8996 15036 9002 15048
rect 9585 15045 9597 15048
rect 9631 15076 9643 15079
rect 10042 15076 10048 15088
rect 9631 15048 10048 15076
rect 9631 15045 9643 15048
rect 9585 15039 9643 15045
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 12437 15079 12495 15085
rect 10244 15048 12020 15076
rect 10244 15020 10272 15048
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 5316 14980 6561 15008
rect 5316 14968 5322 14980
rect 6549 14977 6561 14980
rect 6595 15008 6607 15011
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 6595 14980 7389 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7926 15008 7932 15020
rect 7377 14971 7435 14977
rect 7760 14980 7932 15008
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14909 1823 14943
rect 2130 14940 2136 14952
rect 2091 14912 2136 14940
rect 1765 14903 1823 14909
rect 1780 14872 1808 14903
rect 2130 14900 2136 14912
rect 2188 14900 2194 14952
rect 4516 14943 4574 14949
rect 4516 14909 4528 14943
rect 4562 14940 4574 14943
rect 5718 14940 5724 14952
rect 4562 14912 5724 14940
rect 4562 14909 4574 14912
rect 4516 14903 4574 14909
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 6270 14940 6276 14952
rect 6231 14912 6276 14940
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 7760 14940 7788 14980
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 8478 15008 8484 15020
rect 8343 14980 8484 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 15008 8631 15011
rect 10226 15008 10232 15020
rect 8619 14980 10232 15008
rect 8619 14977 8631 14980
rect 8573 14971 8631 14977
rect 8588 14940 8616 14971
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11425 15011 11483 15017
rect 11425 15008 11437 15011
rect 11204 14980 11437 15008
rect 11204 14968 11210 14980
rect 11425 14977 11437 14980
rect 11471 14977 11483 15011
rect 11698 15008 11704 15020
rect 11659 14980 11704 15008
rect 11425 14971 11483 14977
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 6512 14912 7788 14940
rect 7852 14912 8616 14940
rect 9217 14943 9275 14949
rect 6512 14900 6518 14912
rect 2961 14875 3019 14881
rect 1780 14844 2820 14872
rect 2792 14813 2820 14844
rect 2961 14841 2973 14875
rect 3007 14872 3019 14875
rect 3142 14872 3148 14884
rect 3007 14844 3148 14872
rect 3007 14841 3019 14844
rect 2961 14835 3019 14841
rect 3142 14832 3148 14844
rect 3200 14872 3206 14884
rect 3421 14875 3479 14881
rect 3421 14872 3433 14875
rect 3200 14844 3433 14872
rect 3200 14832 3206 14844
rect 3421 14841 3433 14844
rect 3467 14841 3479 14875
rect 3421 14835 3479 14841
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 5813 14875 5871 14881
rect 5813 14872 5825 14875
rect 5408 14844 5825 14872
rect 5408 14832 5414 14844
rect 5813 14841 5825 14844
rect 5859 14872 5871 14875
rect 6365 14875 6423 14881
rect 5859 14844 6316 14872
rect 5859 14841 5871 14844
rect 5813 14835 5871 14841
rect 2777 14807 2835 14813
rect 2777 14773 2789 14807
rect 2823 14804 2835 14807
rect 3513 14807 3571 14813
rect 3513 14804 3525 14807
rect 2823 14776 3525 14804
rect 2823 14773 2835 14776
rect 2777 14767 2835 14773
rect 3513 14773 3525 14776
rect 3559 14804 3571 14807
rect 3970 14804 3976 14816
rect 3559 14776 3976 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 5902 14804 5908 14816
rect 5863 14776 5908 14804
rect 5902 14764 5908 14776
rect 5960 14764 5966 14816
rect 6288 14804 6316 14844
rect 6365 14841 6377 14875
rect 6411 14872 6423 14875
rect 7006 14872 7012 14884
rect 6411 14844 7012 14872
rect 6411 14841 6423 14844
rect 6365 14835 6423 14841
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 7852 14872 7880 14912
rect 9217 14909 9229 14943
rect 9263 14940 9275 14943
rect 10962 14940 10968 14952
rect 9263 14912 10968 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 11882 14940 11888 14952
rect 11287 14912 11888 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 11992 14940 12020 15048
rect 12437 15045 12449 15079
rect 12483 15076 12495 15079
rect 14752 15076 14780 15116
rect 15746 15104 15752 15116
rect 15804 15144 15810 15156
rect 16114 15144 16120 15156
rect 15804 15116 16120 15144
rect 15804 15104 15810 15116
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 16209 15147 16267 15153
rect 16209 15113 16221 15147
rect 16255 15144 16267 15147
rect 16298 15144 16304 15156
rect 16255 15116 16304 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 17865 15147 17923 15153
rect 17865 15113 17877 15147
rect 17911 15144 17923 15147
rect 17911 15116 19012 15144
rect 17911 15113 17923 15116
rect 17865 15107 17923 15113
rect 15838 15076 15844 15088
rect 12483 15048 13860 15076
rect 14752 15048 15844 15076
rect 12483 15045 12495 15048
rect 12437 15039 12495 15045
rect 12250 14968 12256 15020
rect 12308 15008 12314 15020
rect 12894 15008 12900 15020
rect 12308 14980 12900 15008
rect 12308 14968 12314 14980
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 15008 13139 15011
rect 13538 15008 13544 15020
rect 13127 14980 13544 15008
rect 13127 14977 13139 14980
rect 13081 14971 13139 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 13832 15008 13860 15048
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 17954 15076 17960 15088
rect 17144 15048 17960 15076
rect 16853 15011 16911 15017
rect 13832 14980 13952 15008
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 11992 14912 12817 14940
rect 12805 14909 12817 14912
rect 12851 14940 12863 14943
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 12851 14912 13277 14940
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 13688 14912 13737 14940
rect 13688 14900 13694 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 13924 14940 13952 14980
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 17144 15008 17172 15048
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 16899 14980 17172 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 17276 14980 17509 15008
rect 17276 14968 17282 14980
rect 17497 14977 17509 14980
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17586 14968 17592 15020
rect 17644 15008 17650 15020
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 17644 14980 18613 15008
rect 17644 14968 17650 14980
rect 18601 14977 18613 14980
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 16117 14943 16175 14949
rect 16117 14940 16129 14943
rect 13924 14912 14228 14940
rect 13817 14903 13875 14909
rect 7239 14844 7880 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7926 14832 7932 14884
rect 7984 14872 7990 14884
rect 12342 14872 12348 14884
rect 7984 14844 12348 14872
rect 7984 14832 7990 14844
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 13832 14872 13860 14903
rect 14200 14884 14228 14912
rect 14844 14912 16129 14940
rect 14090 14881 14096 14884
rect 14084 14872 14096 14881
rect 13464 14844 13860 14872
rect 14051 14844 14096 14872
rect 6454 14804 6460 14816
rect 6288 14776 6460 14804
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7800 14776 8033 14804
rect 7800 14764 7806 14776
rect 8021 14773 8033 14776
rect 8067 14773 8079 14807
rect 8021 14767 8079 14773
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 8386 14804 8392 14816
rect 8159 14776 8392 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11882 14804 11888 14816
rect 11379 14776 11888 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11882 14764 11888 14776
rect 11940 14804 11946 14816
rect 11977 14807 12035 14813
rect 11977 14804 11989 14807
rect 11940 14776 11989 14804
rect 11940 14764 11946 14776
rect 11977 14773 11989 14776
rect 12023 14773 12035 14807
rect 11977 14767 12035 14773
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 13464 14804 13492 14844
rect 14084 14835 14096 14844
rect 14090 14832 14096 14835
rect 14148 14832 14154 14884
rect 14182 14832 14188 14884
rect 14240 14832 14246 14884
rect 12124 14776 13492 14804
rect 13541 14807 13599 14813
rect 12124 14764 12130 14776
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 14642 14804 14648 14816
rect 13587 14776 14648 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 14642 14764 14648 14776
rect 14700 14804 14706 14816
rect 14844 14804 14872 14912
rect 16117 14909 16129 14912
rect 16163 14909 16175 14943
rect 16666 14940 16672 14952
rect 16117 14903 16175 14909
rect 16500 14912 16672 14940
rect 16500 14872 16528 14912
rect 16666 14900 16672 14912
rect 16724 14900 16730 14952
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14940 17463 14943
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17451 14912 17877 14940
rect 17451 14909 17463 14912
rect 17405 14903 17463 14909
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 18417 14943 18475 14949
rect 18417 14909 18429 14943
rect 18463 14940 18475 14943
rect 18690 14940 18696 14952
rect 18463 14912 18696 14940
rect 18463 14909 18475 14912
rect 18417 14903 18475 14909
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 18984 14949 19012 15116
rect 19058 15104 19064 15156
rect 19116 15144 19122 15156
rect 21358 15144 21364 15156
rect 19116 15116 19161 15144
rect 21319 15116 21364 15144
rect 19116 15104 19122 15116
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 15008 20407 15011
rect 20438 15008 20444 15020
rect 20395 14980 20444 15008
rect 20395 14977 20407 14980
rect 20349 14971 20407 14977
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 20898 15008 20904 15020
rect 20859 14980 20904 15008
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14940 19027 14943
rect 19058 14940 19064 14952
rect 19015 14912 19064 14940
rect 19015 14909 19027 14912
rect 18969 14903 19027 14909
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 19150 14900 19156 14952
rect 19208 14940 19214 14952
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 19208 14912 20085 14940
rect 19208 14900 19214 14912
rect 20073 14909 20085 14912
rect 20119 14909 20131 14943
rect 20622 14940 20628 14952
rect 20583 14912 20628 14940
rect 20073 14903 20131 14909
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 21177 14943 21235 14949
rect 21177 14909 21189 14943
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 15948 14844 16528 14872
rect 16577 14875 16635 14881
rect 14700 14776 14872 14804
rect 15197 14807 15255 14813
rect 14700 14764 14706 14776
rect 15197 14773 15209 14807
rect 15243 14804 15255 14807
rect 15286 14804 15292 14816
rect 15243 14776 15292 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 15948 14813 15976 14844
rect 16577 14841 16589 14875
rect 16623 14872 16635 14875
rect 16623 14844 18092 14872
rect 16623 14841 16635 14844
rect 16577 14835 16635 14841
rect 18064 14813 18092 14844
rect 18230 14832 18236 14884
rect 18288 14872 18294 14884
rect 18509 14875 18567 14881
rect 18509 14872 18521 14875
rect 18288 14844 18521 14872
rect 18288 14832 18294 14844
rect 18509 14841 18521 14844
rect 18555 14872 18567 14875
rect 20714 14872 20720 14884
rect 18555 14844 20720 14872
rect 18555 14841 18567 14844
rect 18509 14835 18567 14841
rect 20714 14832 20720 14844
rect 20772 14832 20778 14884
rect 15933 14807 15991 14813
rect 15933 14804 15945 14807
rect 15436 14776 15945 14804
rect 15436 14764 15442 14776
rect 15933 14773 15945 14776
rect 15979 14773 15991 14807
rect 15933 14767 15991 14773
rect 16669 14807 16727 14813
rect 16669 14773 16681 14807
rect 16715 14804 16727 14807
rect 17037 14807 17095 14813
rect 17037 14804 17049 14807
rect 16715 14776 17049 14804
rect 16715 14773 16727 14776
rect 16669 14767 16727 14773
rect 17037 14773 17049 14776
rect 17083 14773 17095 14807
rect 17037 14767 17095 14773
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14773 18107 14807
rect 18049 14767 18107 14773
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 21192 14804 21220 14903
rect 20496 14776 21220 14804
rect 20496 14764 20502 14776
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2317 14603 2375 14609
rect 2317 14569 2329 14603
rect 2363 14600 2375 14603
rect 2774 14600 2780 14612
rect 2363 14572 2780 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 8202 14600 8208 14612
rect 7340 14572 8208 14600
rect 7340 14560 7346 14572
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 8757 14603 8815 14609
rect 8757 14600 8769 14603
rect 8444 14572 8769 14600
rect 8444 14560 8450 14572
rect 8757 14569 8769 14572
rect 8803 14569 8815 14603
rect 8757 14563 8815 14569
rect 9217 14603 9275 14609
rect 9217 14569 9229 14603
rect 9263 14600 9275 14603
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 9263 14572 9689 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 10100 14572 10149 14600
rect 10100 14560 10106 14572
rect 10137 14569 10149 14572
rect 10183 14600 10195 14603
rect 10502 14600 10508 14612
rect 10183 14572 10508 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12434 14600 12440 14612
rect 12299 14572 12440 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 4080 14504 5396 14532
rect 4080 14476 4108 14504
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14433 1823 14467
rect 1765 14427 1823 14433
rect 1780 14396 1808 14427
rect 1854 14424 1860 14476
rect 1912 14464 1918 14476
rect 2133 14467 2191 14473
rect 2133 14464 2145 14467
rect 1912 14436 2145 14464
rect 1912 14424 1918 14436
rect 2133 14433 2145 14436
rect 2179 14433 2191 14467
rect 4062 14464 4068 14476
rect 4023 14436 4068 14464
rect 2133 14427 2191 14433
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4332 14467 4390 14473
rect 4332 14464 4344 14467
rect 4212 14436 4344 14464
rect 4212 14424 4218 14436
rect 4332 14433 4344 14436
rect 4378 14464 4390 14467
rect 5258 14464 5264 14476
rect 4378 14436 5264 14464
rect 4378 14433 4390 14436
rect 4332 14427 4390 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 2314 14396 2320 14408
rect 1780 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 5368 14396 5396 14504
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 5782 14535 5840 14541
rect 5782 14532 5794 14535
rect 5592 14504 5794 14532
rect 5592 14492 5598 14504
rect 5782 14501 5794 14504
rect 5828 14501 5840 14535
rect 5782 14495 5840 14501
rect 7552 14535 7610 14541
rect 7552 14501 7564 14535
rect 7598 14532 7610 14535
rect 7598 14504 10364 14532
rect 7598 14501 7610 14504
rect 7552 14495 7610 14501
rect 7190 14464 7196 14476
rect 6932 14436 7196 14464
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 5368 14368 5549 14396
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 6932 14337 6960 14436
rect 7190 14424 7196 14436
rect 7248 14464 7254 14476
rect 7567 14464 7595 14495
rect 9122 14464 9128 14476
rect 7248 14436 7595 14464
rect 9083 14436 9128 14464
rect 7248 14424 7254 14436
rect 9122 14424 9128 14436
rect 9180 14424 9186 14476
rect 9490 14424 9496 14476
rect 9548 14464 9554 14476
rect 9766 14464 9772 14476
rect 9548 14436 9772 14464
rect 9548 14424 9554 14436
rect 9766 14424 9772 14436
rect 9824 14464 9830 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9824 14436 10057 14464
rect 9824 14424 9830 14436
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 10336 14408 10364 14504
rect 10410 14492 10416 14544
rect 10468 14532 10474 14544
rect 12268 14532 12296 14563
rect 12434 14560 12440 14572
rect 12492 14600 12498 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 12492 14572 14197 14600
rect 12492 14560 12498 14572
rect 14185 14569 14197 14572
rect 14231 14569 14243 14603
rect 14185 14563 14243 14569
rect 14369 14603 14427 14609
rect 14369 14569 14381 14603
rect 14415 14600 14427 14603
rect 19150 14600 19156 14612
rect 14415 14572 19156 14600
rect 14415 14569 14427 14572
rect 14369 14563 14427 14569
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 19889 14603 19947 14609
rect 19889 14569 19901 14603
rect 19935 14600 19947 14603
rect 20622 14600 20628 14612
rect 19935 14572 20628 14600
rect 19935 14569 19947 14572
rect 19889 14563 19947 14569
rect 10468 14504 12296 14532
rect 16936 14535 16994 14541
rect 10468 14492 10474 14504
rect 16936 14501 16948 14535
rect 16982 14532 16994 14535
rect 19812 14532 19840 14563
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 21085 14603 21143 14609
rect 21085 14569 21097 14603
rect 21131 14600 21143 14603
rect 21174 14600 21180 14612
rect 21131 14572 21180 14600
rect 21131 14569 21143 14572
rect 21085 14563 21143 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 16982 14504 20484 14532
rect 16982 14501 16994 14504
rect 16936 14495 16994 14501
rect 12980 14467 13038 14473
rect 12980 14433 12992 14467
rect 13026 14464 13038 14467
rect 13538 14464 13544 14476
rect 13026 14436 13544 14464
rect 13026 14433 13038 14436
rect 12980 14427 13038 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 14734 14464 14740 14476
rect 14695 14436 14740 14464
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16574 14464 16580 14476
rect 16071 14436 16580 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 16724 14436 18429 14464
rect 16724 14424 16730 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 18684 14467 18742 14473
rect 18684 14433 18696 14467
rect 18730 14464 18742 14467
rect 19426 14464 19432 14476
rect 18730 14436 19432 14464
rect 18730 14433 18742 14436
rect 18684 14427 18742 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19702 14424 19708 14476
rect 19760 14464 19766 14476
rect 20257 14467 20315 14473
rect 20257 14464 20269 14467
rect 19760 14436 20269 14464
rect 19760 14424 19766 14436
rect 20257 14433 20269 14436
rect 20303 14433 20315 14467
rect 20257 14427 20315 14433
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8680 14368 9321 14396
rect 8680 14337 8708 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 10318 14396 10324 14408
rect 10279 14368 10324 14396
rect 9309 14359 9367 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 10612 14368 12357 14396
rect 6917 14331 6975 14337
rect 6917 14297 6929 14331
rect 6963 14297 6975 14331
rect 6917 14291 6975 14297
rect 8665 14331 8723 14337
rect 8665 14297 8677 14331
rect 8711 14297 8723 14331
rect 8665 14291 8723 14297
rect 5445 14263 5503 14269
rect 5445 14229 5457 14263
rect 5491 14260 5503 14263
rect 5718 14260 5724 14272
rect 5491 14232 5724 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 8202 14220 8208 14272
rect 8260 14260 8266 14272
rect 8680 14260 8708 14291
rect 8260 14232 8708 14260
rect 8260 14220 8266 14232
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10612 14260 10640 14368
rect 12345 14365 12357 14368
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12713 14399 12771 14405
rect 12492 14368 12537 14396
rect 12492 14356 12498 14368
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 10870 14288 10876 14340
rect 10928 14328 10934 14340
rect 12066 14328 12072 14340
rect 10928 14300 12072 14328
rect 10928 14288 10934 14300
rect 12066 14288 12072 14300
rect 12124 14328 12130 14340
rect 12728 14328 12756 14359
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 13780 14368 14841 14396
rect 13780 14356 13786 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 15286 14396 15292 14408
rect 15059 14368 15292 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15488 14368 16129 14396
rect 12124 14300 12756 14328
rect 12124 14288 12130 14300
rect 10100 14232 10640 14260
rect 11885 14263 11943 14269
rect 10100 14220 10106 14232
rect 11885 14229 11897 14263
rect 11931 14260 11943 14263
rect 12526 14260 12532 14272
rect 11931 14232 12532 14260
rect 11931 14229 11943 14232
rect 11885 14223 11943 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 14090 14260 14096 14272
rect 14051 14232 14096 14260
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 14642 14220 14648 14272
rect 14700 14260 14706 14272
rect 15488 14269 15516 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 16298 14396 16304 14408
rect 16211 14368 16304 14396
rect 16117 14359 16175 14365
rect 16132 14328 16160 14359
rect 16298 14356 16304 14368
rect 16356 14396 16362 14408
rect 18230 14396 18236 14408
rect 16356 14368 16620 14396
rect 18191 14368 18236 14396
rect 16356 14356 16362 14368
rect 16482 14328 16488 14340
rect 16132 14300 16488 14328
rect 16482 14288 16488 14300
rect 16540 14288 16546 14340
rect 15473 14263 15531 14269
rect 15473 14260 15485 14263
rect 14700 14232 15485 14260
rect 14700 14220 14706 14232
rect 15473 14229 15485 14232
rect 15519 14229 15531 14263
rect 15654 14260 15660 14272
rect 15615 14232 15660 14260
rect 15473 14223 15531 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 16592 14260 16620 14368
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 20456 14405 20484 14504
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21174 14464 21180 14476
rect 20947 14436 21180 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 20349 14399 20407 14405
rect 20349 14396 20361 14399
rect 19576 14368 20361 14396
rect 19576 14356 19582 14368
rect 20349 14365 20361 14368
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 18049 14263 18107 14269
rect 18049 14260 18061 14263
rect 16592 14232 18061 14260
rect 18049 14229 18061 14232
rect 18095 14229 18107 14263
rect 18049 14223 18107 14229
rect 19610 14220 19616 14272
rect 19668 14260 19674 14272
rect 20438 14260 20444 14272
rect 19668 14232 20444 14260
rect 19668 14220 19674 14232
rect 20438 14220 20444 14232
rect 20496 14260 20502 14272
rect 21269 14263 21327 14269
rect 21269 14260 21281 14263
rect 20496 14232 21281 14260
rect 20496 14220 20502 14232
rect 21269 14229 21281 14232
rect 21315 14229 21327 14263
rect 21269 14223 21327 14229
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 3513 14059 3571 14065
rect 3513 14025 3525 14059
rect 3559 14056 3571 14059
rect 4246 14056 4252 14068
rect 3559 14028 4252 14056
rect 3559 14025 3571 14028
rect 3513 14019 3571 14025
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 4856 14028 5181 14056
rect 4856 14016 4862 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 5718 14056 5724 14068
rect 5169 14019 5227 14025
rect 5276 14028 5724 14056
rect 5276 13988 5304 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7064 14028 8340 14056
rect 7064 14016 7070 14028
rect 6822 13988 6828 14000
rect 4172 13960 5304 13988
rect 5644 13960 6828 13988
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2314 13920 2320 13932
rect 2275 13892 2320 13920
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 4172 13929 4200 13960
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13920 5043 13923
rect 5258 13920 5264 13932
rect 5031 13892 5264 13920
rect 5031 13889 5043 13892
rect 4985 13883 5043 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 5644 13929 5672 13960
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 8312 13988 8340 14028
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8536 14028 8769 14056
rect 8536 14016 8542 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 8938 14056 8944 14068
rect 8899 14028 8944 14056
rect 8757 14019 8815 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9122 14056 9128 14068
rect 9083 14028 9128 14056
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 10428 14028 11928 14056
rect 10428 13988 10456 14028
rect 8312 13960 10456 13988
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5718 13880 5724 13932
rect 5776 13920 5782 13932
rect 9674 13920 9680 13932
rect 5776 13892 5821 13920
rect 8680 13892 9680 13920
rect 5776 13880 5782 13892
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 3326 13852 3332 13864
rect 2179 13824 3332 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13852 4031 13855
rect 4614 13852 4620 13864
rect 4019 13824 4620 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 5902 13852 5908 13864
rect 5583 13824 5908 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 7340 13824 7389 13852
rect 7340 13812 7346 13824
rect 7377 13821 7389 13824
rect 7423 13852 7435 13855
rect 7644 13855 7702 13861
rect 7423 13824 7604 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 3881 13787 3939 13793
rect 3881 13753 3893 13787
rect 3927 13784 3939 13787
rect 4706 13784 4712 13796
rect 3927 13756 4384 13784
rect 4667 13756 4712 13784
rect 3927 13753 3939 13756
rect 3881 13747 3939 13753
rect 4356 13725 4384 13756
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 7576 13784 7604 13824
rect 7644 13821 7656 13855
rect 7690 13852 7702 13855
rect 8202 13852 8208 13864
rect 7690 13824 8208 13852
rect 7690 13821 7702 13824
rect 7644 13815 7702 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8680 13852 8708 13892
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10318 13920 10324 13932
rect 9815 13892 10324 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 10502 13920 10508 13932
rect 10463 13892 10508 13920
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 10735 13892 11008 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 8312 13824 8708 13852
rect 8312 13784 8340 13824
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 8812 13824 9505 13852
rect 8812 13812 8818 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 10410 13852 10416 13864
rect 9631 13824 10416 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 7576 13756 8340 13784
rect 9508 13784 9536 13815
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 10870 13852 10876 13864
rect 10831 13824 10876 13852
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 10980 13852 11008 13892
rect 11900 13852 11928 14028
rect 13280 14028 14473 14056
rect 12805 13991 12863 13997
rect 12805 13957 12817 13991
rect 12851 13957 12863 13991
rect 12805 13951 12863 13957
rect 12710 13852 12716 13864
rect 10980 13824 11100 13852
rect 11900 13824 12716 13852
rect 10042 13784 10048 13796
rect 9508 13756 10048 13784
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 11072 13784 11100 13824
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 12820 13852 12848 13951
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 13280 13929 13308 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 14792 14028 14933 14056
rect 14792 14016 14798 14028
rect 14921 14025 14933 14028
rect 14967 14025 14979 14059
rect 14921 14019 14979 14025
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 17126 14056 17132 14068
rect 16540 14028 17132 14056
rect 16540 14016 16546 14028
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 19518 14056 19524 14068
rect 19479 14028 19524 14056
rect 19518 14016 19524 14028
rect 19576 14016 19582 14068
rect 21082 14056 21088 14068
rect 21043 14028 21088 14056
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 13538 13988 13544 14000
rect 13372 13960 13544 13988
rect 13372 13929 13400 13960
rect 13538 13948 13544 13960
rect 13596 13988 13602 14000
rect 13596 13960 16344 13988
rect 13596 13948 13602 13960
rect 16316 13932 16344 13960
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 18046 13988 18052 14000
rect 16448 13960 18052 13988
rect 16448 13948 16454 13960
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 19426 13988 19432 14000
rect 19387 13960 19432 13988
rect 19426 13948 19432 13960
rect 19484 13988 19490 14000
rect 20622 13988 20628 14000
rect 19484 13960 20628 13988
rect 19484 13948 19490 13960
rect 13265 13923 13323 13929
rect 13265 13920 13277 13923
rect 12952 13892 13277 13920
rect 12952 13880 12958 13892
rect 13265 13889 13277 13892
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 14148 13892 14289 13920
rect 14148 13880 14154 13892
rect 14277 13889 14289 13892
rect 14323 13920 14335 13923
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 14323 13892 15485 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 16298 13920 16304 13932
rect 16259 13892 16304 13920
rect 15473 13883 15531 13889
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 20088 13929 20116 13960
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19208 13892 19993 13920
rect 19208 13880 19214 13892
rect 19981 13889 19993 13892
rect 20027 13889 20039 13923
rect 19981 13883 20039 13889
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13889 20131 13923
rect 20073 13883 20131 13889
rect 14182 13852 14188 13864
rect 12820 13824 14044 13852
rect 11146 13793 11152 13796
rect 11140 13784 11152 13793
rect 11072 13756 11152 13784
rect 11140 13747 11152 13756
rect 11146 13744 11152 13747
rect 11204 13744 11210 13796
rect 13173 13787 13231 13793
rect 13173 13753 13185 13787
rect 13219 13784 13231 13787
rect 13906 13784 13912 13796
rect 13219 13756 13912 13784
rect 13219 13753 13231 13756
rect 13173 13747 13231 13753
rect 13906 13744 13912 13756
rect 13964 13744 13970 13796
rect 14016 13793 14044 13824
rect 14108 13824 14188 13852
rect 14108 13793 14136 13824
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15289 13855 15347 13861
rect 14875 13824 15240 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15212 13796 15240 13824
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15654 13852 15660 13864
rect 15335 13824 15660 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17880 13824 18061 13852
rect 14001 13787 14059 13793
rect 14001 13753 14013 13787
rect 14047 13753 14059 13787
rect 14001 13747 14059 13753
rect 14093 13787 14151 13793
rect 14093 13753 14105 13787
rect 14139 13753 14151 13787
rect 15194 13784 15200 13796
rect 15107 13756 15200 13784
rect 14093 13747 14151 13753
rect 15194 13744 15200 13756
rect 15252 13784 15258 13796
rect 16117 13787 16175 13793
rect 16117 13784 16129 13787
rect 15252 13756 16129 13784
rect 15252 13744 15258 13756
rect 16117 13753 16129 13756
rect 16163 13784 16175 13787
rect 16390 13784 16396 13796
rect 16163 13756 16396 13784
rect 16163 13753 16175 13756
rect 16117 13747 16175 13753
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 16574 13784 16580 13796
rect 16535 13756 16580 13784
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 16666 13744 16672 13796
rect 16724 13784 16730 13796
rect 17880 13784 17908 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 20349 13855 20407 13861
rect 20349 13852 20361 13855
rect 19392 13824 20361 13852
rect 19392 13812 19398 13824
rect 20349 13821 20361 13824
rect 20395 13821 20407 13855
rect 20349 13815 20407 13821
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13852 20683 13855
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 20671 13824 20913 13852
rect 20671 13821 20683 13824
rect 20625 13815 20683 13821
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 16724 13756 17908 13784
rect 16724 13744 16730 13756
rect 18138 13744 18144 13796
rect 18196 13784 18202 13796
rect 18316 13787 18374 13793
rect 18316 13784 18328 13787
rect 18196 13756 18328 13784
rect 18196 13744 18202 13756
rect 18316 13753 18328 13756
rect 18362 13784 18374 13787
rect 19794 13784 19800 13796
rect 18362 13756 19800 13784
rect 18362 13753 18374 13756
rect 18316 13747 18374 13753
rect 19794 13744 19800 13756
rect 19852 13744 19858 13796
rect 4341 13719 4399 13725
rect 4341 13685 4353 13719
rect 4387 13685 4399 13719
rect 4798 13716 4804 13728
rect 4759 13688 4804 13716
rect 4341 13679 4399 13685
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 7374 13676 7380 13728
rect 7432 13716 7438 13728
rect 8754 13716 8760 13728
rect 7432 13688 8760 13716
rect 7432 13676 7438 13688
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 9824 13688 10425 13716
rect 9824 13676 9830 13688
rect 10413 13685 10425 13688
rect 10459 13685 10471 13719
rect 12250 13716 12256 13728
rect 12211 13688 12256 13716
rect 10413 13679 10471 13685
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 13633 13719 13691 13725
rect 13633 13685 13645 13719
rect 13679 13716 13691 13719
rect 13722 13716 13728 13728
rect 13679 13688 13728 13716
rect 13679 13685 13691 13688
rect 13633 13679 13691 13685
rect 13722 13676 13728 13688
rect 13780 13676 13786 13728
rect 15381 13719 15439 13725
rect 15381 13685 15393 13719
rect 15427 13716 15439 13719
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15427 13688 15761 13716
rect 15427 13685 15439 13688
rect 15381 13679 15439 13685
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 16209 13719 16267 13725
rect 16209 13685 16221 13719
rect 16255 13716 16267 13719
rect 16945 13719 17003 13725
rect 16945 13716 16957 13719
rect 16255 13688 16957 13716
rect 16255 13685 16267 13688
rect 16209 13679 16267 13685
rect 16945 13685 16957 13688
rect 16991 13716 17003 13719
rect 17126 13716 17132 13728
rect 16991 13688 17132 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 19886 13716 19892 13728
rect 19847 13688 19892 13716
rect 19886 13676 19892 13688
rect 19944 13676 19950 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 3697 13515 3755 13521
rect 3697 13481 3709 13515
rect 3743 13512 3755 13515
rect 4154 13512 4160 13524
rect 3743 13484 4160 13512
rect 3743 13481 3755 13484
rect 3697 13475 3755 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 4764 13484 5457 13512
rect 4764 13472 4770 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5445 13475 5503 13481
rect 5997 13515 6055 13521
rect 5997 13481 6009 13515
rect 6043 13481 6055 13515
rect 5997 13475 6055 13481
rect 4246 13444 4252 13456
rect 4159 13416 4252 13444
rect 4246 13404 4252 13416
rect 4304 13444 4310 13456
rect 4798 13444 4804 13456
rect 4304 13416 4804 13444
rect 4304 13404 4310 13416
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 5077 13447 5135 13453
rect 5077 13444 5089 13447
rect 4908 13416 5089 13444
rect 2584 13379 2642 13385
rect 2584 13345 2596 13379
rect 2630 13376 2642 13379
rect 2958 13376 2964 13388
rect 2630 13348 2964 13376
rect 2630 13345 2642 13348
rect 2584 13339 2642 13345
rect 2958 13336 2964 13348
rect 3016 13336 3022 13388
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4908 13376 4936 13416
rect 5077 13413 5089 13416
rect 5123 13444 5135 13447
rect 5721 13447 5779 13453
rect 5721 13444 5733 13447
rect 5123 13416 5733 13444
rect 5123 13413 5135 13416
rect 5077 13407 5135 13413
rect 5721 13413 5733 13416
rect 5767 13413 5779 13447
rect 6012 13444 6040 13475
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7190 13512 7196 13524
rect 6972 13484 7196 13512
rect 6972 13472 6978 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7285 13515 7343 13521
rect 7285 13481 7297 13515
rect 7331 13512 7343 13515
rect 7374 13512 7380 13524
rect 7331 13484 7380 13512
rect 7331 13481 7343 13484
rect 7285 13475 7343 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 7653 13515 7711 13521
rect 7653 13481 7665 13515
rect 7699 13512 7711 13515
rect 7742 13512 7748 13524
rect 7699 13484 7748 13512
rect 7699 13481 7711 13484
rect 7653 13475 7711 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8754 13512 8760 13524
rect 8715 13484 8760 13512
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9766 13512 9772 13524
rect 9727 13484 9772 13512
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10229 13515 10287 13521
rect 10229 13481 10241 13515
rect 10275 13512 10287 13515
rect 10410 13512 10416 13524
rect 10275 13484 10416 13512
rect 10275 13481 10287 13484
rect 10229 13475 10287 13481
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 14182 13512 14188 13524
rect 11020 13484 13768 13512
rect 14143 13484 14188 13512
rect 11020 13472 11026 13484
rect 8021 13447 8079 13453
rect 8021 13444 8033 13447
rect 6012 13416 8033 13444
rect 5721 13407 5779 13413
rect 8021 13413 8033 13416
rect 8067 13413 8079 13447
rect 10042 13444 10048 13456
rect 8021 13407 8079 13413
rect 8588 13416 8800 13444
rect 10003 13416 10048 13444
rect 4396 13348 4936 13376
rect 4985 13379 5043 13385
rect 4396 13336 4402 13348
rect 4985 13345 4997 13379
rect 5031 13345 5043 13379
rect 4985 13339 5043 13345
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 2317 13311 2375 13317
rect 2317 13308 2329 13311
rect 1728 13280 2329 13308
rect 1728 13268 1734 13280
rect 2317 13277 2329 13280
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 4433 13175 4491 13181
rect 4433 13172 4445 13175
rect 4396 13144 4445 13172
rect 4396 13132 4402 13144
rect 4433 13141 4445 13144
rect 4479 13172 4491 13175
rect 5000 13172 5028 13339
rect 5258 13308 5264 13320
rect 5219 13280 5264 13308
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5736 13240 5764 13407
rect 6362 13376 6368 13388
rect 6323 13348 6368 13376
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 8588 13376 8616 13416
rect 6564 13348 8616 13376
rect 8665 13379 8723 13385
rect 5902 13268 5908 13320
rect 5960 13308 5966 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 5960 13280 6469 13308
rect 5960 13268 5966 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6564 13240 6592 13348
rect 8665 13345 8677 13379
rect 8711 13345 8723 13379
rect 8772 13376 8800 13416
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10505 13447 10563 13453
rect 10505 13413 10517 13447
rect 10551 13444 10563 13447
rect 10594 13444 10600 13456
rect 10551 13416 10600 13444
rect 10551 13413 10563 13416
rect 10505 13407 10563 13413
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 12066 13404 12072 13456
rect 12124 13444 12130 13456
rect 12124 13416 12572 13444
rect 12124 13404 12130 13416
rect 12434 13376 12440 13388
rect 8772 13348 12440 13376
rect 8665 13339 8723 13345
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13308 6699 13311
rect 7282 13308 7288 13320
rect 6687 13280 7288 13308
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 7282 13268 7288 13280
rect 7340 13308 7346 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7340 13280 7389 13308
rect 7340 13268 7346 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 5736 13212 6592 13240
rect 6825 13243 6883 13249
rect 6825 13209 6837 13243
rect 6871 13240 6883 13243
rect 8128 13240 8156 13271
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8260 13280 8305 13308
rect 8260 13268 8266 13280
rect 6871 13212 8156 13240
rect 8680 13240 8708 13339
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 12544 13376 12572 13416
rect 12612 13379 12670 13385
rect 12612 13376 12624 13379
rect 12544 13348 12624 13376
rect 12612 13345 12624 13348
rect 12658 13376 12670 13379
rect 13740 13376 13768 13484
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 14734 13472 14740 13524
rect 14792 13512 14798 13524
rect 19521 13515 19579 13521
rect 14792 13484 19472 13512
rect 14792 13472 14798 13484
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 14645 13447 14703 13453
rect 14645 13444 14657 13447
rect 14056 13416 14657 13444
rect 14056 13404 14062 13416
rect 14645 13413 14657 13416
rect 14691 13413 14703 13447
rect 14645 13407 14703 13413
rect 15286 13404 15292 13456
rect 15344 13444 15350 13456
rect 15534 13447 15592 13453
rect 15534 13444 15546 13447
rect 15344 13416 15546 13444
rect 15344 13404 15350 13416
rect 15534 13413 15546 13416
rect 15580 13413 15592 13447
rect 15534 13407 15592 13413
rect 16666 13404 16672 13456
rect 16724 13444 16730 13456
rect 17954 13444 17960 13456
rect 16724 13416 17960 13444
rect 16724 13404 16730 13416
rect 17954 13404 17960 13416
rect 18012 13404 18018 13456
rect 19444 13444 19472 13484
rect 19521 13481 19533 13515
rect 19567 13512 19579 13515
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 19567 13484 19993 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 20438 13512 20444 13524
rect 20399 13484 20444 13512
rect 19981 13475 20039 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 21174 13444 21180 13456
rect 19444 13416 20944 13444
rect 21135 13416 21180 13444
rect 17120 13379 17178 13385
rect 12658 13348 13400 13376
rect 13740 13348 16436 13376
rect 12658 13345 12670 13348
rect 12612 13339 12670 13345
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 11698 13308 11704 13320
rect 9272 13280 11704 13308
rect 9272 13268 9278 13280
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 12342 13308 12348 13320
rect 12303 13280 12348 13308
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 11790 13240 11796 13252
rect 8680 13212 11796 13240
rect 6871 13209 6883 13212
rect 6825 13203 6883 13209
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 13372 13240 13400 13348
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13504 13280 14289 13308
rect 13504 13268 13510 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 15286 13308 15292 13320
rect 14424 13280 14469 13308
rect 15247 13280 15292 13308
rect 14424 13268 14430 13280
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16408 13240 16436 13348
rect 17120 13345 17132 13379
rect 17166 13376 17178 13379
rect 17494 13376 17500 13388
rect 17166 13348 17500 13376
rect 17166 13345 17178 13348
rect 17120 13339 17178 13345
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 20349 13379 20407 13385
rect 19812 13348 20300 13376
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16853 13311 16911 13317
rect 16853 13308 16865 13311
rect 16632 13280 16865 13308
rect 16632 13268 16638 13280
rect 16853 13277 16865 13280
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18782 13308 18788 13320
rect 18012 13280 18788 13308
rect 18012 13268 18018 13280
rect 18782 13268 18788 13280
rect 18840 13308 18846 13320
rect 18969 13311 19027 13317
rect 18969 13308 18981 13311
rect 18840 13280 18981 13308
rect 18840 13268 18846 13280
rect 18969 13277 18981 13280
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 19242 13268 19248 13320
rect 19300 13308 19306 13320
rect 19812 13317 19840 13348
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19300 13280 19625 13308
rect 19300 13268 19306 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 13372 13212 15148 13240
rect 16408 13212 16804 13240
rect 15120 13184 15148 13212
rect 4479 13144 5028 13172
rect 4479 13141 4491 13144
rect 4433 13135 4491 13141
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 7708 13144 8493 13172
rect 7708 13132 7714 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 10502 13132 10508 13184
rect 10560 13172 10566 13184
rect 11882 13172 11888 13184
rect 10560 13144 11888 13172
rect 10560 13132 10566 13144
rect 11882 13132 11888 13144
rect 11940 13172 11946 13184
rect 13538 13172 13544 13184
rect 11940 13144 13544 13172
rect 11940 13132 11946 13144
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 13722 13172 13728 13184
rect 13683 13144 13728 13172
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 13817 13175 13875 13181
rect 13817 13141 13829 13175
rect 13863 13172 13875 13175
rect 14734 13172 14740 13184
rect 13863 13144 14740 13172
rect 13863 13141 13875 13144
rect 13817 13135 13875 13141
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 15102 13132 15108 13184
rect 15160 13172 15166 13184
rect 16669 13175 16727 13181
rect 16669 13172 16681 13175
rect 15160 13144 16681 13172
rect 15160 13132 15166 13144
rect 16669 13141 16681 13144
rect 16715 13141 16727 13175
rect 16776 13172 16804 13212
rect 18046 13200 18052 13252
rect 18104 13240 18110 13252
rect 19153 13243 19211 13249
rect 18104 13212 19104 13240
rect 18104 13200 18110 13212
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 16776 13144 18245 13172
rect 16669 13135 16727 13141
rect 18233 13141 18245 13144
rect 18279 13172 18291 13175
rect 18690 13172 18696 13184
rect 18279 13144 18696 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 19076 13172 19104 13212
rect 19153 13209 19165 13243
rect 19199 13240 19211 13243
rect 19702 13240 19708 13252
rect 19199 13212 19708 13240
rect 19199 13209 19211 13212
rect 19153 13203 19211 13209
rect 19702 13200 19708 13212
rect 19760 13200 19766 13252
rect 20272 13240 20300 13348
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 20806 13376 20812 13388
rect 20395 13348 20812 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 20916 13385 20944 13416
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 20901 13379 20959 13385
rect 20901 13345 20913 13379
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 20438 13268 20444 13320
rect 20496 13308 20502 13320
rect 20533 13311 20591 13317
rect 20533 13308 20545 13311
rect 20496 13280 20545 13308
rect 20496 13268 20502 13280
rect 20533 13277 20545 13280
rect 20579 13277 20591 13311
rect 20533 13271 20591 13277
rect 20622 13240 20628 13252
rect 20272 13212 20628 13240
rect 20622 13200 20628 13212
rect 20680 13200 20686 13252
rect 20990 13172 20996 13184
rect 19076 13144 20996 13172
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1397 12971 1455 12977
rect 1397 12937 1409 12971
rect 1443 12968 1455 12971
rect 1578 12968 1584 12980
rect 1443 12940 1584 12968
rect 1443 12937 1455 12940
rect 1397 12931 1455 12937
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 3694 12928 3700 12980
rect 3752 12968 3758 12980
rect 3881 12971 3939 12977
rect 3881 12968 3893 12971
rect 3752 12940 3893 12968
rect 3752 12928 3758 12940
rect 3881 12937 3893 12940
rect 3927 12937 3939 12971
rect 3881 12931 3939 12937
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 4120 12940 9536 12968
rect 4120 12928 4126 12940
rect 5166 12860 5172 12912
rect 5224 12900 5230 12912
rect 5902 12900 5908 12912
rect 5224 12872 5908 12900
rect 5224 12860 5230 12872
rect 5902 12860 5908 12872
rect 5960 12860 5966 12912
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 2056 12764 2084 12795
rect 2498 12792 2504 12844
rect 2556 12832 2562 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2556 12804 2789 12832
rect 2556 12792 2562 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 3786 12792 3792 12844
rect 3844 12832 3850 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 3844 12804 4077 12832
rect 3844 12792 3850 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 5316 12804 5365 12832
rect 5316 12792 5322 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 6362 12792 6368 12844
rect 6420 12832 6426 12844
rect 6457 12835 6515 12841
rect 6457 12832 6469 12835
rect 6420 12804 6469 12832
rect 6420 12792 6426 12804
rect 6457 12801 6469 12804
rect 6503 12801 6515 12835
rect 6457 12795 6515 12801
rect 8110 12792 8116 12844
rect 8168 12832 8174 12844
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 8168 12804 8309 12832
rect 8168 12792 8174 12804
rect 8297 12801 8309 12804
rect 8343 12832 8355 12835
rect 9508 12832 9536 12940
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11204 12940 11345 12968
rect 11204 12928 11210 12940
rect 11333 12937 11345 12940
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 12437 12971 12495 12977
rect 12437 12968 12449 12971
rect 11756 12940 12449 12968
rect 11756 12928 11762 12940
rect 12437 12937 12449 12940
rect 12483 12937 12495 12971
rect 13446 12968 13452 12980
rect 13407 12940 13452 12968
rect 12437 12931 12495 12937
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13538 12928 13544 12980
rect 13596 12968 13602 12980
rect 18782 12968 18788 12980
rect 13596 12940 18788 12968
rect 13596 12928 13602 12940
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 19061 12971 19119 12977
rect 19061 12968 19073 12971
rect 19024 12940 19073 12968
rect 19024 12928 19030 12940
rect 19061 12937 19073 12940
rect 19107 12937 19119 12971
rect 19242 12968 19248 12980
rect 19203 12940 19248 12968
rect 19061 12931 19119 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 19886 12928 19892 12980
rect 19944 12968 19950 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 19944 12940 20085 12968
rect 19944 12928 19950 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 9861 12903 9919 12909
rect 9861 12869 9873 12903
rect 9907 12900 9919 12903
rect 9950 12900 9956 12912
rect 9907 12872 9956 12900
rect 9907 12869 9919 12872
rect 9861 12863 9919 12869
rect 9950 12860 9956 12872
rect 10008 12860 10014 12912
rect 12713 12903 12771 12909
rect 12713 12900 12725 12903
rect 10980 12872 12725 12900
rect 8343 12804 8616 12832
rect 9508 12804 10088 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 2958 12764 2964 12776
rect 2056 12736 2964 12764
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 6871 12736 8493 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7300 12708 7328 12736
rect 8481 12733 8493 12736
rect 8527 12733 8539 12767
rect 8588 12764 8616 12804
rect 8588 12736 8984 12764
rect 8481 12727 8539 12733
rect 2593 12699 2651 12705
rect 2593 12665 2605 12699
rect 2639 12696 2651 12699
rect 3050 12696 3056 12708
rect 2639 12668 3056 12696
rect 2639 12665 2651 12668
rect 2593 12659 2651 12665
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 5261 12699 5319 12705
rect 5261 12665 5273 12699
rect 5307 12696 5319 12699
rect 6086 12696 6092 12708
rect 5307 12668 6092 12696
rect 5307 12665 5319 12668
rect 5261 12659 5319 12665
rect 6086 12656 6092 12668
rect 6144 12656 6150 12708
rect 6270 12656 6276 12708
rect 6328 12696 6334 12708
rect 7070 12699 7128 12705
rect 7070 12696 7082 12699
rect 6328 12668 7082 12696
rect 6328 12656 6334 12668
rect 7070 12665 7082 12668
rect 7116 12665 7128 12699
rect 7070 12659 7128 12665
rect 7282 12656 7288 12708
rect 7340 12656 7346 12708
rect 7558 12656 7564 12708
rect 7616 12696 7622 12708
rect 8110 12696 8116 12708
rect 7616 12668 8116 12696
rect 7616 12656 7622 12668
rect 8110 12656 8116 12668
rect 8168 12656 8174 12708
rect 8754 12705 8760 12708
rect 8748 12696 8760 12705
rect 8220 12668 8760 12696
rect 1762 12628 1768 12640
rect 1723 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 1857 12631 1915 12637
rect 1857 12597 1869 12631
rect 1903 12628 1915 12631
rect 2225 12631 2283 12637
rect 2225 12628 2237 12631
rect 1903 12600 2237 12628
rect 1903 12597 1915 12600
rect 1857 12591 1915 12597
rect 2225 12597 2237 12600
rect 2271 12597 2283 12631
rect 2682 12628 2688 12640
rect 2643 12600 2688 12628
rect 2225 12591 2283 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 4798 12628 4804 12640
rect 4759 12600 4804 12628
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 8220 12637 8248 12668
rect 8748 12659 8760 12668
rect 8754 12656 8760 12659
rect 8812 12656 8818 12708
rect 5169 12631 5227 12637
rect 5169 12628 5181 12631
rect 4948 12600 5181 12628
rect 4948 12588 4954 12600
rect 5169 12597 5181 12600
rect 5215 12597 5227 12631
rect 5169 12591 5227 12597
rect 8205 12631 8263 12637
rect 8205 12597 8217 12631
rect 8251 12597 8263 12631
rect 8956 12628 8984 12736
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9674 12764 9680 12776
rect 9180 12736 9680 12764
rect 9180 12724 9186 12736
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 9824 12736 9965 12764
rect 9824 12724 9830 12736
rect 9953 12733 9965 12736
rect 9999 12733 10011 12767
rect 10060 12764 10088 12804
rect 10980 12764 11008 12872
rect 12713 12869 12725 12872
rect 12759 12869 12771 12903
rect 12713 12863 12771 12869
rect 12805 12903 12863 12909
rect 12805 12869 12817 12903
rect 12851 12900 12863 12903
rect 13630 12900 13636 12912
rect 12851 12872 13636 12900
rect 12851 12869 12863 12872
rect 12805 12863 12863 12869
rect 13630 12860 13636 12872
rect 13688 12900 13694 12912
rect 14553 12903 14611 12909
rect 14553 12900 14565 12903
rect 13688 12872 14565 12900
rect 13688 12860 13694 12872
rect 14553 12869 14565 12872
rect 14599 12869 14611 12903
rect 14553 12863 14611 12869
rect 18049 12903 18107 12909
rect 18049 12869 18061 12903
rect 18095 12900 18107 12903
rect 19702 12900 19708 12912
rect 18095 12872 19708 12900
rect 18095 12869 18107 12872
rect 18049 12863 18107 12869
rect 19702 12860 19708 12872
rect 19760 12860 19766 12912
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 11756 12804 11897 12832
rect 11756 12792 11762 12804
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 12066 12832 12072 12844
rect 12027 12804 12072 12832
rect 11885 12795 11943 12801
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 13722 12792 13728 12844
rect 13780 12832 13786 12844
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13780 12804 14013 12832
rect 13780 12792 13786 12804
rect 14001 12801 14013 12804
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15160 12804 15393 12832
rect 15160 12792 15166 12804
rect 15381 12801 15393 12804
rect 15427 12832 15439 12835
rect 15470 12832 15476 12844
rect 15427 12804 15476 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 17552 12804 18613 12832
rect 17552 12792 17558 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 19794 12832 19800 12844
rect 19755 12804 19800 12832
rect 18601 12795 18659 12801
rect 19794 12792 19800 12804
rect 19852 12832 19858 12844
rect 20438 12832 20444 12844
rect 19852 12804 20444 12832
rect 19852 12792 19858 12804
rect 20438 12792 20444 12804
rect 20496 12832 20502 12844
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20496 12804 20637 12832
rect 20496 12792 20502 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 20806 12792 20812 12844
rect 20864 12832 20870 12844
rect 20901 12835 20959 12841
rect 20901 12832 20913 12835
rect 20864 12804 20913 12832
rect 20864 12792 20870 12804
rect 20901 12801 20913 12804
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 10060 12736 11008 12764
rect 9953 12727 10011 12733
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 11848 12736 13001 12764
rect 11848 12724 11854 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 13814 12764 13820 12776
rect 13775 12736 13820 12764
rect 12989 12727 13047 12733
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 14461 12767 14519 12773
rect 14461 12733 14473 12767
rect 14507 12764 14519 12767
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 14507 12736 14565 12764
rect 14507 12733 14519 12736
rect 14461 12727 14519 12733
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 14553 12727 14611 12733
rect 14660 12736 15301 12764
rect 10220 12699 10278 12705
rect 10220 12665 10232 12699
rect 10266 12696 10278 12699
rect 10962 12696 10968 12708
rect 10266 12668 10968 12696
rect 10266 12665 10278 12668
rect 10220 12659 10278 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 14660 12705 14688 12736
rect 15289 12733 15301 12736
rect 15335 12764 15347 12767
rect 15335 12736 17356 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 13909 12699 13967 12705
rect 13909 12696 13921 12699
rect 11440 12668 13921 12696
rect 10502 12628 10508 12640
rect 8956 12600 10508 12628
rect 8205 12591 8263 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 11440 12637 11468 12668
rect 13909 12665 13921 12668
rect 13955 12665 13967 12699
rect 14645 12699 14703 12705
rect 14645 12696 14657 12699
rect 13909 12659 13967 12665
rect 14016 12668 14657 12696
rect 11425 12631 11483 12637
rect 11425 12597 11437 12631
rect 11471 12597 11483 12631
rect 11790 12628 11796 12640
rect 11751 12600 11796 12628
rect 11425 12591 11483 12597
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 12713 12631 12771 12637
rect 12713 12597 12725 12631
rect 12759 12628 12771 12631
rect 14016 12628 14044 12668
rect 14645 12665 14657 12668
rect 14691 12665 14703 12699
rect 14645 12659 14703 12665
rect 15197 12699 15255 12705
rect 15197 12665 15209 12699
rect 15243 12696 15255 12699
rect 15657 12699 15715 12705
rect 15657 12696 15669 12699
rect 15243 12668 15669 12696
rect 15243 12665 15255 12668
rect 15197 12659 15255 12665
rect 15657 12665 15669 12668
rect 15703 12665 15715 12699
rect 15657 12659 15715 12665
rect 12759 12600 14044 12628
rect 12759 12597 12771 12600
rect 12713 12591 12771 12597
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 14277 12631 14335 12637
rect 14277 12628 14289 12631
rect 14148 12600 14289 12628
rect 14148 12588 14154 12600
rect 14277 12597 14289 12600
rect 14323 12597 14335 12631
rect 14277 12591 14335 12597
rect 14734 12588 14740 12640
rect 14792 12628 14798 12640
rect 14829 12631 14887 12637
rect 14829 12628 14841 12631
rect 14792 12600 14841 12628
rect 14792 12588 14798 12600
rect 14829 12597 14841 12600
rect 14875 12597 14887 12631
rect 17328 12628 17356 12736
rect 17770 12724 17776 12776
rect 17828 12764 17834 12776
rect 18966 12764 18972 12776
rect 17828 12736 18972 12764
rect 17828 12724 17834 12736
rect 18966 12724 18972 12736
rect 19024 12764 19030 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19024 12736 19625 12764
rect 19024 12724 19030 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 20441 12699 20499 12705
rect 18196 12668 20392 12696
rect 18196 12656 18202 12668
rect 18046 12628 18052 12640
rect 17328 12600 18052 12628
rect 14829 12591 14887 12597
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18414 12628 18420 12640
rect 18375 12600 18420 12628
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18509 12631 18567 12637
rect 18509 12597 18521 12631
rect 18555 12628 18567 12631
rect 18598 12628 18604 12640
rect 18555 12600 18604 12628
rect 18555 12597 18567 12600
rect 18509 12591 18567 12597
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 19426 12628 19432 12640
rect 18932 12600 19432 12628
rect 18932 12588 18938 12600
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 19705 12631 19763 12637
rect 19705 12597 19717 12631
rect 19751 12628 19763 12631
rect 20070 12628 20076 12640
rect 19751 12600 20076 12628
rect 19751 12597 19763 12600
rect 19705 12591 19763 12597
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 20364 12628 20392 12668
rect 20441 12665 20453 12699
rect 20487 12696 20499 12699
rect 20714 12696 20720 12708
rect 20487 12668 20720 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 20714 12656 20720 12668
rect 20772 12696 20778 12708
rect 21361 12699 21419 12705
rect 21361 12696 21373 12699
rect 20772 12668 21373 12696
rect 20772 12656 20778 12668
rect 21361 12665 21373 12668
rect 21407 12665 21419 12699
rect 21361 12659 21419 12665
rect 20533 12631 20591 12637
rect 20533 12628 20545 12631
rect 20364 12600 20545 12628
rect 20533 12597 20545 12600
rect 20579 12628 20591 12631
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 20579 12600 21189 12628
rect 20579 12597 20591 12600
rect 20533 12591 20591 12597
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 21177 12591 21235 12597
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 2958 12424 2964 12436
rect 2919 12396 2964 12424
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3421 12427 3479 12433
rect 3108 12396 3153 12424
rect 3108 12384 3114 12396
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 3694 12424 3700 12436
rect 3467 12396 3700 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 3786 12384 3792 12436
rect 3844 12384 3850 12436
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 4798 12424 4804 12436
rect 4571 12396 4804 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 7745 12427 7803 12433
rect 7745 12393 7757 12427
rect 7791 12424 7803 12427
rect 9122 12424 9128 12436
rect 7791 12396 9128 12424
rect 7791 12393 7803 12396
rect 7745 12387 7803 12393
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 9548 12396 12388 12424
rect 9548 12384 9554 12396
rect 2498 12316 2504 12368
rect 2556 12316 2562 12368
rect 3513 12359 3571 12365
rect 3513 12325 3525 12359
rect 3559 12356 3571 12359
rect 3804 12356 3832 12384
rect 3559 12328 3832 12356
rect 5160 12359 5218 12365
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 5160 12325 5172 12359
rect 5206 12356 5218 12359
rect 5258 12356 5264 12368
rect 5206 12328 5264 12356
rect 5206 12325 5218 12328
rect 5160 12319 5218 12325
rect 5258 12316 5264 12328
rect 5316 12316 5322 12368
rect 6730 12316 6736 12368
rect 6788 12356 6794 12368
rect 7558 12356 7564 12368
rect 6788 12328 7564 12356
rect 6788 12316 6794 12328
rect 7558 12316 7564 12328
rect 7616 12356 7622 12368
rect 7653 12359 7711 12365
rect 7653 12356 7665 12359
rect 7616 12328 7665 12356
rect 7616 12316 7622 12328
rect 7653 12325 7665 12328
rect 7699 12325 7711 12359
rect 7653 12319 7711 12325
rect 8380 12359 8438 12365
rect 8380 12325 8392 12359
rect 8426 12356 8438 12359
rect 8478 12356 8484 12368
rect 8426 12328 8484 12356
rect 8426 12325 8438 12328
rect 8380 12319 8438 12325
rect 8478 12316 8484 12328
rect 8536 12316 8542 12368
rect 8754 12316 8760 12368
rect 8812 12356 8818 12368
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 8812 12328 9873 12356
rect 8812 12316 8818 12328
rect 9861 12325 9873 12328
rect 9907 12325 9919 12359
rect 10413 12359 10471 12365
rect 10413 12356 10425 12359
rect 9861 12319 9919 12325
rect 10051 12328 10425 12356
rect 1848 12291 1906 12297
rect 1848 12257 1860 12291
rect 1894 12288 1906 12291
rect 2222 12288 2228 12300
rect 1894 12260 2228 12288
rect 1894 12257 1906 12260
rect 1848 12251 1906 12257
rect 2222 12248 2228 12260
rect 2280 12288 2286 12300
rect 2516 12288 2544 12316
rect 2280 12260 2544 12288
rect 2280 12248 2286 12260
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 3844 12260 4445 12288
rect 3844 12248 3850 12260
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 7340 12260 8125 12288
rect 7340 12248 7346 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 10051 12288 10079 12328
rect 10413 12325 10425 12328
rect 10459 12325 10471 12359
rect 10413 12319 10471 12325
rect 10502 12316 10508 12368
rect 10560 12316 10566 12368
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 11241 12359 11299 12365
rect 11241 12356 11253 12359
rect 11020 12328 11253 12356
rect 11020 12316 11026 12328
rect 11241 12325 11253 12328
rect 11287 12356 11299 12359
rect 11977 12359 12035 12365
rect 11977 12356 11989 12359
rect 11287 12328 11989 12356
rect 11287 12325 11299 12328
rect 11241 12319 11299 12325
rect 11977 12325 11989 12328
rect 12023 12325 12035 12359
rect 11977 12319 12035 12325
rect 9272 12260 10079 12288
rect 10321 12291 10379 12297
rect 9272 12248 9278 12260
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10520 12288 10548 12316
rect 10367 12260 10732 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 2682 12180 2688 12232
rect 2740 12220 2746 12232
rect 3697 12223 3755 12229
rect 3697 12220 3709 12223
rect 2740 12192 3709 12220
rect 2740 12180 2746 12192
rect 3697 12189 3709 12192
rect 3743 12220 3755 12223
rect 4522 12220 4528 12232
rect 3743 12192 4528 12220
rect 3743 12189 3755 12192
rect 3697 12183 3755 12189
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 3326 12112 3332 12164
rect 3384 12152 3390 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 3384 12124 4077 12152
rect 3384 12112 3390 12124
rect 4065 12121 4077 12124
rect 4111 12121 4123 12155
rect 4065 12115 4123 12121
rect 4724 12084 4752 12183
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4856 12192 4905 12220
rect 4856 12180 4862 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12220 7987 12223
rect 8018 12220 8024 12232
rect 7975 12192 8024 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 9907 12192 10609 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6822 12152 6828 12164
rect 6052 12124 6828 12152
rect 6052 12112 6058 12124
rect 6822 12112 6828 12124
rect 6880 12112 6886 12164
rect 9493 12155 9551 12161
rect 9493 12121 9505 12155
rect 9539 12152 9551 12155
rect 9539 12124 10180 12152
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 6270 12084 6276 12096
rect 4724 12056 6276 12084
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 7285 12087 7343 12093
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 8478 12084 8484 12096
rect 7331 12056 8484 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9766 12084 9772 12096
rect 9180 12056 9772 12084
rect 9180 12044 9186 12056
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 9953 12087 10011 12093
rect 9953 12053 9965 12087
rect 9999 12084 10011 12087
rect 10042 12084 10048 12096
rect 9999 12056 10048 12084
rect 9999 12053 10011 12056
rect 9953 12047 10011 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10152 12084 10180 12124
rect 10226 12084 10232 12096
rect 10152 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10704 12084 10732 12260
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 11149 12291 11207 12297
rect 11149 12288 11161 12291
rect 10928 12260 11161 12288
rect 10928 12248 10934 12260
rect 11149 12257 11161 12260
rect 11195 12288 11207 12291
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11195 12260 12173 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12360 12288 12388 12396
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 13722 12424 13728 12436
rect 12860 12396 13728 12424
rect 12860 12384 12866 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14001 12427 14059 12433
rect 14001 12424 14013 12427
rect 13872 12396 14013 12424
rect 13872 12384 13878 12396
rect 14001 12393 14013 12396
rect 14047 12393 14059 12427
rect 14001 12387 14059 12393
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 16390 12424 16396 12436
rect 14415 12396 16396 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16577 12427 16635 12433
rect 16577 12393 16589 12427
rect 16623 12424 16635 12427
rect 18049 12427 18107 12433
rect 18049 12424 18061 12427
rect 16623 12396 18061 12424
rect 16623 12393 16635 12396
rect 16577 12387 16635 12393
rect 18049 12393 18061 12396
rect 18095 12393 18107 12427
rect 18049 12387 18107 12393
rect 18414 12384 18420 12436
rect 18472 12424 18478 12436
rect 18509 12427 18567 12433
rect 18509 12424 18521 12427
rect 18472 12396 18521 12424
rect 18472 12384 18478 12396
rect 18509 12393 18521 12396
rect 18555 12393 18567 12427
rect 19334 12424 19340 12436
rect 19295 12396 19340 12424
rect 18509 12387 18567 12393
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 19702 12424 19708 12436
rect 19663 12396 19708 12424
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 20070 12384 20076 12436
rect 20128 12424 20134 12436
rect 20165 12427 20223 12433
rect 20165 12424 20177 12427
rect 20128 12396 20177 12424
rect 20128 12384 20134 12396
rect 20165 12393 20177 12396
rect 20211 12424 20223 12427
rect 20254 12424 20260 12436
rect 20211 12396 20260 12424
rect 20211 12393 20223 12396
rect 20165 12387 20223 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 14642 12356 14648 12368
rect 12697 12328 14648 12356
rect 12697 12288 12725 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 18748 12328 19932 12356
rect 18748 12316 18754 12328
rect 12802 12297 12808 12300
rect 12796 12288 12808 12297
rect 12360 12260 12725 12288
rect 12763 12260 12808 12288
rect 12161 12251 12219 12257
rect 12796 12251 12808 12260
rect 12802 12248 12808 12251
rect 12860 12248 12866 12300
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 13412 12260 14473 12288
rect 13412 12248 13418 12260
rect 14461 12257 14473 12260
rect 14507 12288 14519 12291
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14507 12260 14841 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 15654 12288 15660 12300
rect 15615 12260 15660 12288
rect 14829 12251 14887 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16206 12288 16212 12300
rect 15795 12260 16212 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 16942 12288 16948 12300
rect 16903 12260 16948 12288
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17954 12288 17960 12300
rect 17915 12260 17960 12288
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18877 12291 18935 12297
rect 18877 12288 18889 12291
rect 18104 12260 18889 12288
rect 18104 12248 18110 12260
rect 18877 12257 18889 12260
rect 18923 12257 18935 12291
rect 18877 12251 18935 12257
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12220 11483 12223
rect 12250 12220 12256 12232
rect 11471 12192 12256 12220
rect 11471 12189 11483 12192
rect 11425 12183 11483 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12492 12192 12541 12220
rect 12492 12180 12498 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 15470 12220 15476 12232
rect 14691 12192 15476 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 15470 12180 15476 12192
rect 15528 12220 15534 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15528 12192 15853 12220
rect 15528 12180 15534 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17267 12192 17448 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 10781 12155 10839 12161
rect 10781 12121 10793 12155
rect 10827 12152 10839 12155
rect 17052 12152 17080 12183
rect 10827 12124 12572 12152
rect 10827 12121 10839 12124
rect 10781 12115 10839 12121
rect 11609 12087 11667 12093
rect 11609 12084 11621 12087
rect 10704 12056 11621 12084
rect 11609 12053 11621 12056
rect 11655 12084 11667 12087
rect 11790 12084 11796 12096
rect 11655 12056 11796 12084
rect 11655 12053 11667 12056
rect 11609 12047 11667 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 12544 12084 12572 12124
rect 13556 12124 17080 12152
rect 13556 12084 13584 12124
rect 13906 12084 13912 12096
rect 12544 12056 13584 12084
rect 13819 12056 13912 12084
rect 13906 12044 13912 12056
rect 13964 12084 13970 12096
rect 14366 12084 14372 12096
rect 13964 12056 14372 12084
rect 13964 12044 13970 12056
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 14918 12044 14924 12096
rect 14976 12084 14982 12096
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 14976 12056 15025 12084
rect 14976 12044 14982 12056
rect 15013 12053 15025 12056
rect 15059 12053 15071 12087
rect 15013 12047 15071 12053
rect 15102 12044 15108 12096
rect 15160 12084 15166 12096
rect 15289 12087 15347 12093
rect 15289 12084 15301 12087
rect 15160 12056 15301 12084
rect 15160 12044 15166 12056
rect 15289 12053 15301 12056
rect 15335 12053 15347 12087
rect 16206 12084 16212 12096
rect 16167 12056 16212 12084
rect 15289 12047 15347 12053
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16390 12084 16396 12096
rect 16351 12056 16396 12084
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 17420 12084 17448 12192
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 17862 12220 17868 12232
rect 17552 12192 17868 12220
rect 17552 12180 17558 12192
rect 17862 12180 17868 12192
rect 17920 12220 17926 12232
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 17920 12192 18153 12220
rect 17920 12180 17926 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18966 12220 18972 12232
rect 18927 12192 18972 12220
rect 18141 12183 18199 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 19150 12220 19156 12232
rect 19111 12192 19156 12220
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 19904 12229 19932 12328
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 17589 12155 17647 12161
rect 17589 12121 17601 12155
rect 17635 12152 17647 12155
rect 19812 12152 19840 12183
rect 17635 12124 19840 12152
rect 17635 12121 17647 12124
rect 17589 12115 17647 12121
rect 19150 12084 19156 12096
rect 16816 12056 19156 12084
rect 16816 12044 16822 12056
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 1857 11883 1915 11889
rect 1857 11880 1869 11883
rect 1820 11852 1869 11880
rect 1820 11840 1826 11852
rect 1857 11849 1869 11852
rect 1903 11849 1915 11883
rect 1857 11843 1915 11849
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4120 11852 5396 11880
rect 4120 11840 4126 11852
rect 5258 11812 5264 11824
rect 5219 11784 5264 11812
rect 5258 11772 5264 11784
rect 5316 11772 5322 11824
rect 5368 11812 5396 11852
rect 6086 11840 6092 11892
rect 6144 11880 6150 11892
rect 8297 11883 8355 11889
rect 8297 11880 8309 11883
rect 6144 11852 8309 11880
rect 6144 11840 6150 11852
rect 8297 11849 8309 11852
rect 8343 11849 8355 11883
rect 8297 11843 8355 11849
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9493 11883 9551 11889
rect 9493 11880 9505 11883
rect 9272 11852 9505 11880
rect 9272 11840 9278 11852
rect 9493 11849 9505 11852
rect 9539 11849 9551 11883
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 9493 11843 9551 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 10008 11852 10272 11880
rect 10008 11840 10014 11852
rect 10042 11812 10048 11824
rect 5368 11784 10048 11812
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2409 11747 2467 11753
rect 2409 11744 2421 11747
rect 2280 11716 2421 11744
rect 2280 11704 2286 11716
rect 2409 11713 2421 11716
rect 2455 11744 2467 11747
rect 2498 11744 2504 11756
rect 2455 11716 2504 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11744 6055 11747
rect 6178 11744 6184 11756
rect 6043 11716 6184 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 6178 11704 6184 11716
rect 6236 11744 6242 11756
rect 8018 11744 8024 11756
rect 6236 11716 8024 11744
rect 6236 11704 6242 11716
rect 8018 11704 8024 11716
rect 8076 11744 8082 11756
rect 8938 11744 8944 11756
rect 8076 11716 8121 11744
rect 8404 11716 8800 11744
rect 8899 11716 8944 11744
rect 8076 11704 8082 11716
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 3881 11679 3939 11685
rect 3881 11676 3893 11679
rect 2188 11648 3893 11676
rect 2188 11636 2194 11648
rect 3881 11645 3893 11648
rect 3927 11676 3939 11679
rect 4522 11676 4528 11688
rect 3927 11648 4528 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 4908 11648 5825 11676
rect 4154 11617 4160 11620
rect 4148 11608 4160 11617
rect 4115 11580 4160 11608
rect 4148 11571 4160 11580
rect 4154 11568 4160 11571
rect 4212 11568 4218 11620
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2372 11512 2417 11540
rect 2372 11500 2378 11512
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4908 11540 4936 11648
rect 5813 11645 5825 11648
rect 5859 11676 5871 11679
rect 6273 11679 6331 11685
rect 6273 11676 6285 11679
rect 5859 11648 6285 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 6273 11645 6285 11648
rect 6319 11645 6331 11679
rect 6273 11639 6331 11645
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7466 11676 7472 11688
rect 7055 11648 7472 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8404 11676 8432 11716
rect 7883 11648 8432 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8536 11648 8677 11676
rect 8536 11636 8542 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8772 11676 8800 11716
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 10134 11744 10140 11756
rect 10095 11716 10140 11744
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10244 11753 10272 11852
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 11882 11880 11888 11892
rect 11112 11852 11888 11880
rect 11112 11840 11118 11852
rect 11882 11840 11888 11852
rect 11940 11880 11946 11892
rect 12894 11880 12900 11892
rect 11940 11852 12900 11880
rect 11940 11840 11946 11852
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 14090 11880 14096 11892
rect 13127 11852 14096 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 14240 11852 14657 11880
rect 14240 11840 14246 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 14918 11840 14924 11892
rect 14976 11880 14982 11892
rect 15654 11880 15660 11892
rect 14976 11852 15660 11880
rect 14976 11840 14982 11852
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16206 11840 16212 11892
rect 16264 11880 16270 11892
rect 17862 11880 17868 11892
rect 16264 11852 17448 11880
rect 17823 11852 17868 11880
rect 16264 11840 16270 11852
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 11790 11812 11796 11824
rect 11296 11784 11796 11812
rect 11296 11772 11302 11784
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 12250 11772 12256 11824
rect 12308 11812 12314 11824
rect 12986 11812 12992 11824
rect 12308 11784 12992 11812
rect 12308 11772 12314 11784
rect 12986 11772 12992 11784
rect 13044 11772 13050 11824
rect 14108 11812 14136 11840
rect 17420 11812 17448 11852
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18509 11883 18567 11889
rect 18509 11849 18521 11883
rect 18555 11880 18567 11883
rect 18598 11880 18604 11892
rect 18555 11852 18604 11880
rect 18555 11849 18567 11852
rect 18509 11843 18567 11849
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 21266 11880 21272 11892
rect 19392 11852 21272 11880
rect 19392 11840 19398 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 19702 11812 19708 11824
rect 14108 11784 15700 11812
rect 17420 11784 19708 11812
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 12066 11744 12072 11756
rect 12027 11716 12072 11744
rect 11149 11707 11207 11713
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 8772 11648 9137 11676
rect 8665 11639 8723 11645
rect 9125 11645 9137 11648
rect 9171 11676 9183 11679
rect 10778 11676 10784 11688
rect 9171 11648 10784 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 10778 11636 10784 11648
rect 10836 11676 10842 11688
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 10836 11648 10885 11676
rect 10836 11636 10842 11648
rect 10873 11645 10885 11648
rect 10919 11676 10931 11679
rect 10919 11648 11100 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 5721 11611 5779 11617
rect 5721 11577 5733 11611
rect 5767 11608 5779 11611
rect 6457 11611 6515 11617
rect 6457 11608 6469 11611
rect 5767 11580 6469 11608
rect 5767 11577 5779 11580
rect 5721 11571 5779 11577
rect 6457 11577 6469 11580
rect 6503 11608 6515 11611
rect 7190 11608 7196 11620
rect 6503 11580 7196 11608
rect 6503 11577 6515 11580
rect 6457 11571 6515 11577
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 7484 11580 8769 11608
rect 4396 11512 4936 11540
rect 4396 11500 4402 11512
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5132 11512 5365 11540
rect 5132 11500 5138 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 7484 11549 7512 11580
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 10965 11611 11023 11617
rect 10965 11608 10977 11611
rect 8757 11571 8815 11577
rect 9324 11580 10977 11608
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7469 11543 7527 11549
rect 7469 11509 7481 11543
rect 7515 11509 7527 11543
rect 7469 11503 7527 11509
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 9324 11549 9352 11580
rect 10965 11577 10977 11580
rect 11011 11577 11023 11611
rect 10965 11571 11023 11577
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7800 11512 7941 11540
rect 7800 11500 7806 11512
rect 7929 11509 7941 11512
rect 7975 11540 7987 11543
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 7975 11512 9321 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 9309 11503 9367 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10502 11540 10508 11552
rect 10463 11512 10508 11540
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 11072 11540 11100 11648
rect 11164 11608 11192 11707
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 12400 11716 13185 11744
rect 12400 11704 12406 11716
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 15102 11744 15108 11756
rect 15063 11716 15108 11744
rect 13173 11707 13231 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11676 11943 11679
rect 12434 11676 12440 11688
rect 11931 11648 12440 11676
rect 11931 11645 11943 11648
rect 11885 11639 11943 11645
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11676 12679 11679
rect 13081 11679 13139 11685
rect 13081 11676 13093 11679
rect 12667 11648 13093 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 13081 11645 13093 11648
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 13440 11679 13498 11685
rect 13440 11645 13452 11679
rect 13486 11676 13498 11679
rect 13906 11676 13912 11688
rect 13486 11648 13912 11676
rect 13486 11645 13498 11648
rect 13440 11639 13498 11645
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 14792 11648 15025 11676
rect 14792 11636 14798 11648
rect 15013 11645 15025 11648
rect 15059 11645 15071 11679
rect 15212 11676 15240 11707
rect 15672 11685 15700 11784
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 19794 11772 19800 11824
rect 19852 11812 19858 11824
rect 19852 11784 20024 11812
rect 19852 11772 19858 11784
rect 18598 11704 18604 11756
rect 18656 11744 18662 11756
rect 18782 11744 18788 11756
rect 18656 11716 18788 11744
rect 18656 11704 18662 11716
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 19150 11744 19156 11756
rect 19111 11716 19156 11744
rect 19150 11704 19156 11716
rect 19208 11704 19214 11756
rect 19886 11744 19892 11756
rect 19847 11716 19892 11744
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 19996 11744 20024 11784
rect 20625 11747 20683 11753
rect 19996 11716 20392 11744
rect 15013 11639 15071 11645
rect 15120 11648 15240 11676
rect 15657 11679 15715 11685
rect 11238 11608 11244 11620
rect 11151 11580 11244 11608
rect 11238 11568 11244 11580
rect 11296 11608 11302 11620
rect 11296 11580 13676 11608
rect 11296 11568 11302 11580
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 11072 11512 11345 11540
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 11514 11540 11520 11552
rect 11475 11512 11520 11540
rect 11333 11503 11391 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 11977 11543 12035 11549
rect 11977 11509 11989 11543
rect 12023 11540 12035 11543
rect 12158 11540 12164 11552
rect 12023 11512 12164 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 12437 11543 12495 11549
rect 12437 11540 12449 11543
rect 12400 11512 12449 11540
rect 12400 11500 12406 11512
rect 12437 11509 12449 11512
rect 12483 11509 12495 11543
rect 13648 11540 13676 11580
rect 13722 11568 13728 11620
rect 13780 11608 13786 11620
rect 15120 11608 15148 11648
rect 15657 11645 15669 11679
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 16485 11679 16543 11685
rect 16485 11645 16497 11679
rect 16531 11676 16543 11679
rect 16574 11676 16580 11688
rect 16531 11648 16580 11676
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 16758 11685 16764 11688
rect 16752 11676 16764 11685
rect 16719 11648 16764 11676
rect 16752 11639 16764 11648
rect 16758 11636 16764 11639
rect 16816 11636 16822 11688
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 20070 11676 20076 11688
rect 17368 11648 20076 11676
rect 17368 11636 17374 11648
rect 20070 11636 20076 11648
rect 20128 11676 20134 11688
rect 20364 11685 20392 11716
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 21542 11744 21548 11756
rect 20671 11716 21548 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 20349 11679 20407 11685
rect 20128 11648 20300 11676
rect 20128 11636 20134 11648
rect 13780 11580 15148 11608
rect 13780 11568 13786 11580
rect 17126 11568 17132 11620
rect 17184 11608 17190 11620
rect 19797 11611 19855 11617
rect 19797 11608 19809 11611
rect 17184 11580 19809 11608
rect 17184 11568 17190 11580
rect 19797 11577 19809 11580
rect 19843 11608 19855 11611
rect 20165 11611 20223 11617
rect 20165 11608 20177 11611
rect 19843 11580 20177 11608
rect 19843 11577 19855 11580
rect 19797 11571 19855 11577
rect 20165 11577 20177 11580
rect 20211 11577 20223 11611
rect 20272 11608 20300 11648
rect 20349 11645 20361 11679
rect 20395 11645 20407 11679
rect 21085 11679 21143 11685
rect 21085 11676 21097 11679
rect 20349 11639 20407 11645
rect 20456 11648 21097 11676
rect 20456 11608 20484 11648
rect 21085 11645 21097 11648
rect 21131 11645 21143 11679
rect 21085 11639 21143 11645
rect 20272 11580 20484 11608
rect 20165 11571 20223 11577
rect 20714 11568 20720 11620
rect 20772 11608 20778 11620
rect 20772 11580 21312 11608
rect 20772 11568 20778 11580
rect 21284 11552 21312 11580
rect 13814 11540 13820 11552
rect 13648 11512 13820 11540
rect 12437 11503 12495 11509
rect 13814 11500 13820 11512
rect 13872 11540 13878 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 13872 11512 14565 11540
rect 13872 11500 13878 11512
rect 14553 11509 14565 11512
rect 14599 11509 14611 11543
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 14553 11503 14611 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 18690 11540 18696 11552
rect 16448 11512 18696 11540
rect 16448 11500 16454 11512
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 18874 11540 18880 11552
rect 18835 11512 18880 11540
rect 18874 11500 18880 11512
rect 18932 11500 18938 11552
rect 18969 11543 19027 11549
rect 18969 11509 18981 11543
rect 19015 11540 19027 11543
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 19015 11512 19349 11540
rect 19015 11509 19027 11512
rect 18969 11503 19027 11509
rect 19337 11509 19349 11512
rect 19383 11509 19395 11543
rect 19702 11540 19708 11552
rect 19615 11512 19708 11540
rect 19337 11503 19395 11509
rect 19702 11500 19708 11512
rect 19760 11540 19766 11552
rect 20622 11540 20628 11552
rect 19760 11512 20628 11540
rect 19760 11500 19766 11512
rect 20622 11500 20628 11512
rect 20680 11540 20686 11552
rect 20901 11543 20959 11549
rect 20901 11540 20913 11543
rect 20680 11512 20913 11540
rect 20680 11500 20686 11512
rect 20901 11509 20913 11512
rect 20947 11509 20959 11543
rect 21266 11540 21272 11552
rect 21227 11512 21272 11540
rect 20901 11503 20959 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2556 11308 2973 11336
rect 2556 11296 2562 11308
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 2961 11299 3019 11305
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3786 11336 3792 11348
rect 3191 11308 3792 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4338 11336 4344 11348
rect 4120 11308 4344 11336
rect 4120 11296 4126 11308
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 4522 11336 4528 11348
rect 4483 11308 4528 11336
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 4801 11339 4859 11345
rect 4801 11305 4813 11339
rect 4847 11336 4859 11339
rect 4890 11336 4896 11348
rect 4847 11308 4896 11336
rect 4847 11305 4859 11308
rect 4801 11299 4859 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5132 11308 5181 11336
rect 5132 11296 5138 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 5169 11299 5227 11305
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 5307 11308 5641 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 5629 11299 5687 11305
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 7193 11339 7251 11345
rect 7193 11336 7205 11339
rect 6604 11308 7205 11336
rect 6604 11296 6610 11308
rect 7193 11305 7205 11308
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 7699 11308 8585 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9079 11308 9689 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 12158 11336 12164 11348
rect 12119 11308 12164 11336
rect 9677 11299 9735 11305
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12575 11308 13093 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13320 11308 13553 11336
rect 13320 11296 13326 11308
rect 13541 11305 13553 11308
rect 13587 11336 13599 11339
rect 13909 11339 13967 11345
rect 13909 11336 13921 11339
rect 13587 11308 13921 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 13909 11305 13921 11308
rect 13955 11305 13967 11339
rect 16942 11336 16948 11348
rect 16903 11308 16948 11336
rect 13909 11299 13967 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17773 11339 17831 11345
rect 17773 11336 17785 11339
rect 17135 11308 17785 11336
rect 2130 11268 2136 11280
rect 1780 11240 2136 11268
rect 1780 11200 1808 11240
rect 2130 11228 2136 11240
rect 2188 11228 2194 11280
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 6089 11271 6147 11277
rect 6089 11268 6101 11271
rect 5592 11240 6101 11268
rect 5592 11228 5598 11240
rect 6089 11237 6101 11240
rect 6135 11268 6147 11271
rect 6457 11271 6515 11277
rect 6457 11268 6469 11271
rect 6135 11240 6469 11268
rect 6135 11237 6147 11240
rect 6089 11231 6147 11237
rect 6457 11237 6469 11240
rect 6503 11237 6515 11271
rect 6457 11231 6515 11237
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 8389 11271 8447 11277
rect 8389 11268 8401 11271
rect 7800 11240 8401 11268
rect 7800 11228 7806 11240
rect 8389 11237 8401 11240
rect 8435 11237 8447 11271
rect 10134 11268 10140 11280
rect 10095 11240 10140 11268
rect 8389 11231 8447 11237
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 12621 11271 12679 11277
rect 12621 11268 12633 11271
rect 10560 11240 12633 11268
rect 10560 11228 10566 11240
rect 12621 11237 12633 11240
rect 12667 11237 12679 11271
rect 12621 11231 12679 11237
rect 12986 11228 12992 11280
rect 13044 11268 13050 11280
rect 15718 11271 15776 11277
rect 15718 11268 15730 11271
rect 13044 11240 15730 11268
rect 13044 11228 13050 11240
rect 15718 11237 15730 11240
rect 15764 11268 15776 11271
rect 17034 11268 17040 11280
rect 15764 11240 17040 11268
rect 15764 11237 15776 11240
rect 15718 11231 15776 11237
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 1688 11172 1808 11200
rect 1848 11203 1906 11209
rect 1578 11132 1584 11144
rect 1491 11104 1584 11132
rect 1578 11092 1584 11104
rect 1636 11132 1642 11144
rect 1688 11132 1716 11172
rect 1848 11169 1860 11203
rect 1894 11200 1906 11203
rect 2682 11200 2688 11212
rect 1894 11172 2688 11200
rect 1894 11169 1906 11172
rect 1848 11163 1906 11169
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 3513 11203 3571 11209
rect 3513 11169 3525 11203
rect 3559 11200 3571 11203
rect 4338 11200 4344 11212
rect 3559 11172 4344 11200
rect 3559 11169 3571 11172
rect 3513 11163 3571 11169
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11200 4767 11203
rect 4755 11172 5948 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 3602 11132 3608 11144
rect 1636 11104 1716 11132
rect 3563 11104 3608 11132
rect 1636 11092 1642 11104
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11132 3847 11135
rect 5258 11132 5264 11144
rect 3835 11104 5264 11132
rect 3835 11101 3847 11104
rect 3789 11095 3847 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5442 11132 5448 11144
rect 5403 11104 5448 11132
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5920 11064 5948 11172
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6052 11172 6097 11200
rect 6052 11160 6058 11172
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7432 11172 7573 11200
rect 7432 11160 7438 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 8938 11200 8944 11212
rect 8899 11172 8944 11200
rect 7561 11163 7619 11169
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9306 11160 9312 11212
rect 9364 11200 9370 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9364 11172 10057 11200
rect 9364 11160 9370 11172
rect 10045 11169 10057 11172
rect 10091 11200 10103 11203
rect 10778 11200 10784 11212
rect 10091 11172 10784 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 10956 11203 11014 11209
rect 10956 11169 10968 11203
rect 11002 11200 11014 11203
rect 11238 11200 11244 11212
rect 11002 11172 11244 11200
rect 11002 11169 11014 11172
rect 10956 11163 11014 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 13354 11200 13360 11212
rect 12636 11172 13360 11200
rect 6178 11132 6184 11144
rect 6139 11104 6184 11132
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 7156 11104 7757 11132
rect 7156 11092 7162 11104
rect 7745 11101 7757 11104
rect 7791 11132 7803 11135
rect 8202 11132 8208 11144
rect 7791 11104 8208 11132
rect 7791 11101 7803 11104
rect 7745 11095 7803 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 10134 11132 10140 11144
rect 9416 11104 10140 11132
rect 6730 11064 6736 11076
rect 4080 11036 4384 11064
rect 5920 11036 6736 11064
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 4080 10996 4108 11036
rect 4246 10996 4252 11008
rect 3844 10968 4108 10996
rect 4207 10968 4252 10996
rect 3844 10956 3850 10968
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 4356 10996 4384 11036
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 6822 11024 6828 11076
rect 6880 11064 6886 11076
rect 9416 11073 9444 11104
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10686 11132 10692 11144
rect 10284 11104 10329 11132
rect 10647 11104 10692 11132
rect 10284 11092 10290 11104
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 9401 11067 9459 11073
rect 9401 11064 9413 11067
rect 6880 11036 9413 11064
rect 6880 11024 6886 11036
rect 9401 11033 9413 11036
rect 9447 11033 9459 11067
rect 12636 11064 12664 11172
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11200 13507 11203
rect 13495 11172 13952 11200
rect 13495 11169 13507 11172
rect 13449 11163 13507 11169
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 13814 11132 13820 11144
rect 13771 11104 13820 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 9401 11027 9459 11033
rect 11900 11036 12664 11064
rect 8662 10996 8668 11008
rect 4356 10968 8668 10996
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 10042 10956 10048 11008
rect 10100 10996 10106 11008
rect 10597 10999 10655 11005
rect 10597 10996 10609 10999
rect 10100 10968 10609 10996
rect 10100 10956 10106 10968
rect 10597 10965 10609 10968
rect 10643 10996 10655 10999
rect 11900 10996 11928 11036
rect 12066 10996 12072 11008
rect 10643 10968 11928 10996
rect 12027 10968 12072 10996
rect 10643 10965 10655 10968
rect 10597 10959 10655 10965
rect 12066 10956 12072 10968
rect 12124 10996 12130 11008
rect 12820 10996 12848 11095
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 13924 11132 13952 11172
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 14550 11200 14556 11212
rect 14424 11172 14556 11200
rect 14424 11160 14430 11172
rect 14550 11160 14556 11172
rect 14608 11200 14614 11212
rect 17135 11200 17163 11308
rect 17773 11305 17785 11308
rect 17819 11336 17831 11339
rect 17862 11336 17868 11348
rect 17819 11308 17868 11336
rect 17819 11305 17831 11308
rect 17773 11299 17831 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 17957 11339 18015 11345
rect 17957 11305 17969 11339
rect 18003 11336 18015 11339
rect 18046 11336 18052 11348
rect 18003 11308 18052 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18233 11339 18291 11345
rect 18233 11305 18245 11339
rect 18279 11336 18291 11339
rect 18966 11336 18972 11348
rect 18279 11308 18972 11336
rect 18279 11305 18291 11308
rect 18233 11299 18291 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 19518 11336 19524 11348
rect 19431 11308 19524 11336
rect 19518 11296 19524 11308
rect 19576 11336 19582 11348
rect 20257 11339 20315 11345
rect 19576 11308 20024 11336
rect 19576 11296 19582 11308
rect 17405 11271 17463 11277
rect 17405 11237 17417 11271
rect 17451 11237 17463 11271
rect 17405 11231 17463 11237
rect 18708 11240 18920 11268
rect 14608 11172 17163 11200
rect 14608 11160 14614 11172
rect 17218 11160 17224 11212
rect 17276 11200 17282 11212
rect 17313 11203 17371 11209
rect 17313 11200 17325 11203
rect 17276 11172 17325 11200
rect 17276 11160 17282 11172
rect 17313 11169 17325 11172
rect 17359 11169 17371 11203
rect 17313 11163 17371 11169
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13924 11104 14197 11132
rect 14185 11101 14197 11104
rect 14231 11132 14243 11135
rect 15286 11132 15292 11144
rect 14231 11104 15292 11132
rect 14231 11101 14243 11104
rect 14185 11095 14243 11101
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 15470 11132 15476 11144
rect 15383 11104 15476 11132
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 17420 11132 17448 11231
rect 18708 11209 18736 11240
rect 18601 11203 18659 11209
rect 18601 11169 18613 11203
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11169 18751 11203
rect 18892 11200 18920 11240
rect 19058 11228 19064 11280
rect 19116 11268 19122 11280
rect 19794 11268 19800 11280
rect 19116 11240 19800 11268
rect 19116 11228 19122 11240
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 18966 11200 18972 11212
rect 18892 11172 18972 11200
rect 18693 11163 18751 11169
rect 16816 11104 17448 11132
rect 16816 11092 16822 11104
rect 17586 11092 17592 11144
rect 17644 11132 17650 11144
rect 17644 11104 17689 11132
rect 17644 11092 17650 11104
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 18616 11132 18644 11163
rect 18966 11160 18972 11172
rect 19024 11200 19030 11212
rect 19334 11200 19340 11212
rect 19024 11172 19340 11200
rect 19024 11160 19030 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 19996 11200 20024 11308
rect 20257 11305 20269 11339
rect 20303 11336 20315 11339
rect 20714 11336 20720 11348
rect 20303 11308 20720 11336
rect 20303 11305 20315 11308
rect 20257 11299 20315 11305
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 21358 11336 21364 11348
rect 21131 11308 21364 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 20070 11228 20076 11280
rect 20128 11268 20134 11280
rect 20349 11271 20407 11277
rect 20349 11268 20361 11271
rect 20128 11240 20361 11268
rect 20128 11228 20134 11240
rect 20349 11237 20361 11240
rect 20395 11237 20407 11271
rect 21269 11271 21327 11277
rect 21269 11268 21281 11271
rect 20349 11231 20407 11237
rect 20456 11240 21281 11268
rect 20456 11200 20484 11240
rect 21269 11237 21281 11240
rect 21315 11237 21327 11271
rect 21269 11231 21327 11237
rect 19484 11172 19529 11200
rect 19996 11172 20484 11200
rect 19484 11160 19490 11172
rect 20530 11160 20536 11212
rect 20588 11200 20594 11212
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20588 11172 20913 11200
rect 20588 11160 20594 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 17920 11104 18644 11132
rect 18708 11104 18889 11132
rect 17920 11092 17926 11104
rect 12124 10968 12848 10996
rect 15488 10996 15516 11092
rect 16850 11064 16856 11076
rect 16811 11036 16856 11064
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 18708 11064 18736 11104
rect 18877 11101 18889 11104
rect 18923 11132 18935 11135
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 18923 11104 19625 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 19613 11101 19625 11104
rect 19659 11132 19671 11135
rect 19886 11132 19892 11144
rect 19659 11104 19892 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 19886 11092 19892 11104
rect 19944 11132 19950 11144
rect 20438 11132 20444 11144
rect 19944 11104 20444 11132
rect 19944 11092 19950 11104
rect 20438 11092 20444 11104
rect 20496 11092 20502 11144
rect 21453 11067 21511 11073
rect 21453 11064 21465 11067
rect 18607 11036 18736 11064
rect 18800 11036 19380 11064
rect 16574 10996 16580 11008
rect 15488 10968 16580 10996
rect 12124 10956 12130 10968
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 17586 10996 17592 11008
rect 17092 10968 17592 10996
rect 17092 10956 17098 10968
rect 17586 10956 17592 10968
rect 17644 10996 17650 11008
rect 18607 10996 18635 11036
rect 17644 10968 18635 10996
rect 17644 10956 17650 10968
rect 18690 10956 18696 11008
rect 18748 10996 18754 11008
rect 18800 10996 18828 11036
rect 19058 10996 19064 11008
rect 18748 10968 18828 10996
rect 19019 10968 19064 10996
rect 18748 10956 18754 10968
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 19352 10996 19380 11036
rect 19720 11036 21465 11064
rect 19426 10996 19432 11008
rect 19352 10968 19432 10996
rect 19426 10956 19432 10968
rect 19484 10996 19490 11008
rect 19720 10996 19748 11036
rect 21453 11033 21465 11036
rect 21499 11033 21511 11067
rect 21453 11027 21511 11033
rect 19886 10996 19892 11008
rect 19484 10968 19748 10996
rect 19847 10968 19892 10996
rect 19484 10956 19490 10968
rect 19886 10956 19892 10968
rect 19944 10956 19950 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2041 10795 2099 10801
rect 2041 10761 2053 10795
rect 2087 10792 2099 10795
rect 2314 10792 2320 10804
rect 2087 10764 2320 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 3513 10795 3571 10801
rect 3513 10761 3525 10795
rect 3559 10792 3571 10795
rect 3602 10792 3608 10804
rect 3559 10764 3608 10792
rect 3559 10761 3571 10764
rect 3513 10755 3571 10761
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4396 10764 5181 10792
rect 4396 10752 4402 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 6917 10795 6975 10801
rect 6917 10792 6929 10795
rect 5408 10764 6929 10792
rect 5408 10752 5414 10764
rect 6917 10761 6929 10764
rect 6963 10792 6975 10795
rect 7006 10792 7012 10804
rect 6963 10764 7012 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 8260 10764 8677 10792
rect 8260 10752 8266 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 8665 10755 8723 10761
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9401 10795 9459 10801
rect 9401 10792 9413 10795
rect 8996 10764 9413 10792
rect 8996 10752 9002 10764
rect 9401 10761 9413 10764
rect 9447 10761 9459 10795
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 9401 10755 9459 10761
rect 9876 10764 10517 10792
rect 4154 10724 4160 10736
rect 4067 10696 4160 10724
rect 2682 10656 2688 10668
rect 2643 10628 2688 10656
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 4080 10665 4108 10696
rect 4154 10684 4160 10696
rect 4212 10724 4218 10736
rect 9306 10724 9312 10736
rect 4212 10696 5488 10724
rect 9267 10696 9312 10724
rect 4212 10684 4218 10696
rect 5460 10668 5488 10696
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4396 10628 4813 10656
rect 4396 10616 4402 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5074 10656 5080 10668
rect 5031 10628 5080 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 9876 10665 9904 10764
rect 10505 10761 10517 10764
rect 10551 10792 10563 10795
rect 11054 10792 11060 10804
rect 10551 10764 11060 10792
rect 10551 10761 10563 10764
rect 10505 10755 10563 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11790 10752 11796 10804
rect 11848 10752 11854 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12492 10764 12537 10792
rect 12636 10764 17540 10792
rect 12492 10752 12498 10764
rect 11808 10724 11836 10752
rect 12636 10724 12664 10764
rect 11808 10696 12664 10724
rect 12894 10684 12900 10736
rect 12952 10724 12958 10736
rect 16758 10724 16764 10736
rect 12952 10696 16764 10724
rect 12952 10684 12958 10696
rect 16758 10684 16764 10696
rect 16816 10684 16822 10736
rect 17512 10724 17540 10764
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18601 10795 18659 10801
rect 18601 10792 18613 10795
rect 18012 10764 18613 10792
rect 18012 10752 18018 10764
rect 18601 10761 18613 10764
rect 18647 10761 18659 10795
rect 18601 10755 18659 10761
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 20441 10795 20499 10801
rect 20441 10792 20453 10795
rect 18932 10764 20453 10792
rect 18932 10752 18938 10764
rect 20441 10761 20453 10764
rect 20487 10761 20499 10795
rect 21450 10792 21456 10804
rect 21411 10764 21456 10792
rect 20441 10755 20499 10761
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 18046 10724 18052 10736
rect 17512 10696 18052 10724
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 19260 10696 19380 10724
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5500 10628 5733 10656
rect 5500 10616 5506 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 10042 10656 10048 10668
rect 9955 10628 10048 10656
rect 9861 10619 9919 10625
rect 10042 10616 10048 10628
rect 10100 10656 10106 10668
rect 10226 10656 10232 10668
rect 10100 10628 10232 10656
rect 10100 10616 10106 10628
rect 10226 10616 10232 10628
rect 10284 10616 10290 10668
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10744 10628 10885 10656
rect 10744 10616 10750 10628
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 10873 10619 10931 10625
rect 12636 10628 13001 10656
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 1995 10560 2513 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2501 10557 2513 10560
rect 2547 10588 2559 10591
rect 3326 10588 3332 10600
rect 2547 10560 3332 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 7282 10588 7288 10600
rect 6972 10560 7288 10588
rect 6972 10548 6978 10560
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7552 10591 7610 10597
rect 7552 10557 7564 10591
rect 7598 10588 7610 10591
rect 9214 10588 9220 10600
rect 7598 10560 9220 10588
rect 7598 10557 7610 10560
rect 7552 10551 7610 10557
rect 8220 10532 8248 10560
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 11140 10591 11198 10597
rect 11140 10557 11152 10591
rect 11186 10588 11198 10591
rect 12066 10588 12072 10600
rect 11186 10560 12072 10588
rect 11186 10557 11198 10560
rect 11140 10551 11198 10557
rect 12066 10548 12072 10560
rect 12124 10588 12130 10600
rect 12636 10588 12664 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14093 10659 14151 10665
rect 14093 10656 14105 10659
rect 13872 10628 14105 10656
rect 13872 10616 13878 10628
rect 14093 10625 14105 10628
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14182 10616 14188 10668
rect 14240 10656 14246 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 14240 10628 15393 10656
rect 14240 10616 14246 10628
rect 15381 10625 15393 10628
rect 15427 10625 15439 10659
rect 15562 10656 15568 10668
rect 15523 10628 15568 10656
rect 15381 10619 15439 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10656 16451 10659
rect 16666 10656 16672 10668
rect 16439 10628 16672 10656
rect 16439 10625 16451 10628
rect 16393 10619 16451 10625
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 17218 10616 17224 10668
rect 17276 10656 17282 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17276 10628 17877 10656
rect 17276 10616 17282 10628
rect 17865 10625 17877 10628
rect 17911 10656 17923 10659
rect 18138 10656 18144 10668
rect 17911 10628 18144 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 19058 10656 19064 10668
rect 19019 10628 19064 10656
rect 19058 10616 19064 10628
rect 19116 10616 19122 10668
rect 19260 10665 19288 10696
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10625 19303 10659
rect 19352 10656 19380 10696
rect 19702 10656 19708 10668
rect 19352 10628 19708 10656
rect 19245 10619 19303 10625
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 20162 10656 20168 10668
rect 20123 10628 20168 10656
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 20438 10616 20444 10668
rect 20496 10656 20502 10668
rect 20993 10659 21051 10665
rect 20993 10656 21005 10659
rect 20496 10628 21005 10656
rect 20496 10616 20502 10628
rect 20993 10625 21005 10628
rect 21039 10625 21051 10659
rect 20993 10619 21051 10625
rect 12124 10560 12664 10588
rect 12124 10548 12130 10560
rect 13170 10548 13176 10600
rect 13228 10588 13234 10600
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13228 10560 13921 10588
rect 13228 10548 13234 10560
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 15746 10548 15752 10600
rect 15804 10588 15810 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15804 10560 16129 10588
rect 15804 10548 15810 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 18012 10560 18061 10588
rect 18012 10548 18018 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19886 10588 19892 10600
rect 19015 10560 19892 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19886 10548 19892 10560
rect 19944 10548 19950 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 20806 10588 20812 10600
rect 20027 10560 20812 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 21266 10588 21272 10600
rect 21227 10560 21272 10588
rect 21266 10548 21272 10560
rect 21324 10548 21330 10600
rect 3881 10523 3939 10529
rect 3881 10489 3893 10523
rect 3927 10520 3939 10523
rect 3927 10492 4384 10520
rect 3927 10489 3939 10492
rect 3881 10483 3939 10489
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 1811 10424 2421 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 2409 10421 2421 10424
rect 2455 10452 2467 10455
rect 2498 10452 2504 10464
rect 2455 10424 2504 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 2866 10452 2872 10464
rect 2827 10424 2872 10452
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 3970 10452 3976 10464
rect 3931 10424 3976 10452
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4356 10461 4384 10492
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 6178 10520 6184 10532
rect 5132 10492 6184 10520
rect 5132 10480 5138 10492
rect 6178 10480 6184 10492
rect 6236 10480 6242 10532
rect 8202 10480 8208 10532
rect 8260 10480 8266 10532
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13265 10523 13323 10529
rect 13265 10520 13277 10523
rect 12851 10492 13277 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13265 10489 13277 10492
rect 13311 10489 13323 10523
rect 16209 10523 16267 10529
rect 16209 10520 16221 10523
rect 13265 10483 13323 10489
rect 14936 10492 16221 10520
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10421 4399 10455
rect 4341 10415 4399 10421
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 5166 10452 5172 10464
rect 4755 10424 5172 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 5718 10452 5724 10464
rect 5675 10424 5724 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5994 10452 6000 10464
rect 5955 10424 6000 10452
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 9769 10455 9827 10461
rect 9769 10421 9781 10455
rect 9815 10452 9827 10455
rect 9858 10452 9864 10464
rect 9815 10424 9864 10452
rect 9815 10421 9827 10424
rect 9769 10415 9827 10421
rect 9858 10412 9864 10424
rect 9916 10452 9922 10464
rect 10226 10452 10232 10464
rect 9916 10424 10232 10452
rect 9916 10412 9922 10424
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11790 10452 11796 10464
rect 10560 10424 11796 10452
rect 10560 10412 10566 10424
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 12216 10424 12265 10452
rect 12216 10412 12222 10424
rect 12253 10421 12265 10424
rect 12299 10421 12311 10455
rect 12253 10415 12311 10421
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13541 10455 13599 10461
rect 13541 10452 13553 10455
rect 12943 10424 13553 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13541 10421 13553 10424
rect 13587 10421 13599 10455
rect 13541 10415 13599 10421
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 14047 10424 14473 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14461 10421 14473 10424
rect 14507 10452 14519 10455
rect 14734 10452 14740 10464
rect 14507 10424 14740 10452
rect 14507 10421 14519 10424
rect 14461 10415 14519 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 14936 10461 14964 10492
rect 16209 10489 16221 10492
rect 16255 10489 16267 10523
rect 20254 10520 20260 10532
rect 16209 10483 16267 10489
rect 16684 10492 20260 10520
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10421 14979 10455
rect 14921 10415 14979 10421
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15654 10452 15660 10464
rect 15335 10424 15660 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 15749 10455 15807 10461
rect 15749 10421 15761 10455
rect 15795 10452 15807 10455
rect 16684 10452 16712 10492
rect 20254 10480 20260 10492
rect 20312 10480 20318 10532
rect 15795 10424 16712 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 18966 10452 18972 10464
rect 17828 10424 18972 10452
rect 17828 10412 17834 10424
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19426 10452 19432 10464
rect 19116 10424 19432 10452
rect 19116 10412 19122 10424
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 19610 10452 19616 10464
rect 19571 10424 19616 10452
rect 19610 10412 19616 10424
rect 19668 10412 19674 10464
rect 20070 10452 20076 10464
rect 20031 10424 20076 10452
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 20714 10452 20720 10464
rect 20404 10424 20720 10452
rect 20404 10412 20410 10424
rect 20714 10412 20720 10424
rect 20772 10452 20778 10464
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 20772 10424 20821 10452
rect 20772 10412 20778 10424
rect 20809 10421 20821 10424
rect 20855 10421 20867 10455
rect 20809 10415 20867 10421
rect 20898 10412 20904 10464
rect 20956 10452 20962 10464
rect 20956 10424 21001 10452
rect 20956 10412 20962 10424
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2222 10248 2228 10260
rect 2087 10220 2228 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 2866 10248 2872 10260
rect 2455 10220 2872 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 3016 10220 3065 10248
rect 3016 10208 3022 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 3053 10211 3111 10217
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 4028 10220 4537 10248
rect 4028 10208 4034 10220
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 4525 10211 4583 10217
rect 4985 10251 5043 10257
rect 4985 10217 4997 10251
rect 5031 10248 5043 10251
rect 5350 10248 5356 10260
rect 5031 10220 5356 10248
rect 5031 10217 5043 10220
rect 4985 10211 5043 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 5500 10220 6929 10248
rect 5500 10208 5506 10220
rect 6917 10217 6929 10220
rect 6963 10248 6975 10251
rect 8846 10248 8852 10260
rect 6963 10220 8852 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9214 10248 9220 10260
rect 9175 10220 9220 10248
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 10318 10248 10324 10260
rect 10275 10220 10324 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 10551 10220 13001 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 12989 10211 13047 10217
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 13228 10220 13369 10248
rect 13228 10208 13234 10220
rect 13357 10217 13369 10220
rect 13403 10217 13415 10251
rect 13357 10211 13415 10217
rect 14369 10251 14427 10257
rect 14369 10217 14381 10251
rect 14415 10248 14427 10251
rect 14550 10248 14556 10260
rect 14415 10220 14556 10248
rect 14415 10217 14427 10220
rect 14369 10211 14427 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 14737 10251 14795 10257
rect 14737 10217 14749 10251
rect 14783 10248 14795 10251
rect 16206 10248 16212 10260
rect 14783 10220 16212 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16666 10248 16672 10260
rect 16627 10220 16672 10248
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17586 10208 17592 10260
rect 17644 10248 17650 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 17644 10220 18153 10248
rect 17644 10208 17650 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 18969 10251 19027 10257
rect 18969 10217 18981 10251
rect 19015 10248 19027 10251
rect 19337 10251 19395 10257
rect 19337 10248 19349 10251
rect 19015 10220 19349 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 19337 10217 19349 10220
rect 19383 10217 19395 10251
rect 19337 10211 19395 10217
rect 2498 10140 2504 10192
rect 2556 10180 2562 10192
rect 3605 10183 3663 10189
rect 3605 10180 3617 10183
rect 2556 10152 3617 10180
rect 2556 10140 2562 10152
rect 3605 10149 3617 10152
rect 3651 10149 3663 10183
rect 4154 10180 4160 10192
rect 4115 10152 4160 10180
rect 3605 10143 3663 10149
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2866 10112 2872 10124
rect 2827 10084 2872 10112
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3620 10112 3648 10143
rect 4154 10140 4160 10152
rect 4212 10140 4218 10192
rect 4249 10183 4307 10189
rect 4249 10149 4261 10183
rect 4295 10180 4307 10183
rect 5534 10180 5540 10192
rect 4295 10152 5540 10180
rect 4295 10149 4307 10152
rect 4249 10143 4307 10149
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 12434 10180 12440 10192
rect 5736 10152 12440 10180
rect 4798 10112 4804 10124
rect 3620 10084 4804 10112
rect 4798 10072 4804 10084
rect 4856 10112 4862 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4856 10084 4905 10112
rect 4856 10072 4862 10084
rect 4893 10081 4905 10084
rect 4939 10081 4951 10115
rect 5736 10112 5764 10152
rect 12434 10140 12440 10152
rect 12492 10140 12498 10192
rect 15562 10189 15568 10192
rect 15556 10180 15568 10189
rect 15028 10152 15568 10180
rect 4893 10075 4951 10081
rect 5184 10084 5764 10112
rect 5804 10115 5862 10121
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 2501 10047 2559 10053
rect 2501 10044 2513 10047
rect 1627 10016 2513 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 2501 10013 2513 10016
rect 2547 10013 2559 10047
rect 2501 10007 2559 10013
rect 2516 9976 2544 10007
rect 2590 10004 2596 10056
rect 2648 10044 2654 10056
rect 4154 10044 4160 10056
rect 2648 10016 2693 10044
rect 3896 10016 4160 10044
rect 2648 10004 2654 10016
rect 3896 9976 3924 10016
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 5074 10044 5080 10056
rect 5035 10016 5080 10044
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 2516 9948 3924 9976
rect 3970 9936 3976 9988
rect 4028 9976 4034 9988
rect 5184 9976 5212 10084
rect 5804 10081 5816 10115
rect 5850 10112 5862 10115
rect 6178 10112 6184 10124
rect 5850 10084 6184 10112
rect 5850 10081 5862 10084
rect 5804 10075 5862 10081
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7558 10112 7564 10124
rect 7423 10084 7564 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 8093 10115 8151 10121
rect 8093 10112 8105 10115
rect 7668 10084 8105 10112
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 4028 9948 5212 9976
rect 4028 9936 4034 9948
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9908 1915 9911
rect 2682 9908 2688 9920
rect 1903 9880 2688 9908
rect 1903 9877 1915 9880
rect 1857 9871 1915 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3292 9880 3801 9908
rect 3292 9868 3298 9880
rect 3789 9877 3801 9880
rect 3835 9908 3847 9911
rect 5353 9911 5411 9917
rect 5353 9908 5365 9911
rect 3835 9880 5365 9908
rect 3835 9877 3847 9880
rect 3789 9871 3847 9877
rect 5353 9877 5365 9880
rect 5399 9877 5411 9911
rect 5552 9908 5580 10007
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7668 10053 7696 10084
rect 8093 10081 8105 10084
rect 8139 10112 8151 10115
rect 10042 10112 10048 10124
rect 8139 10084 10048 10112
rect 8139 10081 8151 10084
rect 8093 10075 8151 10081
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10112 10471 10115
rect 10594 10112 10600 10124
rect 10459 10084 10600 10112
rect 10459 10081 10471 10084
rect 10413 10075 10471 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 10870 10112 10876 10124
rect 10831 10084 10876 10112
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 12894 10112 12900 10124
rect 12855 10084 12900 10112
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 14366 10112 14372 10124
rect 13096 10084 14372 10112
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 7064 10016 7481 10044
rect 7064 10004 7070 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 10502 10044 10508 10056
rect 7837 10007 7895 10013
rect 8864 10016 10508 10044
rect 6638 9936 6644 9988
rect 6696 9976 6702 9988
rect 6696 9948 7236 9976
rect 6696 9936 6702 9948
rect 6914 9908 6920 9920
rect 5552 9880 6920 9908
rect 5353 9871 5411 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7208 9908 7236 9948
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 7742 9976 7748 9988
rect 7340 9948 7748 9976
rect 7340 9936 7346 9948
rect 7742 9936 7748 9948
rect 7800 9976 7806 9988
rect 7852 9976 7880 10007
rect 7800 9948 7880 9976
rect 7800 9936 7806 9948
rect 8864 9908 8892 10016
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 10612 10044 10640 10072
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10612 10016 10977 10044
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 11146 10044 11152 10056
rect 11107 10016 11152 10044
rect 10965 10007 11023 10013
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 13096 10044 13124 10084
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 12452 10016 13124 10044
rect 13173 10047 13231 10053
rect 9122 9936 9128 9988
rect 9180 9976 9186 9988
rect 12452 9976 12480 10016
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13814 10044 13820 10056
rect 13219 10016 13820 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 15028 10053 15056 10152
rect 15556 10143 15568 10152
rect 15562 10140 15568 10143
rect 15620 10140 15626 10192
rect 16684 10180 16712 10208
rect 17006 10183 17064 10189
rect 17006 10180 17018 10183
rect 16684 10152 17018 10180
rect 17006 10149 17018 10152
rect 17052 10149 17064 10183
rect 17006 10143 17064 10149
rect 18877 10183 18935 10189
rect 18877 10149 18889 10183
rect 18923 10180 18935 10183
rect 19610 10180 19616 10192
rect 18923 10152 19616 10180
rect 18923 10149 18935 10152
rect 18877 10143 18935 10149
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 20530 10180 20536 10192
rect 20491 10152 20536 10180
rect 20530 10140 20536 10152
rect 20588 10140 20594 10192
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10112 15347 10115
rect 16574 10112 16580 10124
rect 15335 10084 16580 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 16574 10072 16580 10084
rect 16632 10112 16638 10124
rect 16761 10115 16819 10121
rect 16761 10112 16773 10115
rect 16632 10084 16773 10112
rect 16632 10072 16638 10084
rect 16761 10081 16773 10084
rect 16807 10112 16819 10115
rect 16850 10112 16856 10124
rect 16807 10084 16856 10112
rect 16807 10081 16819 10084
rect 16761 10075 16819 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 19518 10112 19524 10124
rect 19208 10084 19524 10112
rect 19208 10072 19214 10084
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 19702 10112 19708 10124
rect 19663 10084 19708 10112
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 20254 10112 20260 10124
rect 20215 10084 20260 10112
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 15013 10047 15071 10053
rect 15013 10013 15025 10047
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 9180 9948 12480 9976
rect 12529 9979 12587 9985
rect 9180 9936 9186 9948
rect 12529 9945 12541 9979
rect 12575 9976 12587 9979
rect 14182 9976 14188 9988
rect 12575 9948 14188 9976
rect 12575 9945 12587 9948
rect 12529 9939 12587 9945
rect 14182 9936 14188 9948
rect 14240 9936 14246 9988
rect 14844 9976 14872 10007
rect 18690 10004 18696 10056
rect 18748 10044 18754 10056
rect 19061 10047 19119 10053
rect 19061 10044 19073 10047
rect 18748 10016 19073 10044
rect 18748 10004 18754 10016
rect 19061 10013 19073 10016
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19392 10016 19809 10044
rect 19392 10004 19398 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20162 10044 20168 10056
rect 20027 10016 20168 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 20898 10004 20904 10056
rect 20956 10004 20962 10056
rect 15194 9976 15200 9988
rect 14844 9948 15200 9976
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 18874 9936 18880 9988
rect 18932 9976 18938 9988
rect 20916 9976 20944 10004
rect 21269 9979 21327 9985
rect 21269 9976 21281 9979
rect 18932 9948 21281 9976
rect 18932 9936 18938 9948
rect 21269 9945 21281 9948
rect 21315 9945 21327 9979
rect 21269 9939 21327 9945
rect 7064 9880 7109 9908
rect 7208 9880 8892 9908
rect 7064 9868 7070 9880
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 12250 9908 12256 9920
rect 9548 9880 12256 9908
rect 9548 9868 9554 9880
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13170 9908 13176 9920
rect 12492 9880 13176 9908
rect 12492 9868 12498 9880
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 18509 9911 18567 9917
rect 18509 9877 18521 9911
rect 18555 9908 18567 9911
rect 20898 9908 20904 9920
rect 18555 9880 20904 9908
rect 18555 9877 18567 9880
rect 18509 9871 18567 9877
rect 20898 9868 20904 9880
rect 20956 9868 20962 9920
rect 21542 9908 21548 9920
rect 21503 9880 21548 9908
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 5994 9704 6000 9716
rect 3200 9676 6000 9704
rect 3200 9664 3206 9676
rect 5994 9664 6000 9676
rect 6052 9704 6058 9716
rect 6546 9704 6552 9716
rect 6052 9676 6552 9704
rect 6052 9664 6058 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 15473 9707 15531 9713
rect 7208 9676 7512 9704
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9605 2099 9639
rect 2041 9599 2099 9605
rect 4249 9639 4307 9645
rect 4249 9605 4261 9639
rect 4295 9605 4307 9639
rect 4249 9599 4307 9605
rect 4617 9639 4675 9645
rect 4617 9605 4629 9639
rect 4663 9636 4675 9639
rect 5718 9636 5724 9648
rect 4663 9608 5724 9636
rect 4663 9605 4675 9608
rect 4617 9599 4675 9605
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 2056 9500 2084 9599
rect 2682 9568 2688 9580
rect 2643 9540 2688 9568
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9537 2927 9571
rect 4264 9568 4292 9599
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 7208 9636 7236 9676
rect 7374 9636 7380 9648
rect 6788 9608 7236 9636
rect 7335 9608 7380 9636
rect 6788 9596 6794 9608
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 7484 9636 7512 9676
rect 15473 9673 15485 9707
rect 15519 9704 15531 9707
rect 15519 9676 15553 9704
rect 15519 9673 15531 9676
rect 15473 9667 15531 9673
rect 12158 9636 12164 9648
rect 7484 9608 8708 9636
rect 5074 9568 5080 9580
rect 4264 9540 5080 9568
rect 2869 9531 2927 9537
rect 1535 9472 2084 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 2130 9460 2136 9512
rect 2188 9500 2194 9512
rect 2884 9500 2912 9531
rect 5074 9528 5080 9540
rect 5132 9568 5138 9580
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 5132 9540 5181 9568
rect 5132 9528 5138 9540
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7837 9571 7895 9577
rect 7837 9568 7849 9571
rect 7064 9540 7849 9568
rect 7064 9528 7070 9540
rect 7837 9537 7849 9540
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8202 9568 8208 9580
rect 8067 9540 8208 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 2188 9472 2912 9500
rect 2188 9460 2194 9472
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 8680 9509 8708 9608
rect 10980 9608 12164 9636
rect 8665 9503 8723 9509
rect 4120 9472 8340 9500
rect 4120 9460 4126 9472
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 2866 9432 2872 9444
rect 1811 9404 2872 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3142 9441 3148 9444
rect 3136 9395 3148 9441
rect 3200 9432 3206 9444
rect 3200 9404 3236 9432
rect 3142 9392 3148 9395
rect 3200 9392 3206 9404
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 4985 9435 5043 9441
rect 4985 9432 4997 9435
rect 4212 9404 4997 9432
rect 4212 9392 4218 9404
rect 4985 9401 4997 9404
rect 5031 9401 5043 9435
rect 6917 9435 6975 9441
rect 6917 9432 6929 9435
rect 4985 9395 5043 9401
rect 5092 9404 6929 9432
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 2004 9336 2421 9364
rect 2004 9324 2010 9336
rect 2409 9333 2421 9336
rect 2455 9333 2467 9367
rect 2409 9327 2467 9333
rect 2501 9367 2559 9373
rect 2501 9333 2513 9367
rect 2547 9364 2559 9367
rect 2774 9364 2780 9376
rect 2547 9336 2780 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 5092 9373 5120 9404
rect 6917 9401 6929 9404
rect 6963 9432 6975 9435
rect 7558 9432 7564 9444
rect 6963 9404 7564 9432
rect 6963 9401 6975 9404
rect 6917 9395 6975 9401
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 7745 9435 7803 9441
rect 7745 9401 7757 9435
rect 7791 9432 7803 9435
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 7791 9404 8217 9432
rect 7791 9401 7803 9404
rect 7745 9395 7803 9401
rect 8205 9401 8217 9404
rect 8251 9401 8263 9435
rect 8312 9432 8340 9472
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9907 9472 9965 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 9953 9469 9965 9472
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 10220 9503 10278 9509
rect 10220 9469 10232 9503
rect 10266 9500 10278 9503
rect 10980 9500 11008 9608
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 15488 9636 15516 9667
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 18046 9704 18052 9716
rect 15896 9676 18052 9704
rect 15896 9664 15902 9676
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 20070 9704 20076 9716
rect 20031 9676 20076 9704
rect 20070 9664 20076 9676
rect 20128 9664 20134 9716
rect 15654 9636 15660 9648
rect 15488 9608 15660 9636
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 16206 9596 16212 9648
rect 16264 9636 16270 9648
rect 16301 9639 16359 9645
rect 16301 9636 16313 9639
rect 16264 9608 16313 9636
rect 16264 9596 16270 9608
rect 16301 9605 16313 9608
rect 16347 9605 16359 9639
rect 19426 9636 19432 9648
rect 19339 9608 19432 9636
rect 16301 9599 16359 9605
rect 19426 9596 19432 9608
rect 19484 9636 19490 9648
rect 20162 9636 20168 9648
rect 19484 9608 20168 9636
rect 19484 9596 19490 9608
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 15746 9568 15752 9580
rect 15528 9540 15752 9568
rect 15528 9528 15534 9540
rect 15746 9528 15752 9540
rect 15804 9568 15810 9580
rect 15933 9571 15991 9577
rect 15933 9568 15945 9571
rect 15804 9540 15945 9568
rect 15804 9528 15810 9540
rect 15933 9537 15945 9540
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9537 16175 9571
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16117 9531 16175 9537
rect 16408 9540 16865 9568
rect 10266 9472 11008 9500
rect 10266 9469 10278 9472
rect 10220 9463 10278 9469
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 12492 9472 13921 9500
rect 12492 9460 12498 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 14176 9503 14234 9509
rect 14176 9469 14188 9503
rect 14222 9500 14234 9503
rect 15838 9500 15844 9512
rect 14222 9472 15844 9500
rect 14222 9469 14234 9472
rect 14176 9463 14234 9469
rect 11054 9432 11060 9444
rect 8312 9404 11060 9432
rect 8205 9395 8263 9401
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 11146 9392 11152 9444
rect 11204 9432 11210 9444
rect 12250 9432 12256 9444
rect 11204 9404 12256 9432
rect 11204 9392 11210 9404
rect 12250 9392 12256 9404
rect 12308 9432 12314 9444
rect 12682 9435 12740 9441
rect 12682 9432 12694 9435
rect 12308 9404 12694 9432
rect 12308 9392 12314 9404
rect 12682 9401 12694 9404
rect 12728 9401 12740 9435
rect 12682 9395 12740 9401
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 3016 9336 4445 9364
rect 3016 9324 3022 9336
rect 4433 9333 4445 9336
rect 4479 9364 4491 9367
rect 5077 9367 5135 9373
rect 5077 9364 5089 9367
rect 4479 9336 5089 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 5077 9333 5089 9336
rect 5123 9333 5135 9367
rect 5077 9327 5135 9333
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8294 9364 8300 9376
rect 7708 9336 8300 9364
rect 7708 9324 7714 9336
rect 8294 9324 8300 9336
rect 8352 9364 8358 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 8352 9336 8493 9364
rect 8352 9324 8358 9336
rect 8481 9333 8493 9336
rect 8527 9364 8539 9367
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 8527 9336 9873 9364
rect 8527 9333 8539 9336
rect 8481 9327 8539 9333
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10962 9364 10968 9376
rect 10008 9336 10968 9364
rect 10008 9324 10014 9336
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11330 9364 11336 9376
rect 11291 9336 11336 9364
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 13814 9364 13820 9376
rect 13727 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9364 13878 9376
rect 14180 9364 14208 9463
rect 15838 9460 15844 9472
rect 15896 9500 15902 9512
rect 16132 9500 16160 9531
rect 16408 9500 16436 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 19852 9540 19901 9568
rect 19852 9528 19858 9540
rect 19889 9537 19901 9540
rect 19935 9537 19947 9571
rect 19889 9531 19947 9537
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9568 21235 9571
rect 21266 9568 21272 9580
rect 21223 9540 21272 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 15896 9472 16436 9500
rect 15896 9460 15902 9472
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 16540 9472 16773 9500
rect 16540 9460 16546 9472
rect 16761 9469 16773 9472
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17920 9472 18061 9500
rect 17920 9460 17926 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 20640 9500 20668 9531
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 20898 9500 20904 9512
rect 18049 9463 18107 9469
rect 18524 9472 20668 9500
rect 20859 9472 20904 9500
rect 18524 9444 18552 9472
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 14734 9392 14740 9444
rect 14792 9432 14798 9444
rect 16666 9432 16672 9444
rect 14792 9404 15792 9432
rect 16627 9404 16672 9432
rect 14792 9392 14798 9404
rect 15764 9376 15792 9404
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 18316 9435 18374 9441
rect 18316 9401 18328 9435
rect 18362 9432 18374 9435
rect 18506 9432 18512 9444
rect 18362 9404 18512 9432
rect 18362 9401 18374 9404
rect 18316 9395 18374 9401
rect 18506 9392 18512 9404
rect 18564 9392 18570 9444
rect 19794 9392 19800 9444
rect 19852 9432 19858 9444
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 19852 9404 20453 9432
rect 19852 9392 19858 9404
rect 20441 9401 20453 9404
rect 20487 9401 20499 9435
rect 20441 9395 20499 9401
rect 13872 9336 14208 9364
rect 15289 9367 15347 9373
rect 13872 9324 13878 9336
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15562 9364 15568 9376
rect 15335 9336 15568 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 15746 9324 15752 9376
rect 15804 9324 15810 9376
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 17126 9364 17132 9376
rect 15887 9336 17132 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 18966 9364 18972 9376
rect 18288 9336 18972 9364
rect 18288 9324 18294 9336
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 20533 9367 20591 9373
rect 20533 9333 20545 9367
rect 20579 9364 20591 9367
rect 20714 9364 20720 9376
rect 20579 9336 20720 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 20714 9324 20720 9336
rect 20772 9364 20778 9376
rect 21542 9364 21548 9376
rect 20772 9336 21548 9364
rect 20772 9324 20778 9336
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 3142 9160 3148 9172
rect 2740 9132 3148 9160
rect 2740 9120 2746 9132
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 7101 9163 7159 9169
rect 7101 9160 7113 9163
rect 6604 9132 7113 9160
rect 6604 9120 6610 9132
rect 7101 9129 7113 9132
rect 7147 9129 7159 9163
rect 7101 9123 7159 9129
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7653 9163 7711 9169
rect 7653 9160 7665 9163
rect 7239 9132 7665 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7653 9129 7665 9132
rect 7699 9160 7711 9163
rect 8386 9160 8392 9172
rect 7699 9132 8392 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8570 9160 8576 9172
rect 8527 9132 8576 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8570 9120 8576 9132
rect 8628 9160 8634 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8628 9132 9045 9160
rect 8628 9120 8634 9132
rect 9033 9129 9045 9132
rect 9079 9160 9091 9163
rect 9398 9160 9404 9172
rect 9079 9132 9404 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9539 9132 10241 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 10229 9129 10241 9132
rect 10275 9160 10287 9163
rect 10594 9160 10600 9172
rect 10275 9132 10600 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 10962 9160 10968 9172
rect 10923 9132 10968 9160
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11057 9163 11115 9169
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 11698 9160 11704 9172
rect 11103 9132 11704 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 12952 9132 13369 9160
rect 12952 9120 12958 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 13725 9163 13783 9169
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 14090 9160 14096 9172
rect 13771 9132 14096 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 14090 9120 14096 9132
rect 14148 9160 14154 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 14148 9132 14197 9160
rect 14148 9120 14154 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 15194 9120 15200 9172
rect 15252 9160 15258 9172
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 15252 9132 15301 9160
rect 15252 9120 15258 9132
rect 15289 9129 15301 9132
rect 15335 9129 15347 9163
rect 15746 9160 15752 9172
rect 15707 9132 15752 9160
rect 15289 9123 15347 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 16117 9163 16175 9169
rect 16117 9129 16129 9163
rect 16163 9160 16175 9163
rect 16574 9160 16580 9172
rect 16163 9132 16580 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 18230 9160 18236 9172
rect 16724 9132 18236 9160
rect 16724 9120 16730 9132
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 18506 9160 18512 9172
rect 18467 9132 18512 9160
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 19981 9163 20039 9169
rect 19981 9160 19993 9163
rect 18708 9132 19993 9160
rect 18708 9104 18736 9132
rect 19981 9129 19993 9132
rect 20027 9129 20039 9163
rect 20990 9160 20996 9172
rect 20951 9132 20996 9160
rect 19981 9123 20039 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 1118 9052 1124 9104
rect 1176 9092 1182 9104
rect 3326 9092 3332 9104
rect 1176 9064 3332 9092
rect 1176 9052 1182 9064
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 3510 9092 3516 9104
rect 3471 9064 3516 9092
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 6638 9092 6644 9104
rect 5132 9064 6644 9092
rect 5132 9052 5138 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 8312 9064 10640 9092
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 1854 9024 1860 9036
rect 1811 8996 1860 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 2032 9027 2090 9033
rect 2032 8993 2044 9027
rect 2078 9024 2090 9027
rect 2866 9024 2872 9036
rect 2078 8996 2872 9024
rect 2078 8993 2090 8996
rect 2032 8987 2090 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 9024 3295 9027
rect 4338 9024 4344 9036
rect 3283 8996 4344 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6822 9024 6828 9036
rect 6227 8996 6828 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 6178 8888 6184 8900
rect 3344 8860 6184 8888
rect 3344 8832 3372 8860
rect 6178 8848 6184 8860
rect 6236 8848 6242 8900
rect 6288 8888 6316 8919
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 7377 8959 7435 8965
rect 6420 8928 6465 8956
rect 6420 8916 6426 8928
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 8312 8956 8340 9064
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 9024 8447 9027
rect 9309 9027 9367 9033
rect 8435 8996 8984 9024
rect 8435 8993 8447 8996
rect 8389 8987 8447 8993
rect 8478 8956 8484 8968
rect 7423 8928 8484 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 8956 8965 8984 8996
rect 9309 8993 9321 9027
rect 9355 9024 9367 9027
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 9355 8996 10149 9024
rect 9355 8993 9367 8996
rect 9309 8987 9367 8993
rect 10137 8993 10149 8996
rect 10183 9024 10195 9027
rect 10318 9024 10324 9036
rect 10183 8996 10324 9024
rect 10183 8993 10195 8996
rect 10137 8987 10195 8993
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 8941 8959 8999 8965
rect 8628 8928 8673 8956
rect 8628 8916 8634 8928
rect 8941 8925 8953 8959
rect 8987 8956 8999 8959
rect 9950 8956 9956 8968
rect 8987 8928 9956 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 9858 8888 9864 8900
rect 6288 8860 9864 8888
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 10428 8888 10456 8919
rect 10612 8888 10640 9064
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 12152 9095 12210 9101
rect 10744 9064 11928 9092
rect 10744 9052 10750 9064
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 11900 9033 11928 9064
rect 12152 9061 12164 9095
rect 12198 9092 12210 9095
rect 18690 9092 18696 9104
rect 12198 9064 18696 9092
rect 12198 9061 12210 9064
rect 12152 9055 12210 9061
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 18868 9095 18926 9101
rect 18868 9061 18880 9095
rect 18914 9092 18926 9095
rect 19426 9092 19432 9104
rect 18914 9064 19432 9092
rect 18914 9061 18926 9064
rect 18868 9055 18926 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 11425 9027 11483 9033
rect 11425 9024 11437 9027
rect 11020 8996 11437 9024
rect 11020 8984 11026 8996
rect 11425 8993 11437 8996
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 12434 9024 12440 9036
rect 11931 8996 12440 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 12434 8984 12440 8996
rect 12492 8984 12498 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15028 8996 15669 9024
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11330 8956 11336 8968
rect 11195 8928 11336 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11164 8888 11192 8919
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13320 8928 13829 8956
rect 13320 8916 13326 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 13909 8959 13967 8965
rect 13909 8925 13921 8959
rect 13955 8925 13967 8959
rect 13909 8919 13967 8925
rect 13924 8888 13952 8919
rect 10428 8860 11192 8888
rect 13280 8860 13952 8888
rect 3326 8780 3332 8832
rect 3384 8780 3390 8832
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 4212 8792 4261 8820
rect 4212 8780 4218 8792
rect 4249 8789 4261 8792
rect 4295 8789 4307 8823
rect 4249 8783 4307 8789
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 4948 8792 5825 8820
rect 4948 8780 4954 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 6733 8823 6791 8829
rect 6733 8789 6745 8823
rect 6779 8820 6791 8823
rect 7282 8820 7288 8832
rect 6779 8792 7288 8820
rect 6779 8789 6791 8792
rect 6733 8783 6791 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8021 8823 8079 8829
rect 8021 8820 8033 8823
rect 7800 8792 8033 8820
rect 7800 8780 7806 8792
rect 8021 8789 8033 8792
rect 8067 8789 8079 8823
rect 9766 8820 9772 8832
rect 9727 8792 9772 8820
rect 8021 8783 8079 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 10284 8792 10609 8820
rect 10284 8780 10290 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 11698 8820 11704 8832
rect 11659 8792 11704 8820
rect 10597 8783 10655 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 13280 8829 13308 8860
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 12308 8792 13277 8820
rect 12308 8780 12314 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 15028 8829 15056 8996
rect 15657 8993 15669 8996
rect 15703 9024 15715 9027
rect 15930 9024 15936 9036
rect 15703 8996 15936 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16482 9024 16488 9036
rect 16443 8996 16488 9024
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 17402 9033 17408 9036
rect 17396 8987 17408 9033
rect 17460 9024 17466 9036
rect 17460 8996 17496 9024
rect 17402 8984 17408 8987
rect 17460 8984 17466 8996
rect 15838 8956 15844 8968
rect 15799 8928 15844 8956
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 18601 8959 18659 8965
rect 18601 8925 18613 8959
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 21174 8956 21180 8968
rect 20579 8928 21180 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 15746 8848 15752 8900
rect 15804 8888 15810 8900
rect 16669 8891 16727 8897
rect 16669 8888 16681 8891
rect 15804 8860 16681 8888
rect 15804 8848 15810 8860
rect 16669 8857 16681 8860
rect 16715 8888 16727 8891
rect 16758 8888 16764 8900
rect 16715 8860 16764 8888
rect 16715 8857 16727 8860
rect 16669 8851 16727 8857
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 14792 8792 15025 8820
rect 14792 8780 14798 8792
rect 15013 8789 15025 8792
rect 15059 8789 15071 8823
rect 15013 8783 15071 8789
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 17144 8820 17172 8919
rect 17862 8820 17868 8832
rect 17000 8792 17868 8820
rect 17000 8780 17006 8792
rect 17862 8780 17868 8792
rect 17920 8820 17926 8832
rect 18616 8820 18644 8919
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 20438 8848 20444 8900
rect 20496 8888 20502 8900
rect 20622 8888 20628 8900
rect 20496 8860 20628 8888
rect 20496 8848 20502 8860
rect 20622 8848 20628 8860
rect 20680 8888 20686 8900
rect 21085 8891 21143 8897
rect 21085 8888 21097 8891
rect 20680 8860 21097 8888
rect 20680 8848 20686 8860
rect 21085 8857 21097 8860
rect 21131 8857 21143 8891
rect 21085 8851 21143 8857
rect 18966 8820 18972 8832
rect 17920 8792 18972 8820
rect 17920 8780 17926 8792
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 20346 8780 20352 8832
rect 20404 8820 20410 8832
rect 21269 8823 21327 8829
rect 21269 8820 21281 8823
rect 20404 8792 21281 8820
rect 20404 8780 20410 8792
rect 21269 8789 21281 8792
rect 21315 8820 21327 8823
rect 21358 8820 21364 8832
rect 21315 8792 21364 8820
rect 21315 8789 21327 8792
rect 21269 8783 21327 8789
rect 21358 8780 21364 8792
rect 21416 8780 21422 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 2832 8588 2877 8616
rect 2832 8576 2838 8588
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 9858 8616 9864 8628
rect 4120 8588 9352 8616
rect 9819 8588 9864 8616
rect 4120 8576 4126 8588
rect 4338 8508 4344 8560
rect 4396 8548 4402 8560
rect 4433 8551 4491 8557
rect 4433 8548 4445 8551
rect 4396 8520 4445 8548
rect 4396 8508 4402 8520
rect 4433 8517 4445 8520
rect 4479 8517 4491 8551
rect 6822 8548 6828 8560
rect 6783 8520 6828 8548
rect 4433 8511 4491 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 7190 8508 7196 8560
rect 7248 8548 7254 8560
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 7248 8520 7665 8548
rect 7248 8508 7254 8520
rect 7653 8517 7665 8520
rect 7699 8517 7711 8551
rect 9324 8548 9352 8588
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 11238 8616 11244 8628
rect 10008 8588 11244 8616
rect 10008 8576 10014 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 12066 8616 12072 8628
rect 11756 8588 12072 8616
rect 11756 8576 11762 8588
rect 12066 8576 12072 8588
rect 12124 8616 12130 8628
rect 13262 8616 13268 8628
rect 12124 8588 13268 8616
rect 12124 8576 12130 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 18598 8576 18604 8628
rect 18656 8616 18662 8628
rect 18877 8619 18935 8625
rect 18656 8588 18828 8616
rect 18656 8576 18662 8588
rect 14642 8548 14648 8560
rect 9324 8520 14648 8548
rect 7653 8511 7711 8517
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 16669 8551 16727 8557
rect 16669 8517 16681 8551
rect 16715 8548 16727 8551
rect 18800 8548 18828 8588
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 19334 8616 19340 8628
rect 18923 8588 19340 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19760 8588 19993 8616
rect 19760 8576 19766 8588
rect 19981 8585 19993 8588
rect 20027 8585 20039 8619
rect 20806 8616 20812 8628
rect 20767 8588 20812 8616
rect 19981 8579 20039 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 16715 8520 18736 8548
rect 18800 8520 19472 8548
rect 16715 8517 16727 8520
rect 16669 8511 16727 8517
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8480 2651 8483
rect 2866 8480 2872 8492
rect 2639 8452 2872 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 2866 8440 2872 8452
rect 2924 8480 2930 8492
rect 3418 8480 3424 8492
rect 2924 8452 3424 8480
rect 2924 8440 2930 8452
rect 3418 8440 3424 8452
rect 3476 8440 3482 8492
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4157 8483 4215 8489
rect 4157 8480 4169 8483
rect 3844 8452 4169 8480
rect 3844 8440 3850 8452
rect 4157 8449 4169 8452
rect 4203 8449 4215 8483
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4157 8443 4215 8449
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5123 8452 5396 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 3694 8412 3700 8424
rect 2363 8384 3700 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 5261 8415 5319 8421
rect 5261 8412 5273 8415
rect 4764 8384 5273 8412
rect 4764 8372 4770 8384
rect 5261 8381 5273 8384
rect 5307 8381 5319 8415
rect 5368 8412 5396 8452
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 7282 8480 7288 8492
rect 6328 8452 6776 8480
rect 7243 8452 7288 8480
rect 6328 8440 6334 8452
rect 6748 8412 6776 8452
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7515 8452 7604 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7576 8412 7604 8452
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 9824 8452 10333 8480
rect 9824 8440 9830 8452
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 10413 8443 10471 8449
rect 10520 8452 16313 8480
rect 5368 8384 6684 8412
rect 6748 8384 7604 8412
rect 5261 8375 5319 8381
rect 2409 8347 2467 8353
rect 2409 8313 2421 8347
rect 2455 8344 2467 8347
rect 2866 8344 2872 8356
rect 2455 8316 2872 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 4065 8347 4123 8353
rect 3191 8316 3648 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 3237 8279 3295 8285
rect 3237 8245 3249 8279
rect 3283 8276 3295 8279
rect 3326 8276 3332 8288
rect 3283 8248 3332 8276
rect 3283 8245 3295 8248
rect 3237 8239 3295 8245
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 3620 8285 3648 8316
rect 4065 8313 4077 8347
rect 4111 8344 4123 8347
rect 4522 8344 4528 8356
rect 4111 8316 4528 8344
rect 4111 8313 4123 8316
rect 4065 8307 4123 8313
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 4801 8347 4859 8353
rect 4801 8313 4813 8347
rect 4847 8344 4859 8347
rect 5528 8347 5586 8353
rect 4847 8316 5488 8344
rect 4847 8313 4859 8316
rect 4801 8307 4859 8313
rect 3605 8279 3663 8285
rect 3605 8245 3617 8279
rect 3651 8245 3663 8279
rect 3970 8276 3976 8288
rect 3883 8248 3976 8276
rect 3605 8239 3663 8245
rect 3970 8236 3976 8248
rect 4028 8276 4034 8288
rect 4338 8276 4344 8288
rect 4028 8248 4344 8276
rect 4028 8236 4034 8248
rect 4338 8236 4344 8248
rect 4396 8236 4402 8288
rect 5460 8276 5488 8316
rect 5528 8313 5540 8347
rect 5574 8344 5586 8347
rect 6362 8344 6368 8356
rect 5574 8316 6368 8344
rect 5574 8313 5586 8316
rect 5528 8307 5586 8313
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 6656 8288 6684 8384
rect 7190 8344 7196 8356
rect 7151 8316 7196 8344
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 7576 8344 7604 8384
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 8260 8384 8401 8412
rect 8260 8372 8266 8384
rect 8389 8381 8401 8384
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 8645 8415 8703 8421
rect 8645 8412 8657 8415
rect 8536 8384 8657 8412
rect 8536 8372 8542 8384
rect 8645 8381 8657 8384
rect 8691 8381 8703 8415
rect 8645 8375 8703 8381
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 10226 8412 10232 8424
rect 9456 8384 10088 8412
rect 10187 8384 10232 8412
rect 9456 8372 9462 8384
rect 9950 8344 9956 8356
rect 7576 8316 9956 8344
rect 5718 8276 5724 8288
rect 5460 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 6638 8276 6644 8288
rect 6551 8248 6644 8276
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 9784 8285 9812 8316
rect 9950 8304 9956 8316
rect 10008 8304 10014 8356
rect 9769 8279 9827 8285
rect 9769 8245 9781 8279
rect 9815 8245 9827 8279
rect 10060 8276 10088 8384
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10428 8344 10456 8443
rect 10192 8316 10456 8344
rect 10192 8304 10198 8316
rect 10520 8276 10548 8452
rect 16301 8449 16313 8452
rect 16347 8480 16359 8483
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 16347 8452 17141 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17402 8480 17408 8492
rect 17359 8452 17408 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 17402 8440 17408 8452
rect 17460 8480 17466 8492
rect 18322 8480 18328 8492
rect 17460 8452 18328 8480
rect 17460 8440 17466 8452
rect 18322 8440 18328 8452
rect 18380 8480 18386 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 18380 8452 18613 8480
rect 18380 8440 18386 8452
rect 18601 8449 18613 8452
rect 18647 8449 18659 8483
rect 18708 8480 18736 8520
rect 19444 8489 19472 8520
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 18708 8452 19349 8480
rect 18601 8443 18659 8449
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 20533 8483 20591 8489
rect 20533 8480 20545 8483
rect 19475 8452 20545 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 20533 8449 20545 8452
rect 20579 8480 20591 8483
rect 21361 8483 21419 8489
rect 21361 8480 21373 8483
rect 20579 8452 21373 8480
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 21361 8449 21373 8452
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 11296 8384 16589 8412
rect 11296 8372 11302 8384
rect 16577 8381 16589 8384
rect 16623 8412 16635 8415
rect 17037 8415 17095 8421
rect 17037 8412 17049 8415
rect 16623 8384 17049 8412
rect 16623 8381 16635 8384
rect 16577 8375 16635 8381
rect 17037 8381 17049 8384
rect 17083 8381 17095 8415
rect 18138 8412 18144 8424
rect 17037 8375 17095 8381
rect 17328 8384 18144 8412
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 17328 8344 17356 8384
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 18230 8372 18236 8424
rect 18288 8412 18294 8424
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 18288 8384 18521 8412
rect 18288 8372 18294 8384
rect 18509 8381 18521 8384
rect 18555 8412 18567 8415
rect 19150 8412 19156 8424
rect 18555 8384 19156 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 19150 8372 19156 8384
rect 19208 8412 19214 8424
rect 19705 8415 19763 8421
rect 19705 8412 19717 8415
rect 19208 8384 19717 8412
rect 19208 8372 19214 8384
rect 19705 8381 19717 8384
rect 19751 8381 19763 8415
rect 19705 8375 19763 8381
rect 20346 8372 20352 8424
rect 20404 8412 20410 8424
rect 20441 8415 20499 8421
rect 20441 8412 20453 8415
rect 20404 8384 20453 8412
rect 20404 8372 20410 8384
rect 20441 8381 20453 8384
rect 20487 8381 20499 8415
rect 21174 8412 21180 8424
rect 21135 8384 21180 8412
rect 20441 8375 20499 8381
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 19245 8347 19303 8353
rect 19245 8344 19257 8347
rect 11020 8316 17356 8344
rect 18064 8316 19257 8344
rect 11020 8304 11026 8316
rect 18064 8285 18092 8316
rect 19245 8313 19257 8316
rect 19291 8313 19303 8347
rect 19245 8307 19303 8313
rect 20990 8304 20996 8356
rect 21048 8344 21054 8356
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 21048 8316 21281 8344
rect 21048 8304 21054 8316
rect 21269 8313 21281 8316
rect 21315 8313 21327 8347
rect 21269 8307 21327 8313
rect 10060 8248 10548 8276
rect 18049 8279 18107 8285
rect 9769 8239 9827 8245
rect 18049 8245 18061 8279
rect 18095 8245 18107 8279
rect 18414 8276 18420 8288
rect 18375 8248 18420 8276
rect 18049 8239 18107 8245
rect 18414 8236 18420 8248
rect 18472 8276 18478 8288
rect 19058 8276 19064 8288
rect 18472 8248 19064 8276
rect 18472 8236 18478 8248
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 20349 8279 20407 8285
rect 20349 8245 20361 8279
rect 20395 8276 20407 8279
rect 20438 8276 20444 8288
rect 20395 8248 20444 8276
rect 20395 8245 20407 8248
rect 20349 8239 20407 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 3418 8072 3424 8084
rect 3379 8044 3424 8072
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4522 8072 4528 8084
rect 4435 8044 4528 8072
rect 4522 8032 4528 8044
rect 4580 8072 4586 8084
rect 5074 8072 5080 8084
rect 4580 8044 5080 8072
rect 4580 8032 4586 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 6089 8075 6147 8081
rect 6089 8041 6101 8075
rect 6135 8072 6147 8075
rect 6362 8072 6368 8084
rect 6135 8044 6368 8072
rect 6135 8041 6147 8044
rect 6089 8035 6147 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 16666 8072 16672 8084
rect 9539 8044 16672 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 2056 7976 4016 8004
rect 1946 7828 1952 7880
rect 2004 7868 2010 7880
rect 2056 7877 2084 7976
rect 2308 7939 2366 7945
rect 2308 7905 2320 7939
rect 2354 7936 2366 7939
rect 3786 7936 3792 7948
rect 2354 7908 3792 7936
rect 2354 7905 2366 7908
rect 2308 7899 2366 7905
rect 3786 7896 3792 7908
rect 3844 7896 3850 7948
rect 3988 7936 4016 7976
rect 6914 7964 6920 8016
rect 6972 8004 6978 8016
rect 15378 8004 15384 8016
rect 6972 7976 15384 8004
rect 6972 7964 6978 7976
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 17212 8007 17270 8013
rect 17212 7973 17224 8007
rect 17258 8004 17270 8007
rect 20254 8004 20260 8016
rect 17258 7976 20260 8004
rect 17258 7973 17270 7976
rect 17212 7967 17270 7973
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 21082 7964 21088 8016
rect 21140 8004 21146 8016
rect 21177 8007 21235 8013
rect 21177 8004 21189 8007
rect 21140 7976 21189 8004
rect 21140 7964 21146 7976
rect 21177 7973 21189 7976
rect 21223 7973 21235 8007
rect 21177 7967 21235 7973
rect 4976 7939 5034 7945
rect 3988 7908 4200 7936
rect 2041 7871 2099 7877
rect 2041 7868 2053 7871
rect 2004 7840 2053 7868
rect 2004 7828 2010 7840
rect 2041 7837 2053 7840
rect 2087 7837 2099 7871
rect 2041 7831 2099 7837
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7868 3571 7871
rect 4062 7868 4068 7880
rect 3559 7840 4068 7868
rect 3559 7837 3571 7840
rect 3513 7831 3571 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4172 7868 4200 7908
rect 4976 7905 4988 7939
rect 5022 7936 5034 7939
rect 5442 7936 5448 7948
rect 5022 7908 5448 7936
rect 5022 7905 5034 7908
rect 4976 7899 5034 7905
rect 5442 7896 5448 7908
rect 5500 7936 5506 7948
rect 6270 7936 6276 7948
rect 5500 7908 6276 7936
rect 5500 7896 5506 7908
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6805 7939 6863 7945
rect 6805 7936 6817 7939
rect 6696 7908 6817 7936
rect 6696 7896 6702 7908
rect 6805 7905 6817 7908
rect 6851 7905 6863 7939
rect 8288 7939 8346 7945
rect 8288 7936 8300 7939
rect 6805 7899 6863 7905
rect 7944 7908 8300 7936
rect 4706 7868 4712 7880
rect 4172 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 7944 7809 7972 7908
rect 8288 7905 8300 7908
rect 8334 7936 8346 7939
rect 8570 7936 8576 7948
rect 8334 7908 8576 7936
rect 8334 7905 8346 7908
rect 8288 7899 8346 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 18046 7936 18052 7948
rect 9364 7908 18052 7936
rect 9364 7896 9370 7908
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 19604 7939 19662 7945
rect 19604 7905 19616 7939
rect 19650 7936 19662 7939
rect 20530 7936 20536 7948
rect 19650 7908 20536 7936
rect 19650 7905 19662 7908
rect 19604 7899 19662 7905
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 20622 7896 20628 7948
rect 20680 7936 20686 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 20680 7908 20913 7936
rect 20680 7896 20686 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 16942 7868 16948 7880
rect 8076 7840 8121 7868
rect 16903 7840 16948 7868
rect 8076 7828 8082 7840
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 19208 7840 19349 7868
rect 19208 7828 19214 7840
rect 19337 7837 19349 7840
rect 19383 7837 19395 7871
rect 19337 7831 19395 7837
rect 7929 7803 7987 7809
rect 4028 7772 4568 7800
rect 4028 7760 4034 7772
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3476 7704 3801 7732
rect 3476 7692 3482 7704
rect 3789 7701 3801 7704
rect 3835 7732 3847 7735
rect 4338 7732 4344 7744
rect 3835 7704 4344 7732
rect 3835 7701 3847 7704
rect 3789 7695 3847 7701
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 4540 7732 4568 7772
rect 7929 7769 7941 7803
rect 7975 7769 7987 7803
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 7929 7763 7987 7769
rect 8956 7772 9505 7800
rect 8956 7732 8984 7772
rect 9493 7769 9505 7772
rect 9539 7769 9551 7803
rect 9493 7763 9551 7769
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 18472 7772 19104 7800
rect 18472 7760 18478 7772
rect 19076 7744 19104 7772
rect 9398 7732 9404 7744
rect 4540 7704 8984 7732
rect 9359 7704 9404 7732
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 18966 7732 18972 7744
rect 16172 7704 18972 7732
rect 16172 7692 16178 7704
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 19116 7704 19161 7732
rect 19116 7692 19122 7704
rect 20254 7692 20260 7744
rect 20312 7732 20318 7744
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 20312 7704 20729 7732
rect 20312 7692 20318 7704
rect 20717 7701 20729 7704
rect 20763 7732 20775 7735
rect 21174 7732 21180 7744
rect 20763 7704 21180 7732
rect 20763 7701 20775 7704
rect 20717 7695 20775 7701
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 2866 7528 2872 7540
rect 2827 7500 2872 7528
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 3694 7528 3700 7540
rect 3655 7500 3700 7528
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 5166 7488 5172 7540
rect 5224 7528 5230 7540
rect 5350 7528 5356 7540
rect 5224 7500 5356 7528
rect 5224 7488 5230 7500
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 7285 7531 7343 7537
rect 7285 7528 7297 7531
rect 6236 7500 7297 7528
rect 6236 7488 6242 7500
rect 7285 7497 7297 7500
rect 7331 7497 7343 7531
rect 7285 7491 7343 7497
rect 8205 7531 8263 7537
rect 8205 7497 8217 7531
rect 8251 7528 8263 7531
rect 8294 7528 8300 7540
rect 8251 7500 8300 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 8294 7488 8300 7500
rect 8352 7528 8358 7540
rect 9306 7528 9312 7540
rect 8352 7500 9312 7528
rect 8352 7488 8358 7500
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 20622 7528 20628 7540
rect 20583 7500 20628 7528
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 2958 7420 2964 7472
rect 3016 7460 3022 7472
rect 3602 7460 3608 7472
rect 3016 7432 3608 7460
rect 3016 7420 3022 7432
rect 3602 7420 3608 7432
rect 3660 7420 3666 7472
rect 5442 7420 5448 7472
rect 5500 7420 5506 7472
rect 20530 7460 20536 7472
rect 20491 7432 20536 7460
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2774 7392 2780 7404
rect 2639 7364 2780 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2774 7352 2780 7364
rect 2832 7392 2838 7404
rect 3142 7392 3148 7404
rect 2832 7364 3148 7392
rect 2832 7352 2838 7364
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 3200 7364 3341 7392
rect 3200 7352 3206 7364
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3786 7392 3792 7404
rect 3559 7364 3792 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3786 7352 3792 7364
rect 3844 7392 3850 7404
rect 4341 7395 4399 7401
rect 4341 7392 4353 7395
rect 3844 7364 4353 7392
rect 3844 7352 3850 7364
rect 4341 7361 4353 7364
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4062 7324 4068 7336
rect 4023 7296 4068 7324
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 4356 7324 4384 7355
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 4856 7364 5365 7392
rect 4856 7352 4862 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5460 7392 5488 7420
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5460 7364 5549 7392
rect 5353 7355 5411 7361
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 6362 7392 6368 7404
rect 6323 7364 6368 7392
rect 5537 7355 5595 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 7742 7392 7748 7404
rect 7703 7364 7748 7392
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 9398 7392 9404 7404
rect 7975 7364 9404 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 7944 7324 7972 7355
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 19150 7392 19156 7404
rect 19111 7364 19156 7392
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 21174 7392 21180 7404
rect 21135 7364 21180 7392
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 4356 7296 7972 7324
rect 19420 7327 19478 7333
rect 19420 7293 19432 7327
rect 19466 7324 19478 7327
rect 19886 7324 19892 7336
rect 19466 7296 19892 7324
rect 19466 7293 19478 7296
rect 19420 7287 19478 7293
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 4246 7256 4252 7268
rect 3252 7228 4252 7256
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7188 2746 7200
rect 3252 7197 3280 7228
rect 4246 7216 4252 7228
rect 4304 7216 4310 7268
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 4908 7228 6193 7256
rect 3237 7191 3295 7197
rect 3237 7188 3249 7191
rect 2740 7160 3249 7188
rect 2740 7148 2746 7160
rect 3237 7157 3249 7160
rect 3283 7157 3295 7191
rect 3237 7151 3295 7157
rect 3602 7148 3608 7200
rect 3660 7188 3666 7200
rect 4157 7191 4215 7197
rect 4157 7188 4169 7191
rect 3660 7160 4169 7188
rect 3660 7148 3666 7160
rect 4157 7157 4169 7160
rect 4203 7157 4215 7191
rect 4614 7188 4620 7200
rect 4575 7160 4620 7188
rect 4157 7151 4215 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 4908 7197 4936 7228
rect 6181 7225 6193 7228
rect 6227 7225 6239 7259
rect 6181 7219 6239 7225
rect 7653 7259 7711 7265
rect 7653 7225 7665 7259
rect 7699 7256 7711 7259
rect 8294 7256 8300 7268
rect 7699 7228 8300 7256
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 21085 7259 21143 7265
rect 21085 7256 21097 7259
rect 20312 7228 21097 7256
rect 20312 7216 20318 7228
rect 21085 7225 21097 7228
rect 21131 7225 21143 7259
rect 21085 7219 21143 7225
rect 4893 7191 4951 7197
rect 4893 7157 4905 7191
rect 4939 7157 4951 7191
rect 4893 7151 4951 7157
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 5224 7160 5273 7188
rect 5224 7148 5230 7160
rect 5261 7157 5273 7160
rect 5307 7188 5319 7191
rect 5350 7188 5356 7200
rect 5307 7160 5356 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 6086 7188 6092 7200
rect 6047 7160 6092 7188
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 20622 7148 20628 7200
rect 20680 7188 20686 7200
rect 20993 7191 21051 7197
rect 20993 7188 21005 7191
rect 20680 7160 21005 7188
rect 20680 7148 20686 7160
rect 20993 7157 21005 7160
rect 21039 7157 21051 7191
rect 20993 7151 21051 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 4614 6944 4620 6996
rect 4672 6984 4678 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4672 6956 5181 6984
rect 4672 6944 4678 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 5169 6947 5227 6953
rect 2314 6876 2320 6928
rect 2372 6876 2378 6928
rect 4341 6919 4399 6925
rect 4341 6885 4353 6919
rect 4387 6916 4399 6919
rect 4798 6916 4804 6928
rect 4387 6888 4804 6916
rect 4387 6885 4399 6888
rect 4341 6879 4399 6885
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 1946 6848 1952 6860
rect 1907 6820 1952 6848
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2216 6851 2274 6857
rect 2216 6817 2228 6851
rect 2262 6848 2274 6851
rect 2332 6848 2360 6876
rect 3421 6851 3479 6857
rect 3421 6848 3433 6851
rect 2262 6820 3433 6848
rect 2262 6817 2274 6820
rect 2216 6811 2274 6817
rect 3421 6817 3433 6820
rect 3467 6817 3479 6851
rect 3421 6811 3479 6817
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 14734 6848 14740 6860
rect 4120 6820 14740 6848
rect 4120 6808 4126 6820
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 20441 6851 20499 6857
rect 20441 6817 20453 6851
rect 20487 6848 20499 6851
rect 20622 6848 20628 6860
rect 20487 6820 20628 6848
rect 20487 6817 20499 6820
rect 20441 6811 20499 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4448 6752 5273 6780
rect 3329 6715 3387 6721
rect 3329 6681 3341 6715
rect 3375 6712 3387 6715
rect 3878 6712 3884 6724
rect 3375 6684 3884 6712
rect 3375 6681 3387 6684
rect 3329 6675 3387 6681
rect 3878 6672 3884 6684
rect 3936 6672 3942 6724
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4448 6721 4476 6752
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5261 6743 5319 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 17954 6780 17960 6792
rect 9088 6752 17960 6780
rect 9088 6740 9094 6752
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 4433 6715 4491 6721
rect 4433 6712 4445 6715
rect 4212 6684 4445 6712
rect 4212 6672 4218 6684
rect 4433 6681 4445 6684
rect 4479 6681 4491 6715
rect 4433 6675 4491 6681
rect 4801 6715 4859 6721
rect 4801 6681 4813 6715
rect 4847 6712 4859 6715
rect 6086 6712 6092 6724
rect 4847 6684 6092 6712
rect 4847 6681 4859 6684
rect 4801 6675 4859 6681
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 3602 6644 3608 6656
rect 3563 6616 3608 6644
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4396 6616 4629 6644
rect 4396 6604 4402 6616
rect 4617 6613 4629 6616
rect 4663 6644 4675 6647
rect 5166 6644 5172 6656
rect 4663 6616 5172 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 11882 6440 11888 6452
rect 4028 6412 11888 6440
rect 4028 6400 4034 6412
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 20254 6440 20260 6452
rect 20215 6412 20260 6440
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 5258 6332 5264 6384
rect 5316 6372 5322 6384
rect 9582 6372 9588 6384
rect 5316 6344 9588 6372
rect 5316 6332 5322 6344
rect 9582 6332 9588 6344
rect 9640 6332 9646 6384
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20588 6276 20821 6304
rect 20588 6264 20594 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 20625 6171 20683 6177
rect 20625 6168 20637 6171
rect 20088 6140 20637 6168
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 20088 6109 20116 6140
rect 20625 6137 20637 6140
rect 20671 6137 20683 6171
rect 20625 6131 20683 6137
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 3384 6072 20085 6100
rect 3384 6060 3390 6072
rect 20073 6069 20085 6072
rect 20119 6069 20131 6103
rect 20073 6063 20131 6069
rect 20530 6060 20536 6112
rect 20588 6100 20594 6112
rect 20717 6103 20775 6109
rect 20717 6100 20729 6103
rect 20588 6072 20729 6100
rect 20588 6060 20594 6072
rect 20717 6069 20729 6072
rect 20763 6100 20775 6103
rect 21085 6103 21143 6109
rect 21085 6100 21097 6103
rect 20763 6072 21097 6100
rect 20763 6069 20775 6072
rect 20717 6063 20775 6069
rect 21085 6069 21097 6072
rect 21131 6069 21143 6103
rect 21085 6063 21143 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 17954 5352 17960 5364
rect 5868 5324 17960 5352
rect 5868 5312 5874 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 6454 5284 6460 5296
rect 4120 5256 6460 5284
rect 4120 5244 4126 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 9640 3080 15700 3108
rect 9640 3068 9646 3080
rect 15672 3049 15700 3080
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 4816 3012 5457 3040
rect 4816 2981 4844 3012
rect 5445 3009 5457 3012
rect 5491 3040 5503 3043
rect 15657 3043 15715 3049
rect 5491 3012 5948 3040
rect 5491 3009 5503 3012
rect 5445 3003 5503 3009
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2941 4859 2975
rect 4801 2935 4859 2941
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 5040 2944 5089 2972
rect 5040 2932 5046 2944
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 5552 2836 5580 2935
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 5813 2975 5871 2981
rect 5813 2972 5825 2975
rect 5684 2944 5825 2972
rect 5684 2932 5690 2944
rect 5813 2941 5825 2944
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 5920 2904 5948 3012
rect 15657 3009 15669 3043
rect 15703 3009 15715 3043
rect 15657 3003 15715 3009
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15519 2944 16037 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 16025 2941 16037 2944
rect 16071 2972 16083 2975
rect 16114 2972 16120 2984
rect 16071 2944 16120 2972
rect 16071 2941 16083 2944
rect 16025 2935 16083 2941
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 20714 2904 20720 2916
rect 5920 2876 20720 2904
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 5552 2808 6193 2836
rect 6181 2805 6193 2808
rect 6227 2836 6239 2839
rect 11238 2836 11244 2848
rect 6227 2808 11244 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 3326 1980 3332 2032
rect 3384 2020 3390 2032
rect 4798 2020 4804 2032
rect 3384 1992 4804 2020
rect 3384 1980 3390 1992
rect 4798 1980 4804 1992
rect 4856 1980 4862 2032
rect 4062 1164 4068 1216
rect 4120 1204 4126 1216
rect 7190 1204 7196 1216
rect 4120 1176 7196 1204
rect 4120 1164 4126 1176
rect 7190 1164 7196 1176
rect 7248 1164 7254 1216
<< via1 >>
rect 4068 21088 4120 21140
rect 6368 21088 6420 21140
rect 2320 20884 2372 20936
rect 3056 20884 3108 20936
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 18604 20544 18656 20596
rect 19708 20544 19760 20596
rect 9680 20476 9732 20528
rect 18052 20476 18104 20528
rect 10048 20408 10100 20460
rect 2228 20340 2280 20392
rect 14096 20340 14148 20392
rect 14648 20340 14700 20392
rect 17132 20383 17184 20392
rect 17132 20349 17141 20383
rect 17141 20349 17175 20383
rect 17175 20349 17184 20383
rect 17132 20340 17184 20349
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 19064 20340 19116 20392
rect 8852 20272 8904 20324
rect 14556 20272 14608 20324
rect 15108 20272 15160 20324
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 2136 20204 2188 20256
rect 7288 20204 7340 20256
rect 9220 20247 9272 20256
rect 9220 20213 9229 20247
rect 9229 20213 9263 20247
rect 9263 20213 9272 20247
rect 9220 20204 9272 20213
rect 13084 20204 13136 20256
rect 17224 20204 17276 20256
rect 20352 20247 20404 20256
rect 20352 20213 20361 20247
rect 20361 20213 20395 20247
rect 20395 20213 20404 20247
rect 20352 20204 20404 20213
rect 21180 20204 21232 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2780 20000 2832 20052
rect 9220 20000 9272 20052
rect 13084 20043 13136 20052
rect 1492 19907 1544 19916
rect 1492 19873 1501 19907
rect 1501 19873 1535 19907
rect 1535 19873 1544 19907
rect 1492 19864 1544 19873
rect 2136 19864 2188 19916
rect 2228 19907 2280 19916
rect 2228 19873 2237 19907
rect 2237 19873 2271 19907
rect 2271 19873 2280 19907
rect 2228 19864 2280 19873
rect 3424 19932 3476 19984
rect 8484 19864 8536 19916
rect 10048 19932 10100 19984
rect 10600 19864 10652 19916
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 14372 20000 14424 20052
rect 14556 20043 14608 20052
rect 14556 20009 14565 20043
rect 14565 20009 14599 20043
rect 14599 20009 14608 20043
rect 14556 20000 14608 20009
rect 15476 20043 15528 20052
rect 15476 20009 15485 20043
rect 15485 20009 15519 20043
rect 15519 20009 15528 20043
rect 15476 20000 15528 20009
rect 15936 20000 15988 20052
rect 17592 20000 17644 20052
rect 18880 20000 18932 20052
rect 20628 20000 20680 20052
rect 12532 19932 12584 19984
rect 17500 19932 17552 19984
rect 3240 19796 3292 19848
rect 9404 19839 9456 19848
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 2412 19703 2464 19712
rect 2412 19669 2421 19703
rect 2421 19669 2455 19703
rect 2455 19669 2464 19703
rect 2412 19660 2464 19669
rect 4068 19660 4120 19712
rect 8300 19660 8352 19712
rect 9404 19805 9413 19839
rect 9413 19805 9447 19839
rect 9447 19805 9456 19839
rect 9404 19796 9456 19805
rect 9772 19796 9824 19848
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 15292 19907 15344 19916
rect 12072 19796 12124 19805
rect 11704 19728 11756 19780
rect 12164 19728 12216 19780
rect 13544 19771 13596 19780
rect 13544 19737 13553 19771
rect 13553 19737 13587 19771
rect 13587 19737 13596 19771
rect 13544 19728 13596 19737
rect 9312 19660 9364 19712
rect 12624 19660 12676 19712
rect 13176 19660 13228 19712
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 16580 19864 16632 19916
rect 19340 19907 19392 19916
rect 15568 19796 15620 19848
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 18052 19796 18104 19848
rect 14556 19728 14608 19780
rect 19248 19796 19300 19848
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 14464 19660 14516 19712
rect 20812 19864 20864 19916
rect 21180 19864 21232 19916
rect 21456 19864 21508 19916
rect 20536 19728 20588 19780
rect 22284 19660 22336 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 3148 19499 3200 19508
rect 3148 19465 3157 19499
rect 3157 19465 3191 19499
rect 3191 19465 3200 19499
rect 3148 19456 3200 19465
rect 3608 19499 3660 19508
rect 3608 19465 3617 19499
rect 3617 19465 3651 19499
rect 3651 19465 3660 19499
rect 3608 19456 3660 19465
rect 6368 19499 6420 19508
rect 6368 19465 6377 19499
rect 6377 19465 6411 19499
rect 6411 19465 6420 19499
rect 6368 19456 6420 19465
rect 9404 19456 9456 19508
rect 10048 19456 10100 19508
rect 10600 19456 10652 19508
rect 14372 19456 14424 19508
rect 16120 19456 16172 19508
rect 18052 19499 18104 19508
rect 18052 19465 18061 19499
rect 18061 19465 18095 19499
rect 18095 19465 18104 19499
rect 18052 19456 18104 19465
rect 20720 19456 20772 19508
rect 20996 19499 21048 19508
rect 20996 19465 21005 19499
rect 21005 19465 21039 19499
rect 21039 19465 21048 19499
rect 20996 19456 21048 19465
rect 21364 19499 21416 19508
rect 21364 19465 21373 19499
rect 21373 19465 21407 19499
rect 21407 19465 21416 19499
rect 21364 19456 21416 19465
rect 2596 19388 2648 19440
rect 1584 19252 1636 19304
rect 204 19184 256 19236
rect 1308 19184 1360 19236
rect 2320 19252 2372 19304
rect 14924 19388 14976 19440
rect 2780 19252 2832 19304
rect 3148 19252 3200 19304
rect 3516 19252 3568 19304
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 6828 19252 6880 19304
rect 7012 19252 7064 19304
rect 9404 19295 9456 19304
rect 9404 19261 9438 19295
rect 9438 19261 9456 19295
rect 9404 19252 9456 19261
rect 10876 19295 10928 19304
rect 10876 19261 10885 19295
rect 10885 19261 10919 19295
rect 10919 19261 10928 19295
rect 10876 19252 10928 19261
rect 12624 19252 12676 19304
rect 16028 19320 16080 19372
rect 17132 19320 17184 19372
rect 18604 19363 18656 19372
rect 18604 19329 18613 19363
rect 18613 19329 18647 19363
rect 18647 19329 18656 19363
rect 18604 19320 18656 19329
rect 1860 19116 1912 19168
rect 2044 19159 2096 19168
rect 2044 19125 2053 19159
rect 2053 19125 2087 19159
rect 2087 19125 2096 19159
rect 2044 19116 2096 19125
rect 3056 19184 3108 19236
rect 4344 19184 4396 19236
rect 7564 19184 7616 19236
rect 2872 19116 2924 19168
rect 8300 19116 8352 19168
rect 10600 19159 10652 19168
rect 10600 19125 10609 19159
rect 10609 19125 10643 19159
rect 10643 19125 10652 19159
rect 12348 19184 12400 19236
rect 13084 19184 13136 19236
rect 10600 19116 10652 19125
rect 12072 19116 12124 19168
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 14372 19159 14424 19168
rect 14372 19125 14381 19159
rect 14381 19125 14415 19159
rect 14415 19125 14424 19159
rect 14372 19116 14424 19125
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 17408 19295 17460 19304
rect 17408 19261 17417 19295
rect 17417 19261 17451 19295
rect 17451 19261 17460 19295
rect 17408 19252 17460 19261
rect 17868 19252 17920 19304
rect 19984 19252 20036 19304
rect 20352 19252 20404 19304
rect 20720 19252 20772 19304
rect 14924 19184 14976 19236
rect 16764 19184 16816 19236
rect 14464 19116 14516 19125
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 15384 19116 15436 19168
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 16304 19116 16356 19168
rect 17960 19184 18012 19236
rect 19708 19184 19760 19236
rect 18052 19116 18104 19168
rect 19524 19116 19576 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1308 18912 1360 18964
rect 1768 18912 1820 18964
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 2964 18912 3016 18964
rect 3148 18912 3200 18964
rect 3792 18912 3844 18964
rect 8300 18912 8352 18964
rect 8852 18912 8904 18964
rect 10600 18912 10652 18964
rect 11336 18912 11388 18964
rect 11980 18912 12032 18964
rect 12072 18912 12124 18964
rect 16120 18912 16172 18964
rect 6828 18887 6880 18896
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 2320 18708 2372 18760
rect 2504 18640 2556 18692
rect 2688 18683 2740 18692
rect 2688 18649 2697 18683
rect 2697 18649 2731 18683
rect 2731 18649 2740 18683
rect 2688 18640 2740 18649
rect 3608 18708 3660 18760
rect 6828 18853 6837 18887
rect 6837 18853 6871 18887
rect 6871 18853 6880 18887
rect 6828 18844 6880 18853
rect 7564 18844 7616 18896
rect 5448 18776 5500 18828
rect 6460 18776 6512 18828
rect 6644 18776 6696 18828
rect 8300 18776 8352 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 9680 18819 9732 18828
rect 8392 18776 8444 18785
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 13912 18887 13964 18896
rect 10600 18776 10652 18828
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 12072 18819 12124 18828
rect 8852 18708 8904 18760
rect 9404 18751 9456 18760
rect 1584 18572 1636 18624
rect 2780 18572 2832 18624
rect 3516 18640 3568 18692
rect 6644 18640 6696 18692
rect 8760 18640 8812 18692
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 9956 18751 10008 18760
rect 9956 18717 9965 18751
rect 9965 18717 9999 18751
rect 9999 18717 10008 18751
rect 9956 18708 10008 18717
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 13912 18853 13946 18887
rect 13946 18853 13964 18887
rect 13912 18844 13964 18853
rect 14464 18844 14516 18896
rect 12900 18819 12952 18828
rect 9588 18640 9640 18692
rect 11336 18751 11388 18760
rect 11336 18717 11345 18751
rect 11345 18717 11379 18751
rect 11379 18717 11388 18751
rect 11336 18708 11388 18717
rect 11980 18708 12032 18760
rect 12348 18751 12400 18760
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 12900 18785 12909 18819
rect 12909 18785 12943 18819
rect 12943 18785 12952 18819
rect 12900 18776 12952 18785
rect 14188 18776 14240 18828
rect 14648 18776 14700 18828
rect 17408 18844 17460 18896
rect 19432 18912 19484 18964
rect 21088 18955 21140 18964
rect 21088 18921 21097 18955
rect 21097 18921 21131 18955
rect 21131 18921 21140 18955
rect 21088 18912 21140 18921
rect 21548 18912 21600 18964
rect 18604 18887 18656 18896
rect 18604 18853 18638 18887
rect 18638 18853 18656 18887
rect 18604 18844 18656 18853
rect 19248 18844 19300 18896
rect 12992 18751 13044 18760
rect 12992 18717 13001 18751
rect 13001 18717 13035 18751
rect 13035 18717 13044 18751
rect 12992 18708 13044 18717
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 15844 18751 15896 18760
rect 13084 18708 13136 18717
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 12532 18683 12584 18692
rect 6000 18572 6052 18624
rect 6184 18615 6236 18624
rect 6184 18581 6193 18615
rect 6193 18581 6227 18615
rect 6227 18581 6236 18615
rect 6184 18572 6236 18581
rect 8484 18572 8536 18624
rect 11704 18572 11756 18624
rect 12532 18649 12541 18683
rect 12541 18649 12575 18683
rect 12575 18649 12584 18683
rect 12532 18640 12584 18649
rect 16764 18776 16816 18828
rect 17500 18776 17552 18828
rect 20168 18819 20220 18828
rect 20168 18785 20177 18819
rect 20177 18785 20211 18819
rect 20211 18785 20220 18819
rect 20168 18776 20220 18785
rect 16672 18708 16724 18760
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 17868 18708 17920 18760
rect 19432 18708 19484 18760
rect 20444 18776 20496 18828
rect 20904 18819 20956 18828
rect 20904 18785 20913 18819
rect 20913 18785 20947 18819
rect 20947 18785 20956 18819
rect 20904 18776 20956 18785
rect 21364 18776 21416 18828
rect 19708 18683 19760 18692
rect 19708 18649 19717 18683
rect 19717 18649 19751 18683
rect 19751 18649 19760 18683
rect 19708 18640 19760 18649
rect 18144 18572 18196 18624
rect 20720 18615 20772 18624
rect 20720 18581 20729 18615
rect 20729 18581 20763 18615
rect 20763 18581 20772 18615
rect 20720 18572 20772 18581
rect 21732 18572 21784 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2872 18368 2924 18420
rect 3424 18368 3476 18420
rect 5724 18368 5776 18420
rect 10416 18368 10468 18420
rect 13912 18411 13964 18420
rect 1032 18300 1084 18352
rect 8116 18300 8168 18352
rect 8300 18300 8352 18352
rect 9588 18300 9640 18352
rect 9956 18300 10008 18352
rect 12256 18300 12308 18352
rect 13912 18377 13921 18411
rect 13921 18377 13955 18411
rect 13955 18377 13964 18411
rect 13912 18368 13964 18377
rect 14372 18368 14424 18420
rect 14464 18411 14516 18420
rect 14464 18377 14473 18411
rect 14473 18377 14507 18411
rect 14507 18377 14516 18411
rect 14464 18368 14516 18377
rect 15568 18368 15620 18420
rect 16028 18411 16080 18420
rect 16028 18377 16037 18411
rect 16037 18377 16071 18411
rect 16071 18377 16080 18411
rect 16028 18368 16080 18377
rect 17500 18411 17552 18420
rect 17500 18377 17509 18411
rect 17509 18377 17543 18411
rect 17543 18377 17552 18411
rect 17500 18368 17552 18377
rect 18052 18411 18104 18420
rect 18052 18377 18061 18411
rect 18061 18377 18095 18411
rect 18095 18377 18104 18411
rect 18052 18368 18104 18377
rect 18696 18368 18748 18420
rect 19248 18411 19300 18420
rect 19248 18377 19257 18411
rect 19257 18377 19291 18411
rect 19291 18377 19300 18411
rect 19248 18368 19300 18377
rect 19340 18368 19392 18420
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 17132 18300 17184 18352
rect 1400 18232 1452 18284
rect 2596 18232 2648 18284
rect 5448 18275 5500 18284
rect 2964 18164 3016 18216
rect 2320 18028 2372 18080
rect 2504 18028 2556 18080
rect 4160 18164 4212 18216
rect 5172 18207 5224 18216
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 5172 18164 5224 18173
rect 5448 18241 5457 18275
rect 5457 18241 5491 18275
rect 5491 18241 5500 18275
rect 5448 18232 5500 18241
rect 6552 18232 6604 18284
rect 7472 18232 7524 18284
rect 7564 18232 7616 18284
rect 8392 18275 8444 18284
rect 8392 18241 8401 18275
rect 8401 18241 8435 18275
rect 8435 18241 8444 18275
rect 8392 18232 8444 18241
rect 8484 18232 8536 18284
rect 10140 18232 10192 18284
rect 11704 18232 11756 18284
rect 12900 18232 12952 18284
rect 16028 18232 16080 18284
rect 6828 18164 6880 18216
rect 6920 18164 6972 18216
rect 3332 18096 3384 18148
rect 4896 18096 4948 18148
rect 3700 18028 3752 18080
rect 6736 18028 6788 18080
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 7656 18071 7708 18080
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 8392 18028 8444 18080
rect 8668 18028 8720 18080
rect 10140 18028 10192 18080
rect 11244 18164 11296 18216
rect 14096 18164 14148 18216
rect 14188 18164 14240 18216
rect 14740 18164 14792 18216
rect 15844 18164 15896 18216
rect 17500 18232 17552 18284
rect 19708 18232 19760 18284
rect 11704 18096 11756 18148
rect 11980 18096 12032 18148
rect 16672 18096 16724 18148
rect 10876 18028 10928 18080
rect 11796 18028 11848 18080
rect 15752 18028 15804 18080
rect 17684 18028 17736 18080
rect 18052 18028 18104 18080
rect 20720 18164 20772 18216
rect 20904 18096 20956 18148
rect 20536 18028 20588 18080
rect 20720 18071 20772 18080
rect 20720 18037 20729 18071
rect 20729 18037 20763 18071
rect 20763 18037 20772 18071
rect 20720 18028 20772 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 5172 17824 5224 17876
rect 6920 17824 6972 17876
rect 7288 17824 7340 17876
rect 7656 17824 7708 17876
rect 8208 17824 8260 17876
rect 8852 17824 8904 17876
rect 9312 17867 9364 17876
rect 9312 17833 9321 17867
rect 9321 17833 9355 17867
rect 9355 17833 9364 17867
rect 9312 17824 9364 17833
rect 11060 17824 11112 17876
rect 1768 17756 1820 17808
rect 5540 17756 5592 17808
rect 6828 17756 6880 17808
rect 13912 17824 13964 17876
rect 15384 17824 15436 17876
rect 15752 17867 15804 17876
rect 15752 17833 15761 17867
rect 15761 17833 15795 17867
rect 15795 17833 15804 17867
rect 15752 17824 15804 17833
rect 17960 17824 18012 17876
rect 21088 17867 21140 17876
rect 21088 17833 21097 17867
rect 21097 17833 21131 17867
rect 21131 17833 21140 17867
rect 21088 17824 21140 17833
rect 17408 17756 17460 17808
rect 17684 17756 17736 17808
rect 18788 17756 18840 17808
rect 19984 17756 20036 17808
rect 4252 17620 4304 17672
rect 6000 17688 6052 17740
rect 6736 17688 6788 17740
rect 7104 17731 7156 17740
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 7840 17620 7892 17672
rect 2320 17484 2372 17536
rect 4804 17484 4856 17536
rect 6368 17484 6420 17536
rect 6460 17484 6512 17536
rect 8484 17552 8536 17604
rect 10876 17688 10928 17740
rect 9772 17663 9824 17672
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 7380 17484 7432 17536
rect 9680 17484 9732 17536
rect 11244 17552 11296 17604
rect 11980 17620 12032 17672
rect 14464 17688 14516 17740
rect 20260 17688 20312 17740
rect 12992 17620 13044 17672
rect 15476 17620 15528 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 13544 17552 13596 17604
rect 13636 17552 13688 17604
rect 17500 17663 17552 17672
rect 17500 17629 17509 17663
rect 17509 17629 17543 17663
rect 17543 17629 17552 17663
rect 20352 17663 20404 17672
rect 17500 17620 17552 17629
rect 20352 17629 20361 17663
rect 20361 17629 20395 17663
rect 20395 17629 20404 17663
rect 20352 17620 20404 17629
rect 11980 17484 12032 17536
rect 12716 17484 12768 17536
rect 13452 17484 13504 17536
rect 17408 17484 17460 17536
rect 20536 17552 20588 17604
rect 17868 17527 17920 17536
rect 17868 17493 17877 17527
rect 17877 17493 17911 17527
rect 17911 17493 17920 17527
rect 17868 17484 17920 17493
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 20168 17484 20220 17536
rect 21088 17484 21140 17536
rect 21364 17484 21416 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2688 17280 2740 17332
rect 2964 17280 3016 17332
rect 6000 17323 6052 17332
rect 4528 17255 4580 17264
rect 4528 17221 4537 17255
rect 4537 17221 4571 17255
rect 4571 17221 4580 17255
rect 4528 17212 4580 17221
rect 2688 17187 2740 17196
rect 2688 17153 2697 17187
rect 2697 17153 2731 17187
rect 2731 17153 2740 17187
rect 2688 17144 2740 17153
rect 2780 17144 2832 17196
rect 2964 17144 3016 17196
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 7840 17280 7892 17332
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 8392 17323 8444 17332
rect 8392 17289 8401 17323
rect 8401 17289 8435 17323
rect 8435 17289 8444 17323
rect 8392 17280 8444 17289
rect 9312 17280 9364 17332
rect 10048 17280 10100 17332
rect 11060 17280 11112 17332
rect 8852 17212 8904 17264
rect 11704 17280 11756 17332
rect 11980 17280 12032 17332
rect 12256 17280 12308 17332
rect 13544 17280 13596 17332
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 3148 17119 3200 17128
rect 3148 17085 3157 17119
rect 3157 17085 3191 17119
rect 3191 17085 3200 17119
rect 3148 17076 3200 17085
rect 5172 17076 5224 17128
rect 6184 17076 6236 17128
rect 8484 17144 8536 17196
rect 9680 17144 9732 17196
rect 9864 17144 9916 17196
rect 9956 17144 10008 17196
rect 10416 17144 10468 17196
rect 10692 17144 10744 17196
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 9312 17119 9364 17128
rect 3976 17008 4028 17060
rect 4528 17008 4580 17060
rect 4804 17008 4856 17060
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 12716 17212 12768 17264
rect 16488 17212 16540 17264
rect 17868 17212 17920 17264
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 13176 17144 13228 17196
rect 13544 17144 13596 17196
rect 13728 17144 13780 17196
rect 7012 17008 7064 17060
rect 7564 17008 7616 17060
rect 8208 17008 8260 17060
rect 6276 16940 6328 16992
rect 8760 16983 8812 16992
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 8760 16940 8812 16949
rect 9680 16940 9732 16992
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 10048 16940 10100 16992
rect 10324 16940 10376 16992
rect 11888 17008 11940 17060
rect 12256 17008 12308 17060
rect 13636 17008 13688 17060
rect 11428 16940 11480 16992
rect 12348 16940 12400 16992
rect 13084 16983 13136 16992
rect 13084 16949 13093 16983
rect 13093 16949 13127 16983
rect 13127 16949 13136 16983
rect 13084 16940 13136 16949
rect 13912 16940 13964 16992
rect 15292 17144 15344 17196
rect 17040 17144 17092 17196
rect 18512 17076 18564 17128
rect 19156 17119 19208 17128
rect 19156 17085 19165 17119
rect 19165 17085 19199 17119
rect 19199 17085 19208 17119
rect 19156 17076 19208 17085
rect 20720 17212 20772 17264
rect 20720 17119 20772 17128
rect 15292 17008 15344 17060
rect 15476 17008 15528 17060
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 19340 17008 19392 17060
rect 20536 17008 20588 17060
rect 14464 16983 14516 16992
rect 14464 16949 14473 16983
rect 14473 16949 14507 16983
rect 14507 16949 14516 16983
rect 14464 16940 14516 16949
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 15568 16940 15620 16949
rect 18972 16940 19024 16992
rect 20904 16940 20956 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 4896 16736 4948 16788
rect 7380 16736 7432 16788
rect 7564 16779 7616 16788
rect 7564 16745 7573 16779
rect 7573 16745 7607 16779
rect 7607 16745 7616 16779
rect 7564 16736 7616 16745
rect 9864 16736 9916 16788
rect 12072 16736 12124 16788
rect 3056 16600 3108 16652
rect 8300 16668 8352 16720
rect 9312 16668 9364 16720
rect 15568 16736 15620 16788
rect 18512 16779 18564 16788
rect 13452 16668 13504 16720
rect 16580 16711 16632 16720
rect 16580 16677 16589 16711
rect 16589 16677 16623 16711
rect 16623 16677 16632 16711
rect 16580 16668 16632 16677
rect 572 16532 624 16584
rect 4160 16600 4212 16652
rect 4344 16600 4396 16652
rect 5816 16643 5868 16652
rect 5816 16609 5825 16643
rect 5825 16609 5859 16643
rect 5859 16609 5868 16643
rect 5816 16600 5868 16609
rect 6184 16643 6236 16652
rect 6184 16609 6193 16643
rect 6193 16609 6227 16643
rect 6227 16609 6236 16643
rect 6184 16600 6236 16609
rect 6460 16643 6512 16652
rect 6460 16609 6494 16643
rect 6494 16609 6512 16643
rect 6460 16600 6512 16609
rect 7012 16600 7064 16652
rect 9772 16600 9824 16652
rect 11704 16643 11756 16652
rect 11704 16609 11738 16643
rect 11738 16609 11756 16643
rect 11704 16600 11756 16609
rect 13084 16600 13136 16652
rect 14648 16600 14700 16652
rect 16304 16643 16356 16652
rect 16304 16609 16313 16643
rect 16313 16609 16347 16643
rect 16347 16609 16356 16643
rect 16304 16600 16356 16609
rect 17500 16600 17552 16652
rect 18512 16745 18521 16779
rect 18521 16745 18555 16779
rect 18555 16745 18564 16779
rect 18512 16736 18564 16745
rect 19708 16736 19760 16788
rect 21088 16779 21140 16788
rect 21088 16745 21097 16779
rect 21097 16745 21131 16779
rect 21131 16745 21140 16779
rect 21088 16736 21140 16745
rect 17776 16668 17828 16720
rect 19156 16668 19208 16720
rect 3884 16532 3936 16584
rect 3976 16532 4028 16584
rect 5908 16532 5960 16584
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 10416 16532 10468 16584
rect 2688 16464 2740 16516
rect 1768 16396 1820 16448
rect 3332 16396 3384 16448
rect 4344 16396 4396 16448
rect 4896 16439 4948 16448
rect 4896 16405 4905 16439
rect 4905 16405 4939 16439
rect 4939 16405 4948 16439
rect 4896 16396 4948 16405
rect 9956 16464 10008 16516
rect 11152 16532 11204 16584
rect 13544 16575 13596 16584
rect 8760 16396 8812 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 12716 16464 12768 16516
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 14280 16575 14332 16584
rect 13544 16532 13596 16541
rect 13728 16507 13780 16516
rect 13728 16473 13737 16507
rect 13737 16473 13771 16507
rect 13771 16473 13780 16507
rect 13728 16464 13780 16473
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 16672 16532 16724 16584
rect 19248 16600 19300 16652
rect 20352 16600 20404 16652
rect 20904 16643 20956 16652
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 20904 16600 20956 16609
rect 19064 16532 19116 16584
rect 11796 16396 11848 16448
rect 13268 16396 13320 16448
rect 13820 16396 13872 16448
rect 13912 16396 13964 16448
rect 14740 16396 14792 16448
rect 15200 16396 15252 16448
rect 18052 16396 18104 16448
rect 19340 16396 19392 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2872 16192 2924 16244
rect 3976 16235 4028 16244
rect 3976 16201 3985 16235
rect 3985 16201 4019 16235
rect 4019 16201 4028 16235
rect 3976 16192 4028 16201
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 5540 16192 5592 16244
rect 7104 16192 7156 16244
rect 11244 16192 11296 16244
rect 11704 16192 11756 16244
rect 12072 16192 12124 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 4160 16167 4212 16176
rect 4160 16133 4169 16167
rect 4169 16133 4203 16167
rect 4203 16133 4212 16167
rect 4160 16124 4212 16133
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 2320 15988 2372 16040
rect 3148 15988 3200 16040
rect 3332 15988 3384 16040
rect 3792 15988 3844 16040
rect 9864 16124 9916 16176
rect 4344 16056 4396 16108
rect 4804 16099 4856 16108
rect 4804 16065 4813 16099
rect 4813 16065 4847 16099
rect 4847 16065 4856 16099
rect 4804 16056 4856 16065
rect 7564 16056 7616 16108
rect 8484 16056 8536 16108
rect 4896 15988 4948 16040
rect 7380 15988 7432 16040
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10048 15988 10100 16040
rect 3884 15920 3936 15972
rect 4988 15920 5040 15972
rect 5172 15852 5224 15904
rect 7564 15852 7616 15904
rect 8852 15920 8904 15972
rect 11796 15988 11848 16040
rect 12072 15988 12124 16040
rect 12716 16031 12768 16040
rect 12716 15997 12750 16031
rect 12750 15997 12768 16031
rect 10416 15963 10468 15972
rect 10416 15929 10450 15963
rect 10450 15929 10468 15963
rect 10416 15920 10468 15929
rect 12716 15988 12768 15997
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 16396 16056 16448 16108
rect 17224 16124 17276 16176
rect 18696 16192 18748 16244
rect 19432 16192 19484 16244
rect 21272 16235 21324 16244
rect 21272 16201 21281 16235
rect 21281 16201 21315 16235
rect 21315 16201 21324 16235
rect 21272 16192 21324 16201
rect 20352 16124 20404 16176
rect 17316 16031 17368 16040
rect 8208 15852 8260 15904
rect 9680 15852 9732 15904
rect 9864 15852 9916 15904
rect 11612 15895 11664 15904
rect 11612 15861 11621 15895
rect 11621 15861 11655 15895
rect 11655 15861 11664 15895
rect 11612 15852 11664 15861
rect 13728 15852 13780 15904
rect 14280 15920 14332 15972
rect 14740 15920 14792 15972
rect 17316 15997 17325 16031
rect 17325 15997 17359 16031
rect 17359 15997 17368 16031
rect 17316 15988 17368 15997
rect 17776 15988 17828 16040
rect 19524 15988 19576 16040
rect 19984 15988 20036 16040
rect 16672 15920 16724 15972
rect 14096 15852 14148 15904
rect 18880 15920 18932 15972
rect 19156 15920 19208 15972
rect 19248 15920 19300 15972
rect 17960 15852 18012 15904
rect 20536 15852 20588 15904
rect 21272 15852 21324 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2780 15648 2832 15700
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 6184 15648 6236 15700
rect 7564 15648 7616 15700
rect 9404 15648 9456 15700
rect 10876 15648 10928 15700
rect 14464 15648 14516 15700
rect 15936 15648 15988 15700
rect 17500 15691 17552 15700
rect 4252 15512 4304 15564
rect 5356 15512 5408 15564
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 5540 15444 5592 15496
rect 5908 15444 5960 15496
rect 8208 15580 8260 15632
rect 7380 15512 7432 15564
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 6276 15444 6328 15496
rect 9956 15555 10008 15564
rect 9956 15521 9990 15555
rect 9990 15521 10008 15555
rect 9956 15512 10008 15521
rect 11704 15580 11756 15632
rect 11796 15580 11848 15632
rect 15200 15580 15252 15632
rect 15752 15623 15804 15632
rect 7380 15419 7432 15428
rect 2136 15308 2188 15360
rect 7380 15385 7389 15419
rect 7389 15385 7423 15419
rect 7423 15385 7432 15419
rect 7380 15376 7432 15385
rect 8208 15376 8260 15428
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 8852 15444 8904 15496
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 11244 15444 11296 15496
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 11152 15376 11204 15428
rect 11888 15376 11940 15428
rect 6736 15308 6788 15360
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 9864 15308 9916 15360
rect 10324 15308 10376 15360
rect 10416 15308 10468 15360
rect 13728 15512 13780 15564
rect 15752 15589 15761 15623
rect 15761 15589 15795 15623
rect 15795 15589 15804 15623
rect 15752 15580 15804 15589
rect 16396 15623 16448 15632
rect 16396 15589 16430 15623
rect 16430 15589 16448 15623
rect 16396 15580 16448 15589
rect 17500 15657 17509 15691
rect 17509 15657 17543 15691
rect 17543 15657 17552 15691
rect 17500 15648 17552 15657
rect 19156 15691 19208 15700
rect 19156 15657 19165 15691
rect 19165 15657 19199 15691
rect 19199 15657 19208 15691
rect 19156 15648 19208 15657
rect 19248 15691 19300 15700
rect 19248 15657 19257 15691
rect 19257 15657 19291 15691
rect 19291 15657 19300 15691
rect 20628 15691 20680 15700
rect 19248 15648 19300 15657
rect 20628 15657 20637 15691
rect 20637 15657 20671 15691
rect 20671 15657 20680 15691
rect 20628 15648 20680 15657
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 21456 15691 21508 15700
rect 21456 15657 21465 15691
rect 21465 15657 21499 15691
rect 21499 15657 21508 15691
rect 21456 15648 21508 15657
rect 18052 15623 18104 15632
rect 17684 15512 17736 15564
rect 18052 15589 18086 15623
rect 18086 15589 18104 15623
rect 18052 15580 18104 15589
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 14740 15444 14792 15453
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 17776 15487 17828 15496
rect 15936 15376 15988 15428
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 16764 15308 16816 15360
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 17960 15308 18012 15360
rect 18696 15308 18748 15360
rect 19340 15512 19392 15564
rect 19064 15444 19116 15496
rect 20444 15555 20496 15564
rect 20444 15521 20453 15555
rect 20453 15521 20487 15555
rect 20487 15521 20496 15555
rect 20444 15512 20496 15521
rect 20904 15555 20956 15564
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 19340 15376 19392 15428
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1952 15147 2004 15156
rect 1952 15113 1961 15147
rect 1961 15113 1995 15147
rect 1995 15113 2004 15147
rect 1952 15104 2004 15113
rect 4988 15104 5040 15156
rect 5540 15104 5592 15156
rect 6368 15104 6420 15156
rect 8208 15104 8260 15156
rect 9496 15104 9548 15156
rect 11796 15104 11848 15156
rect 11888 15104 11940 15156
rect 15752 15147 15804 15156
rect 3148 15036 3200 15088
rect 4068 15036 4120 15088
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 3976 14968 4028 15020
rect 7472 15036 7524 15088
rect 8944 15036 8996 15088
rect 10048 15036 10100 15088
rect 5264 14968 5316 15020
rect 2136 14943 2188 14952
rect 2136 14909 2145 14943
rect 2145 14909 2179 14943
rect 2179 14909 2188 14943
rect 2136 14900 2188 14909
rect 5724 14900 5776 14952
rect 6276 14943 6328 14952
rect 6276 14909 6285 14943
rect 6285 14909 6319 14943
rect 6319 14909 6328 14943
rect 6276 14900 6328 14909
rect 6460 14900 6512 14952
rect 7932 14968 7984 15020
rect 8484 14968 8536 15020
rect 10232 14968 10284 15020
rect 11152 14968 11204 15020
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 3148 14832 3200 14884
rect 5356 14832 5408 14884
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 5908 14807 5960 14816
rect 5908 14773 5917 14807
rect 5917 14773 5951 14807
rect 5951 14773 5960 14807
rect 5908 14764 5960 14773
rect 7012 14832 7064 14884
rect 10968 14900 11020 14952
rect 11888 14900 11940 14952
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 16120 15104 16172 15156
rect 16304 15104 16356 15156
rect 12256 14968 12308 15020
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 13544 14968 13596 15020
rect 15844 15036 15896 15088
rect 13636 14900 13688 14952
rect 17960 15036 18012 15088
rect 17224 14968 17276 15020
rect 17592 15011 17644 15020
rect 17592 14977 17601 15011
rect 17601 14977 17635 15011
rect 17635 14977 17644 15011
rect 17592 14968 17644 14977
rect 7932 14832 7984 14884
rect 12348 14832 12400 14884
rect 14096 14875 14148 14884
rect 6460 14764 6512 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 7748 14764 7800 14816
rect 8392 14764 8444 14816
rect 11888 14764 11940 14816
rect 12072 14764 12124 14816
rect 14096 14841 14130 14875
rect 14130 14841 14148 14875
rect 14096 14832 14148 14841
rect 14188 14832 14240 14884
rect 14648 14764 14700 14816
rect 16672 14900 16724 14952
rect 18696 14900 18748 14952
rect 19064 15147 19116 15156
rect 19064 15113 19073 15147
rect 19073 15113 19107 15147
rect 19107 15113 19116 15147
rect 21364 15147 21416 15156
rect 19064 15104 19116 15113
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 20444 14968 20496 15020
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 19064 14900 19116 14952
rect 19156 14900 19208 14952
rect 20628 14943 20680 14952
rect 20628 14909 20637 14943
rect 20637 14909 20671 14943
rect 20671 14909 20680 14943
rect 20628 14900 20680 14909
rect 15292 14764 15344 14816
rect 15384 14764 15436 14816
rect 18236 14832 18288 14884
rect 20720 14832 20772 14884
rect 20444 14764 20496 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2780 14560 2832 14612
rect 7288 14560 7340 14612
rect 8208 14560 8260 14612
rect 8392 14560 8444 14612
rect 10048 14560 10100 14612
rect 10508 14560 10560 14612
rect 1860 14424 1912 14476
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 4160 14424 4212 14476
rect 5264 14424 5316 14476
rect 2320 14356 2372 14408
rect 5540 14492 5592 14544
rect 7196 14424 7248 14476
rect 9128 14467 9180 14476
rect 9128 14433 9137 14467
rect 9137 14433 9171 14467
rect 9171 14433 9180 14467
rect 9128 14424 9180 14433
rect 9496 14424 9548 14476
rect 9772 14424 9824 14476
rect 10416 14492 10468 14544
rect 12440 14560 12492 14612
rect 19156 14560 19208 14612
rect 20628 14560 20680 14612
rect 21180 14560 21232 14612
rect 13544 14424 13596 14476
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 16580 14424 16632 14476
rect 16672 14467 16724 14476
rect 16672 14433 16681 14467
rect 16681 14433 16715 14467
rect 16715 14433 16724 14467
rect 16672 14424 16724 14433
rect 19432 14424 19484 14476
rect 19708 14424 19760 14476
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 5724 14220 5776 14272
rect 8208 14220 8260 14272
rect 10048 14220 10100 14272
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 10876 14288 10928 14340
rect 12072 14288 12124 14340
rect 13728 14356 13780 14408
rect 15292 14356 15344 14408
rect 12532 14220 12584 14272
rect 14096 14263 14148 14272
rect 14096 14229 14105 14263
rect 14105 14229 14139 14263
rect 14139 14229 14148 14263
rect 14096 14220 14148 14229
rect 14648 14220 14700 14272
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 18236 14399 18288 14408
rect 16304 14356 16356 14365
rect 16488 14288 16540 14340
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 19524 14356 19576 14408
rect 21180 14424 21232 14476
rect 19616 14220 19668 14272
rect 20444 14220 20496 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 4252 14016 4304 14068
rect 4804 14016 4856 14068
rect 5724 14016 5776 14068
rect 7012 14016 7064 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 5264 13880 5316 13932
rect 6828 13948 6880 14000
rect 8484 14016 8536 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 9128 14059 9180 14068
rect 9128 14025 9137 14059
rect 9137 14025 9171 14059
rect 9171 14025 9180 14059
rect 9128 14016 9180 14025
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 3332 13812 3384 13864
rect 4620 13812 4672 13864
rect 5908 13812 5960 13864
rect 7288 13812 7340 13864
rect 4712 13787 4764 13796
rect 4712 13753 4721 13787
rect 4721 13753 4755 13787
rect 4755 13753 4764 13787
rect 4712 13744 4764 13753
rect 8208 13812 8260 13864
rect 9680 13880 9732 13932
rect 10324 13880 10376 13932
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 8760 13812 8812 13864
rect 10416 13812 10468 13864
rect 10876 13855 10928 13864
rect 10876 13821 10885 13855
rect 10885 13821 10919 13855
rect 10919 13821 10928 13855
rect 10876 13812 10928 13821
rect 10048 13744 10100 13796
rect 12716 13812 12768 13864
rect 12900 13880 12952 13932
rect 14740 14016 14792 14068
rect 16488 14016 16540 14068
rect 17132 14016 17184 14068
rect 19524 14059 19576 14068
rect 19524 14025 19533 14059
rect 19533 14025 19567 14059
rect 19567 14025 19576 14059
rect 19524 14016 19576 14025
rect 21088 14059 21140 14068
rect 21088 14025 21097 14059
rect 21097 14025 21131 14059
rect 21131 14025 21140 14059
rect 21088 14016 21140 14025
rect 13544 13948 13596 14000
rect 16396 13948 16448 14000
rect 18052 13948 18104 14000
rect 19432 13991 19484 14000
rect 19432 13957 19441 13991
rect 19441 13957 19475 13991
rect 19475 13957 19484 13991
rect 19432 13948 19484 13957
rect 14096 13880 14148 13932
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 19156 13880 19208 13932
rect 20628 13948 20680 14000
rect 11152 13787 11204 13796
rect 11152 13753 11186 13787
rect 11186 13753 11204 13787
rect 11152 13744 11204 13753
rect 13912 13744 13964 13796
rect 14188 13812 14240 13864
rect 15660 13812 15712 13864
rect 15200 13744 15252 13796
rect 16396 13744 16448 13796
rect 16580 13787 16632 13796
rect 16580 13753 16589 13787
rect 16589 13753 16623 13787
rect 16623 13753 16632 13787
rect 16580 13744 16632 13753
rect 16672 13744 16724 13796
rect 19340 13812 19392 13864
rect 18144 13744 18196 13796
rect 19800 13744 19852 13796
rect 4804 13719 4856 13728
rect 4804 13685 4813 13719
rect 4813 13685 4847 13719
rect 4847 13685 4856 13719
rect 4804 13676 4856 13685
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 7380 13676 7432 13728
rect 8760 13676 8812 13728
rect 9772 13676 9824 13728
rect 12256 13719 12308 13728
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 13728 13676 13780 13728
rect 17132 13676 17184 13728
rect 19892 13719 19944 13728
rect 19892 13685 19901 13719
rect 19901 13685 19935 13719
rect 19935 13685 19944 13719
rect 19892 13676 19944 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 4160 13472 4212 13524
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 4712 13472 4764 13524
rect 4252 13447 4304 13456
rect 4252 13413 4261 13447
rect 4261 13413 4295 13447
rect 4295 13413 4304 13447
rect 4252 13404 4304 13413
rect 4804 13404 4856 13456
rect 2964 13336 3016 13388
rect 4344 13336 4396 13388
rect 6920 13472 6972 13524
rect 7196 13515 7248 13524
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 7380 13472 7432 13524
rect 7748 13472 7800 13524
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 9772 13515 9824 13524
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 10416 13472 10468 13524
rect 10968 13472 11020 13524
rect 14188 13515 14240 13524
rect 10048 13447 10100 13456
rect 1676 13268 1728 13320
rect 4344 13132 4396 13184
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 5908 13268 5960 13320
rect 10048 13413 10057 13447
rect 10057 13413 10091 13447
rect 10091 13413 10100 13447
rect 10048 13404 10100 13413
rect 10600 13404 10652 13456
rect 12072 13404 12124 13456
rect 7288 13268 7340 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 12440 13336 12492 13388
rect 14188 13481 14197 13515
rect 14197 13481 14231 13515
rect 14231 13481 14240 13515
rect 14188 13472 14240 13481
rect 14740 13472 14792 13524
rect 14004 13404 14056 13456
rect 15292 13404 15344 13456
rect 16672 13404 16724 13456
rect 17960 13404 18012 13456
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 21180 13447 21232 13456
rect 9220 13268 9272 13320
rect 11704 13268 11756 13320
rect 12348 13311 12400 13320
rect 12348 13277 12357 13311
rect 12357 13277 12391 13311
rect 12391 13277 12400 13311
rect 12348 13268 12400 13277
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 13452 13268 13504 13320
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 15292 13311 15344 13320
rect 14372 13268 14424 13277
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 17500 13336 17552 13388
rect 16580 13268 16632 13320
rect 17960 13268 18012 13320
rect 18788 13268 18840 13320
rect 19248 13268 19300 13320
rect 7656 13132 7708 13184
rect 10508 13132 10560 13184
rect 11888 13132 11940 13184
rect 13544 13132 13596 13184
rect 13728 13175 13780 13184
rect 13728 13141 13737 13175
rect 13737 13141 13771 13175
rect 13771 13141 13780 13175
rect 13728 13132 13780 13141
rect 14740 13132 14792 13184
rect 15108 13132 15160 13184
rect 18052 13200 18104 13252
rect 18696 13132 18748 13184
rect 19708 13200 19760 13252
rect 20812 13336 20864 13388
rect 21180 13413 21189 13447
rect 21189 13413 21223 13447
rect 21223 13413 21232 13447
rect 21180 13404 21232 13413
rect 20444 13268 20496 13320
rect 20628 13200 20680 13252
rect 20996 13132 21048 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1584 12928 1636 12980
rect 3700 12928 3752 12980
rect 4068 12928 4120 12980
rect 5172 12860 5224 12912
rect 5908 12903 5960 12912
rect 5908 12869 5917 12903
rect 5917 12869 5951 12903
rect 5951 12869 5960 12903
rect 5908 12860 5960 12869
rect 2504 12792 2556 12844
rect 3792 12792 3844 12844
rect 5264 12792 5316 12844
rect 6368 12792 6420 12844
rect 8116 12792 8168 12844
rect 11152 12928 11204 12980
rect 11704 12928 11756 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 13544 12928 13596 12980
rect 18788 12928 18840 12980
rect 18972 12928 19024 12980
rect 19248 12971 19300 12980
rect 19248 12937 19257 12971
rect 19257 12937 19291 12971
rect 19291 12937 19300 12971
rect 19248 12928 19300 12937
rect 19892 12928 19944 12980
rect 9956 12860 10008 12912
rect 2964 12724 3016 12776
rect 3056 12656 3108 12708
rect 6092 12656 6144 12708
rect 6276 12656 6328 12708
rect 7288 12656 7340 12708
rect 7564 12656 7616 12708
rect 8116 12656 8168 12708
rect 8760 12699 8812 12708
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 2688 12631 2740 12640
rect 2688 12597 2697 12631
rect 2697 12597 2731 12631
rect 2731 12597 2740 12631
rect 2688 12588 2740 12597
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 4896 12588 4948 12640
rect 8760 12665 8794 12699
rect 8794 12665 8812 12699
rect 8760 12656 8812 12665
rect 9128 12724 9180 12776
rect 9680 12724 9732 12776
rect 9772 12724 9824 12776
rect 13636 12860 13688 12912
rect 19708 12860 19760 12912
rect 11704 12792 11756 12844
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 13728 12792 13780 12844
rect 15108 12792 15160 12844
rect 15476 12792 15528 12844
rect 17500 12792 17552 12844
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 20444 12792 20496 12844
rect 20812 12792 20864 12844
rect 11796 12724 11848 12776
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 10968 12656 11020 12708
rect 10508 12588 10560 12640
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 14096 12588 14148 12640
rect 14740 12588 14792 12640
rect 17776 12724 17828 12776
rect 18972 12724 19024 12776
rect 18144 12656 18196 12708
rect 18052 12588 18104 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 18604 12588 18656 12640
rect 18880 12588 18932 12640
rect 19432 12588 19484 12640
rect 20076 12588 20128 12640
rect 20720 12656 20772 12708
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 2964 12427 3016 12436
rect 2964 12393 2973 12427
rect 2973 12393 3007 12427
rect 3007 12393 3016 12427
rect 2964 12384 3016 12393
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 3700 12384 3752 12436
rect 3792 12384 3844 12436
rect 4804 12384 4856 12436
rect 9128 12384 9180 12436
rect 9496 12384 9548 12436
rect 2504 12316 2556 12368
rect 5264 12316 5316 12368
rect 6736 12316 6788 12368
rect 7564 12316 7616 12368
rect 8484 12316 8536 12368
rect 8760 12316 8812 12368
rect 2228 12248 2280 12300
rect 3792 12248 3844 12300
rect 7288 12248 7340 12300
rect 9220 12248 9272 12300
rect 10508 12316 10560 12368
rect 10968 12316 11020 12368
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 2688 12180 2740 12232
rect 4528 12180 4580 12232
rect 3332 12112 3384 12164
rect 4804 12180 4856 12232
rect 8024 12180 8076 12232
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 6000 12112 6052 12164
rect 6828 12112 6880 12164
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 8484 12044 8536 12096
rect 9128 12044 9180 12096
rect 9772 12044 9824 12096
rect 10048 12044 10100 12096
rect 10232 12044 10284 12096
rect 10876 12248 10928 12300
rect 12808 12384 12860 12436
rect 13728 12384 13780 12436
rect 13820 12384 13872 12436
rect 16396 12384 16448 12436
rect 18420 12384 18472 12436
rect 19340 12427 19392 12436
rect 19340 12393 19349 12427
rect 19349 12393 19383 12427
rect 19383 12393 19392 12427
rect 19340 12384 19392 12393
rect 19708 12427 19760 12436
rect 19708 12393 19717 12427
rect 19717 12393 19751 12427
rect 19751 12393 19760 12427
rect 19708 12384 19760 12393
rect 20076 12384 20128 12436
rect 20260 12384 20312 12436
rect 14648 12316 14700 12368
rect 18696 12316 18748 12368
rect 12808 12291 12860 12300
rect 12808 12257 12842 12291
rect 12842 12257 12860 12291
rect 12808 12248 12860 12257
rect 13360 12248 13412 12300
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 16212 12248 16264 12300
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 17960 12291 18012 12300
rect 17960 12257 17969 12291
rect 17969 12257 18003 12291
rect 18003 12257 18012 12291
rect 17960 12248 18012 12257
rect 18052 12248 18104 12300
rect 12256 12180 12308 12232
rect 12440 12180 12492 12232
rect 15476 12180 15528 12232
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 14372 12044 14424 12096
rect 14924 12044 14976 12096
rect 15108 12044 15160 12096
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 16764 12044 16816 12096
rect 17500 12180 17552 12232
rect 17868 12180 17920 12232
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 19156 12223 19208 12232
rect 19156 12189 19165 12223
rect 19165 12189 19199 12223
rect 19199 12189 19208 12223
rect 19156 12180 19208 12189
rect 19156 12044 19208 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 1768 11840 1820 11892
rect 4068 11840 4120 11892
rect 5264 11815 5316 11824
rect 5264 11781 5273 11815
rect 5273 11781 5307 11815
rect 5307 11781 5316 11815
rect 5264 11772 5316 11781
rect 6092 11840 6144 11892
rect 9220 11840 9272 11892
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 9956 11840 10008 11892
rect 10048 11772 10100 11824
rect 2228 11704 2280 11756
rect 2504 11704 2556 11756
rect 6184 11704 6236 11756
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8944 11747 8996 11756
rect 8024 11704 8076 11713
rect 2136 11636 2188 11688
rect 4528 11636 4580 11688
rect 4160 11611 4212 11620
rect 4160 11577 4194 11611
rect 4194 11577 4212 11611
rect 4160 11568 4212 11577
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 2320 11500 2372 11509
rect 4344 11500 4396 11552
rect 7472 11636 7524 11688
rect 8484 11636 8536 11688
rect 8944 11713 8953 11747
rect 8953 11713 8987 11747
rect 8987 11713 8996 11747
rect 8944 11704 8996 11713
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 11060 11840 11112 11892
rect 11888 11840 11940 11892
rect 12900 11840 12952 11892
rect 14096 11840 14148 11892
rect 14188 11840 14240 11892
rect 14924 11840 14976 11892
rect 15660 11840 15712 11892
rect 16212 11840 16264 11892
rect 17868 11883 17920 11892
rect 11244 11772 11296 11824
rect 11796 11772 11848 11824
rect 12256 11772 12308 11824
rect 12992 11772 13044 11824
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 18604 11840 18656 11892
rect 19340 11840 19392 11892
rect 21272 11840 21324 11892
rect 12072 11747 12124 11756
rect 10784 11636 10836 11688
rect 7196 11568 7248 11620
rect 5080 11500 5132 11552
rect 6736 11500 6788 11552
rect 7748 11500 7800 11552
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 10508 11543 10560 11552
rect 10508 11509 10517 11543
rect 10517 11509 10551 11543
rect 10551 11509 10560 11543
rect 10508 11500 10560 11509
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 12348 11704 12400 11756
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 12440 11636 12492 11688
rect 13912 11636 13964 11688
rect 14740 11636 14792 11688
rect 19708 11772 19760 11824
rect 19800 11772 19852 11824
rect 18604 11704 18656 11756
rect 18788 11704 18840 11756
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 19156 11704 19208 11713
rect 19892 11747 19944 11756
rect 19892 11713 19901 11747
rect 19901 11713 19935 11747
rect 19935 11713 19944 11747
rect 19892 11704 19944 11713
rect 11244 11568 11296 11620
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 12164 11500 12216 11552
rect 12348 11500 12400 11552
rect 13728 11568 13780 11620
rect 16580 11636 16632 11688
rect 16764 11679 16816 11688
rect 16764 11645 16798 11679
rect 16798 11645 16816 11679
rect 16764 11636 16816 11645
rect 17316 11636 17368 11688
rect 20076 11636 20128 11688
rect 21548 11704 21600 11756
rect 17132 11568 17184 11620
rect 20720 11568 20772 11620
rect 13820 11500 13872 11552
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 16396 11500 16448 11552
rect 18696 11500 18748 11552
rect 18880 11543 18932 11552
rect 18880 11509 18889 11543
rect 18889 11509 18923 11543
rect 18923 11509 18932 11543
rect 18880 11500 18932 11509
rect 19708 11543 19760 11552
rect 19708 11509 19717 11543
rect 19717 11509 19751 11543
rect 19751 11509 19760 11543
rect 19708 11500 19760 11509
rect 20628 11500 20680 11552
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2504 11296 2556 11348
rect 3792 11296 3844 11348
rect 4068 11296 4120 11348
rect 4344 11296 4396 11348
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 4896 11296 4948 11348
rect 5080 11296 5132 11348
rect 6552 11296 6604 11348
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 13268 11296 13320 11348
rect 16948 11339 17000 11348
rect 16948 11305 16957 11339
rect 16957 11305 16991 11339
rect 16991 11305 17000 11339
rect 16948 11296 17000 11305
rect 2136 11228 2188 11280
rect 5540 11228 5592 11280
rect 7748 11228 7800 11280
rect 10140 11271 10192 11280
rect 10140 11237 10149 11271
rect 10149 11237 10183 11271
rect 10183 11237 10192 11271
rect 10140 11228 10192 11237
rect 10508 11228 10560 11280
rect 12992 11228 13044 11280
rect 17040 11228 17092 11280
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 2688 11160 2740 11212
rect 4344 11160 4396 11212
rect 3608 11135 3660 11144
rect 1584 11092 1636 11101
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 5264 11092 5316 11144
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 7380 11160 7432 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9312 11160 9364 11212
rect 10784 11160 10836 11212
rect 11244 11160 11296 11212
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 7104 11092 7156 11144
rect 8208 11092 8260 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 3792 10956 3844 11008
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 6736 11024 6788 11076
rect 6828 11024 6880 11076
rect 10140 11092 10192 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10692 11135 10744 11144
rect 10232 11092 10284 11101
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 13360 11160 13412 11212
rect 8668 10956 8720 11008
rect 10048 10956 10100 11008
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 13820 11092 13872 11144
rect 14372 11160 14424 11212
rect 14556 11160 14608 11212
rect 17868 11296 17920 11348
rect 18052 11296 18104 11348
rect 18972 11296 19024 11348
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 17224 11160 17276 11212
rect 15292 11092 15344 11144
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 16764 11092 16816 11144
rect 19064 11228 19116 11280
rect 19800 11228 19852 11280
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 17868 11092 17920 11144
rect 18972 11160 19024 11212
rect 19340 11160 19392 11212
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 20720 11296 20772 11348
rect 21364 11296 21416 11348
rect 20076 11228 20128 11280
rect 19432 11160 19484 11169
rect 20536 11160 20588 11212
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 19892 11092 19944 11144
rect 20444 11135 20496 11144
rect 20444 11101 20453 11135
rect 20453 11101 20487 11135
rect 20487 11101 20496 11135
rect 20444 11092 20496 11101
rect 12072 10956 12124 10965
rect 16580 10956 16632 11008
rect 17040 10956 17092 11008
rect 17592 10956 17644 11008
rect 18696 10956 18748 11008
rect 19064 10999 19116 11008
rect 19064 10965 19073 10999
rect 19073 10965 19107 10999
rect 19107 10965 19116 10999
rect 19064 10956 19116 10965
rect 19432 10956 19484 11008
rect 19892 10999 19944 11008
rect 19892 10965 19901 10999
rect 19901 10965 19935 10999
rect 19935 10965 19944 10999
rect 19892 10956 19944 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2320 10752 2372 10804
rect 3608 10752 3660 10804
rect 4344 10752 4396 10804
rect 5356 10752 5408 10804
rect 7012 10752 7064 10804
rect 8208 10752 8260 10804
rect 8944 10752 8996 10804
rect 2688 10659 2740 10668
rect 2688 10625 2697 10659
rect 2697 10625 2731 10659
rect 2731 10625 2740 10659
rect 2688 10616 2740 10625
rect 4160 10684 4212 10736
rect 9312 10727 9364 10736
rect 9312 10693 9321 10727
rect 9321 10693 9355 10727
rect 9355 10693 9364 10727
rect 9312 10684 9364 10693
rect 4344 10616 4396 10668
rect 5080 10616 5132 10668
rect 5448 10616 5500 10668
rect 11060 10752 11112 10804
rect 11796 10752 11848 10804
rect 12440 10795 12492 10804
rect 12440 10761 12449 10795
rect 12449 10761 12483 10795
rect 12483 10761 12492 10795
rect 12440 10752 12492 10761
rect 12900 10684 12952 10736
rect 16764 10727 16816 10736
rect 16764 10693 16773 10727
rect 16773 10693 16807 10727
rect 16807 10693 16816 10727
rect 16764 10684 16816 10693
rect 17960 10752 18012 10804
rect 18880 10752 18932 10804
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 18052 10684 18104 10736
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 10232 10616 10284 10668
rect 10692 10616 10744 10668
rect 3332 10548 3384 10600
rect 6920 10548 6972 10600
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 9220 10548 9272 10600
rect 12072 10548 12124 10600
rect 13820 10616 13872 10668
rect 14188 10616 14240 10668
rect 15568 10659 15620 10668
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 16672 10616 16724 10668
rect 17224 10616 17276 10668
rect 18144 10616 18196 10668
rect 19064 10659 19116 10668
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 19708 10616 19760 10668
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 20444 10616 20496 10668
rect 13176 10548 13228 10600
rect 15752 10548 15804 10600
rect 17960 10548 18012 10600
rect 19892 10548 19944 10600
rect 20812 10548 20864 10600
rect 21272 10591 21324 10600
rect 21272 10557 21281 10591
rect 21281 10557 21315 10591
rect 21315 10557 21324 10591
rect 21272 10548 21324 10557
rect 2504 10412 2556 10464
rect 2872 10455 2924 10464
rect 2872 10421 2881 10455
rect 2881 10421 2915 10455
rect 2915 10421 2924 10455
rect 2872 10412 2924 10421
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 5080 10480 5132 10532
rect 6184 10480 6236 10532
rect 8208 10480 8260 10532
rect 5172 10412 5224 10464
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 5724 10412 5776 10464
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 9864 10412 9916 10464
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 10508 10412 10560 10464
rect 11796 10412 11848 10464
rect 12164 10412 12216 10464
rect 14740 10412 14792 10464
rect 15660 10412 15712 10464
rect 20260 10480 20312 10532
rect 17776 10412 17828 10464
rect 18972 10412 19024 10464
rect 19064 10412 19116 10464
rect 19432 10412 19484 10464
rect 19616 10455 19668 10464
rect 19616 10421 19625 10455
rect 19625 10421 19659 10455
rect 19659 10421 19668 10455
rect 19616 10412 19668 10421
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 20076 10412 20128 10421
rect 20352 10412 20404 10464
rect 20720 10412 20772 10464
rect 20904 10455 20956 10464
rect 20904 10421 20913 10455
rect 20913 10421 20947 10455
rect 20947 10421 20956 10455
rect 20904 10412 20956 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2228 10208 2280 10260
rect 2872 10208 2924 10260
rect 2964 10208 3016 10260
rect 3976 10208 4028 10260
rect 5356 10251 5408 10260
rect 5356 10217 5365 10251
rect 5365 10217 5399 10251
rect 5399 10217 5408 10251
rect 5356 10208 5408 10217
rect 5448 10208 5500 10260
rect 8852 10208 8904 10260
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 10324 10208 10376 10260
rect 13176 10208 13228 10260
rect 14556 10208 14608 10260
rect 16212 10208 16264 10260
rect 16672 10251 16724 10260
rect 16672 10217 16681 10251
rect 16681 10217 16715 10251
rect 16715 10217 16724 10251
rect 16672 10208 16724 10217
rect 17592 10208 17644 10260
rect 2504 10140 2556 10192
rect 4160 10183 4212 10192
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 2872 10115 2924 10124
rect 2872 10081 2881 10115
rect 2881 10081 2915 10115
rect 2915 10081 2924 10115
rect 2872 10072 2924 10081
rect 4160 10149 4169 10183
rect 4169 10149 4203 10183
rect 4203 10149 4212 10183
rect 4160 10140 4212 10149
rect 5540 10140 5592 10192
rect 4804 10072 4856 10124
rect 12440 10140 12492 10192
rect 15568 10183 15620 10192
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 4160 10004 4212 10056
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 3976 9936 4028 9988
rect 6184 10072 6236 10124
rect 7564 10072 7616 10124
rect 2688 9868 2740 9920
rect 3240 9868 3292 9920
rect 7012 10004 7064 10056
rect 10048 10072 10100 10124
rect 10600 10072 10652 10124
rect 10876 10115 10928 10124
rect 10876 10081 10885 10115
rect 10885 10081 10919 10115
rect 10919 10081 10928 10115
rect 10876 10072 10928 10081
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 6644 9936 6696 9988
rect 6920 9868 6972 9920
rect 7012 9911 7064 9920
rect 7012 9877 7021 9911
rect 7021 9877 7055 9911
rect 7055 9877 7064 9911
rect 7288 9936 7340 9988
rect 7748 9936 7800 9988
rect 10508 10004 10560 10056
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 14372 10072 14424 10124
rect 9128 9936 9180 9988
rect 13820 10004 13872 10056
rect 15568 10149 15602 10183
rect 15602 10149 15620 10183
rect 15568 10140 15620 10149
rect 19616 10140 19668 10192
rect 20536 10183 20588 10192
rect 20536 10149 20545 10183
rect 20545 10149 20579 10183
rect 20579 10149 20588 10183
rect 20536 10140 20588 10149
rect 16580 10072 16632 10124
rect 16856 10072 16908 10124
rect 19156 10072 19208 10124
rect 19524 10072 19576 10124
rect 19708 10115 19760 10124
rect 19708 10081 19717 10115
rect 19717 10081 19751 10115
rect 19751 10081 19760 10115
rect 19708 10072 19760 10081
rect 20260 10115 20312 10124
rect 20260 10081 20269 10115
rect 20269 10081 20303 10115
rect 20303 10081 20312 10115
rect 20260 10072 20312 10081
rect 14188 9936 14240 9988
rect 18696 10004 18748 10056
rect 19340 10004 19392 10056
rect 20168 10004 20220 10056
rect 20904 10004 20956 10056
rect 15200 9936 15252 9988
rect 18880 9936 18932 9988
rect 7012 9868 7064 9877
rect 9496 9868 9548 9920
rect 12256 9868 12308 9920
rect 12440 9868 12492 9920
rect 13176 9868 13228 9920
rect 20904 9868 20956 9920
rect 21548 9911 21600 9920
rect 21548 9877 21557 9911
rect 21557 9877 21591 9911
rect 21591 9877 21600 9911
rect 21548 9868 21600 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 3148 9664 3200 9716
rect 6000 9664 6052 9716
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 2688 9571 2740 9580
rect 2688 9537 2697 9571
rect 2697 9537 2731 9571
rect 2731 9537 2740 9571
rect 2688 9528 2740 9537
rect 5724 9596 5776 9648
rect 6736 9596 6788 9648
rect 7380 9639 7432 9648
rect 7380 9605 7389 9639
rect 7389 9605 7423 9639
rect 7423 9605 7432 9639
rect 7380 9596 7432 9605
rect 2136 9460 2188 9512
rect 5080 9528 5132 9580
rect 7012 9528 7064 9580
rect 8208 9528 8260 9580
rect 4068 9460 4120 9512
rect 2872 9392 2924 9444
rect 3148 9435 3200 9444
rect 3148 9401 3182 9435
rect 3182 9401 3200 9435
rect 3148 9392 3200 9401
rect 4160 9392 4212 9444
rect 1952 9324 2004 9376
rect 2780 9324 2832 9376
rect 2964 9324 3016 9376
rect 7564 9392 7616 9444
rect 12164 9596 12216 9648
rect 15844 9664 15896 9716
rect 18052 9664 18104 9716
rect 20076 9707 20128 9716
rect 20076 9673 20085 9707
rect 20085 9673 20119 9707
rect 20119 9673 20128 9707
rect 20076 9664 20128 9673
rect 15660 9596 15712 9648
rect 16212 9596 16264 9648
rect 19432 9639 19484 9648
rect 19432 9605 19441 9639
rect 19441 9605 19475 9639
rect 19475 9605 19484 9639
rect 19432 9596 19484 9605
rect 20168 9596 20220 9648
rect 15476 9528 15528 9580
rect 15752 9528 15804 9580
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 11060 9392 11112 9444
rect 11152 9392 11204 9444
rect 12256 9392 12308 9444
rect 7656 9324 7708 9376
rect 8300 9324 8352 9376
rect 9956 9324 10008 9376
rect 10968 9324 11020 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 15844 9460 15896 9512
rect 19800 9528 19852 9580
rect 16488 9460 16540 9512
rect 17868 9460 17920 9512
rect 21272 9528 21324 9580
rect 20904 9503 20956 9512
rect 20904 9469 20913 9503
rect 20913 9469 20947 9503
rect 20947 9469 20956 9503
rect 20904 9460 20956 9469
rect 14740 9392 14792 9444
rect 16672 9435 16724 9444
rect 16672 9401 16681 9435
rect 16681 9401 16715 9435
rect 16715 9401 16724 9435
rect 16672 9392 16724 9401
rect 18512 9392 18564 9444
rect 19800 9392 19852 9444
rect 13820 9324 13872 9333
rect 15568 9324 15620 9376
rect 15752 9324 15804 9376
rect 17132 9367 17184 9376
rect 17132 9333 17141 9367
rect 17141 9333 17175 9367
rect 17175 9333 17184 9367
rect 17132 9324 17184 9333
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 18236 9324 18288 9376
rect 18972 9324 19024 9376
rect 20720 9324 20772 9376
rect 21548 9367 21600 9376
rect 21548 9333 21557 9367
rect 21557 9333 21591 9367
rect 21591 9333 21600 9367
rect 21548 9324 21600 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 2688 9120 2740 9172
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 6552 9120 6604 9172
rect 8392 9120 8444 9172
rect 8576 9120 8628 9172
rect 9404 9120 9456 9172
rect 10600 9120 10652 9172
rect 10968 9163 11020 9172
rect 10968 9129 10977 9163
rect 10977 9129 11011 9163
rect 11011 9129 11020 9163
rect 10968 9120 11020 9129
rect 11704 9120 11756 9172
rect 12900 9120 12952 9172
rect 14096 9120 14148 9172
rect 15200 9120 15252 9172
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 16580 9120 16632 9172
rect 16672 9120 16724 9172
rect 18236 9120 18288 9172
rect 18512 9163 18564 9172
rect 18512 9129 18521 9163
rect 18521 9129 18555 9163
rect 18555 9129 18564 9163
rect 18512 9120 18564 9129
rect 20996 9163 21048 9172
rect 20996 9129 21005 9163
rect 21005 9129 21039 9163
rect 21039 9129 21048 9163
rect 20996 9120 21048 9129
rect 1124 9052 1176 9104
rect 3332 9052 3384 9104
rect 3516 9095 3568 9104
rect 3516 9061 3525 9095
rect 3525 9061 3559 9095
rect 3559 9061 3568 9095
rect 3516 9052 3568 9061
rect 5080 9052 5132 9104
rect 6644 9052 6696 9104
rect 1860 8984 1912 9036
rect 2872 8984 2924 9036
rect 4344 8984 4396 9036
rect 6828 8984 6880 9036
rect 6184 8848 6236 8900
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 8484 8916 8536 8968
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 10324 8984 10376 9036
rect 8576 8916 8628 8925
rect 9956 8916 10008 8968
rect 9864 8848 9916 8900
rect 10692 9052 10744 9104
rect 10968 8984 11020 9036
rect 18696 9052 18748 9104
rect 19432 9052 19484 9104
rect 12440 8984 12492 9036
rect 11336 8916 11388 8968
rect 13268 8916 13320 8968
rect 3332 8780 3384 8832
rect 4160 8780 4212 8832
rect 4896 8780 4948 8832
rect 7288 8780 7340 8832
rect 7748 8780 7800 8832
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 10232 8780 10284 8832
rect 11704 8823 11756 8832
rect 11704 8789 11713 8823
rect 11713 8789 11747 8823
rect 11747 8789 11756 8823
rect 11704 8780 11756 8789
rect 12256 8780 12308 8832
rect 14740 8780 14792 8832
rect 15936 8984 15988 9036
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 17408 9027 17460 9036
rect 17408 8993 17442 9027
rect 17442 8993 17460 9027
rect 17408 8984 17460 8993
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 15752 8848 15804 8900
rect 16764 8848 16816 8900
rect 16948 8780 17000 8832
rect 17868 8780 17920 8832
rect 21180 8916 21232 8968
rect 20444 8848 20496 8900
rect 20628 8848 20680 8900
rect 18972 8780 19024 8832
rect 20352 8780 20404 8832
rect 21364 8780 21416 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 4068 8576 4120 8628
rect 9864 8619 9916 8628
rect 4344 8508 4396 8560
rect 6828 8551 6880 8560
rect 6828 8517 6837 8551
rect 6837 8517 6871 8551
rect 6871 8517 6880 8551
rect 6828 8508 6880 8517
rect 7196 8508 7248 8560
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 9956 8576 10008 8628
rect 11244 8576 11296 8628
rect 11704 8576 11756 8628
rect 12072 8576 12124 8628
rect 13268 8619 13320 8628
rect 13268 8585 13277 8619
rect 13277 8585 13311 8619
rect 13311 8585 13320 8619
rect 13268 8576 13320 8585
rect 18604 8576 18656 8628
rect 14648 8508 14700 8560
rect 19340 8576 19392 8628
rect 19708 8576 19760 8628
rect 20812 8619 20864 8628
rect 20812 8585 20821 8619
rect 20821 8585 20855 8619
rect 20855 8585 20864 8619
rect 20812 8576 20864 8585
rect 2872 8440 2924 8492
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 3792 8440 3844 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 3700 8372 3752 8424
rect 4712 8372 4764 8424
rect 6276 8440 6328 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 9772 8440 9824 8492
rect 2872 8304 2924 8356
rect 3332 8236 3384 8288
rect 4528 8304 4580 8356
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 4344 8236 4396 8288
rect 6368 8304 6420 8356
rect 7196 8347 7248 8356
rect 7196 8313 7205 8347
rect 7205 8313 7239 8347
rect 7239 8313 7248 8347
rect 7196 8304 7248 8313
rect 8208 8372 8260 8424
rect 8484 8372 8536 8424
rect 9404 8372 9456 8424
rect 10232 8415 10284 8424
rect 5724 8236 5776 8288
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 9956 8304 10008 8356
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 10140 8304 10192 8356
rect 17408 8440 17460 8492
rect 18328 8440 18380 8492
rect 11244 8372 11296 8424
rect 10968 8304 11020 8356
rect 18144 8372 18196 8424
rect 18236 8372 18288 8424
rect 19156 8372 19208 8424
rect 20352 8372 20404 8424
rect 21180 8415 21232 8424
rect 21180 8381 21189 8415
rect 21189 8381 21223 8415
rect 21223 8381 21232 8415
rect 21180 8372 21232 8381
rect 20996 8304 21048 8356
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 19064 8236 19116 8288
rect 20444 8236 20496 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 5080 8032 5132 8084
rect 6368 8032 6420 8084
rect 16672 8032 16724 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 1952 7828 2004 7880
rect 3792 7896 3844 7948
rect 6920 7964 6972 8016
rect 15384 7964 15436 8016
rect 20260 7964 20312 8016
rect 21088 7964 21140 8016
rect 4068 7828 4120 7880
rect 5448 7896 5500 7948
rect 6276 7896 6328 7948
rect 6644 7896 6696 7948
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 3976 7760 4028 7812
rect 8576 7896 8628 7948
rect 9312 7896 9364 7948
rect 18052 7896 18104 7948
rect 20536 7896 20588 7948
rect 20628 7896 20680 7948
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 16948 7871 17000 7880
rect 8024 7828 8076 7837
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 19156 7828 19208 7880
rect 3424 7692 3476 7744
rect 4344 7692 4396 7744
rect 18420 7760 18472 7812
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 16120 7692 16172 7744
rect 18972 7692 19024 7744
rect 19064 7735 19116 7744
rect 19064 7701 19073 7735
rect 19073 7701 19107 7735
rect 19107 7701 19116 7735
rect 19064 7692 19116 7701
rect 20260 7692 20312 7744
rect 21180 7692 21232 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 3700 7531 3752 7540
rect 3700 7497 3709 7531
rect 3709 7497 3743 7531
rect 3743 7497 3752 7531
rect 3700 7488 3752 7497
rect 5172 7488 5224 7540
rect 5356 7488 5408 7540
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 6184 7488 6236 7540
rect 8300 7488 8352 7540
rect 9312 7488 9364 7540
rect 20628 7531 20680 7540
rect 20628 7497 20637 7531
rect 20637 7497 20671 7531
rect 20671 7497 20680 7531
rect 20628 7488 20680 7497
rect 2964 7420 3016 7472
rect 3608 7420 3660 7472
rect 5448 7420 5500 7472
rect 20536 7463 20588 7472
rect 20536 7429 20545 7463
rect 20545 7429 20579 7463
rect 20579 7429 20588 7463
rect 20536 7420 20588 7429
rect 2780 7352 2832 7404
rect 3148 7352 3200 7404
rect 3792 7352 3844 7404
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 4804 7352 4856 7404
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 9404 7352 9456 7404
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 19892 7284 19944 7336
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 4252 7216 4304 7268
rect 2688 7148 2740 7157
rect 3608 7148 3660 7200
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 8300 7216 8352 7268
rect 20260 7216 20312 7268
rect 5172 7148 5224 7200
rect 5356 7148 5408 7200
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 6092 7148 6144 7157
rect 20628 7148 20680 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 4620 6944 4672 6996
rect 2320 6876 2372 6928
rect 4804 6876 4856 6928
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 4068 6808 4120 6860
rect 14740 6808 14792 6860
rect 20628 6808 20680 6860
rect 3884 6672 3936 6724
rect 4160 6672 4212 6724
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 9036 6740 9088 6792
rect 17960 6740 18012 6792
rect 6092 6672 6144 6724
rect 3608 6647 3660 6656
rect 3608 6613 3617 6647
rect 3617 6613 3651 6647
rect 3651 6613 3660 6647
rect 3608 6604 3660 6613
rect 4344 6604 4396 6656
rect 5172 6604 5224 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 3976 6400 4028 6452
rect 11888 6400 11940 6452
rect 20260 6443 20312 6452
rect 20260 6409 20269 6443
rect 20269 6409 20303 6443
rect 20303 6409 20312 6443
rect 20260 6400 20312 6409
rect 5264 6332 5316 6384
rect 9588 6332 9640 6384
rect 20536 6264 20588 6316
rect 3332 6060 3384 6112
rect 20536 6060 20588 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 5816 5312 5868 5364
rect 17960 5312 18012 5364
rect 4068 5244 4120 5296
rect 6460 5244 6512 5296
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 9588 3068 9640 3120
rect 4988 2932 5040 2984
rect 5632 2932 5684 2984
rect 16120 2932 16172 2984
rect 20720 2864 20772 2916
rect 11244 2796 11296 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 3332 1980 3384 2032
rect 4804 1980 4856 2032
rect 4068 1164 4120 1216
rect 7196 1164 7248 1216
<< metal2 >>
rect 202 22200 258 23000
rect 570 22200 626 23000
rect 1030 22200 1086 23000
rect 1398 22200 1454 23000
rect 1858 22200 1914 23000
rect 2318 22200 2374 23000
rect 2686 22200 2742 23000
rect 2778 22672 2834 22681
rect 2778 22607 2834 22616
rect 216 19242 244 22200
rect 204 19236 256 19242
rect 204 19178 256 19184
rect 584 16590 612 22200
rect 1044 18358 1072 22200
rect 1308 19236 1360 19242
rect 1308 19178 1360 19184
rect 1320 18970 1348 19178
rect 1308 18964 1360 18970
rect 1308 18906 1360 18912
rect 1032 18352 1084 18358
rect 1032 18294 1084 18300
rect 1412 18290 1440 22200
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1504 19922 1532 20198
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 572 16584 624 16590
rect 572 16526 624 16532
rect 1124 9104 1176 9110
rect 1124 9046 1176 9052
rect 1136 241 1164 9046
rect 1504 5817 1532 19858
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 18630 1624 19246
rect 1688 19009 1716 19654
rect 1872 19258 1900 22200
rect 2332 20942 2360 22200
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 2148 19922 2176 20198
rect 2240 19922 2268 20334
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 1950 19408 2006 19417
rect 1950 19343 2006 19352
rect 1780 19230 1900 19258
rect 1674 19000 1730 19009
rect 1780 18970 1808 19230
rect 1860 19168 1912 19174
rect 1858 19136 1860 19145
rect 1912 19136 1914 19145
rect 1858 19071 1914 19080
rect 1964 18970 1992 19343
rect 2042 19272 2098 19281
rect 2042 19207 2098 19216
rect 2056 19174 2084 19207
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 1674 18935 1730 18944
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1950 18864 2006 18873
rect 1768 18828 1820 18834
rect 1950 18799 2006 18808
rect 1768 18770 1820 18776
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1780 17814 1808 18770
rect 1964 18426 1992 18799
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1950 18048 2006 18057
rect 1950 17983 2006 17992
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1964 17338 1992 17983
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1950 17096 2006 17105
rect 1950 17031 2006 17040
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 16046 1808 16390
rect 1964 16250 1992 17031
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1950 16144 2006 16153
rect 1950 16079 2006 16088
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1964 15706 1992 16079
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 1950 15192 2006 15201
rect 1950 15127 1952 15136
rect 2004 15127 2006 15136
rect 1952 15098 2004 15104
rect 2148 14958 2176 15302
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 1950 14648 2006 14657
rect 1950 14583 1952 14592
rect 2004 14583 2006 14592
rect 1952 14554 2004 14560
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1872 13938 1900 14418
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 12986 1624 13806
rect 1676 13320 1728 13326
rect 2240 13297 2268 19858
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2332 18766 2360 19246
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2424 18193 2452 19654
rect 2596 19440 2648 19446
rect 2594 19408 2596 19417
rect 2648 19408 2650 19417
rect 2594 19343 2650 19352
rect 2700 18850 2728 22200
rect 2792 20058 2820 22607
rect 2962 22264 3018 22273
rect 2962 22199 3018 22208
rect 3146 22200 3202 23000
rect 3606 22200 3662 23000
rect 3974 22200 4030 23000
rect 4434 22200 4490 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6550 22200 6606 23000
rect 7010 22200 7066 23000
rect 7378 22200 7434 23000
rect 7838 22200 7894 23000
rect 8206 22200 8262 23000
rect 8666 22200 8722 23000
rect 9126 22200 9182 23000
rect 9494 22200 9550 23000
rect 9954 22200 10010 23000
rect 10414 22200 10470 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12070 22200 12126 23000
rect 12530 22200 12586 23000
rect 12898 22200 12954 23000
rect 13358 22200 13414 23000
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14646 22200 14702 23000
rect 15106 22200 15162 23000
rect 15474 22200 15530 23000
rect 15934 22200 15990 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17590 22200 17646 23000
rect 18050 22200 18106 23000
rect 18510 22200 18566 23000
rect 18878 22200 18934 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20166 22200 20222 23000
rect 20626 22200 20682 23000
rect 20994 22200 21050 23000
rect 21086 22264 21142 22273
rect 2870 20768 2926 20777
rect 2870 20703 2926 20712
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2778 19816 2834 19825
rect 2778 19751 2834 19760
rect 2792 19310 2820 19751
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2884 19174 2912 20703
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2976 18970 3004 22199
rect 3160 21842 3188 22200
rect 3160 21814 3372 21842
rect 3146 21720 3202 21729
rect 3146 21655 3202 21664
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 3068 19242 3096 20878
rect 3160 19514 3188 21655
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 3160 18970 3188 19246
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 2608 18822 2728 18850
rect 2504 18692 2556 18698
rect 2504 18634 2556 18640
rect 2410 18184 2466 18193
rect 2410 18119 2466 18128
rect 2516 18086 2544 18634
rect 2608 18290 2636 18822
rect 2686 18728 2742 18737
rect 2686 18663 2688 18672
rect 2740 18663 2742 18672
rect 2688 18634 2740 18640
rect 2780 18624 2832 18630
rect 2832 18572 2912 18578
rect 2780 18566 2912 18572
rect 2792 18550 2912 18566
rect 2778 18456 2834 18465
rect 2884 18426 2912 18550
rect 2778 18391 2834 18400
rect 2872 18420 2924 18426
rect 2596 18284 2648 18290
rect 2596 18226 2648 18232
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2332 17542 2360 18022
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2792 17354 2820 18391
rect 2872 18362 2924 18368
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2870 17504 2926 17513
rect 2870 17439 2926 17448
rect 2700 17338 2820 17354
rect 2688 17332 2820 17338
rect 2740 17326 2820 17332
rect 2688 17274 2740 17280
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2700 16522 2728 17138
rect 2792 16794 2820 17138
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2778 16552 2834 16561
rect 2688 16516 2740 16522
rect 2778 16487 2834 16496
rect 2688 16458 2740 16464
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 15026 2360 15982
rect 2792 15706 2820 16487
rect 2884 16250 2912 17439
rect 2976 17338 3004 18158
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2976 17202 3004 17274
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2976 16640 3004 17138
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3056 16652 3108 16658
rect 2976 16612 3056 16640
rect 3056 16594 3108 16600
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 3160 16046 3188 17070
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2778 15600 2834 15609
rect 2778 15535 2834 15544
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2792 14618 2820 15535
rect 3160 15094 3188 15982
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3148 14884 3200 14890
rect 3148 14826 3200 14832
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 13938 2360 14350
rect 2870 14240 2926 14249
rect 2870 14175 2926 14184
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2778 13832 2834 13841
rect 2778 13767 2834 13776
rect 1676 13262 1728 13268
rect 2226 13288 2282 13297
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1584 12232 1636 12238
rect 1688 12220 1716 13262
rect 2226 13223 2282 13232
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1636 12192 1716 12220
rect 1584 12174 1636 12180
rect 1596 11150 1624 12174
rect 1780 11898 1808 12582
rect 2516 12374 2544 12786
rect 2686 12744 2742 12753
rect 2686 12679 2742 12688
rect 2700 12646 2728 12679
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 2240 11762 2268 12242
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2148 11286 2176 11630
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 9897 1716 10066
rect 1674 9888 1730 9897
rect 1674 9823 1730 9832
rect 2148 9518 2176 11222
rect 2240 10266 2268 11494
rect 2332 10810 2360 11494
rect 2516 11354 2544 11698
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2700 11218 2728 12174
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2700 10674 2728 11154
rect 2688 10668 2740 10674
rect 2608 10628 2688 10656
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2516 10198 2544 10406
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2608 10062 2636 10628
rect 2688 10610 2740 10616
rect 2792 10282 2820 13767
rect 2884 10690 2912 14175
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2976 12782 3004 13330
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2976 12442 3004 12718
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3068 12442 3096 12650
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3160 12322 3188 14826
rect 3068 12294 3188 12322
rect 2884 10662 3004 10690
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2700 10254 2820 10282
rect 2884 10266 2912 10406
rect 2976 10266 3004 10662
rect 2872 10260 2924 10266
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2700 9926 2728 10254
rect 2872 10202 2924 10208
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2136 9512 2188 9518
rect 1872 9460 2136 9466
rect 1872 9454 2188 9460
rect 1872 9438 2176 9454
rect 1872 9042 1900 9438
rect 2148 9389 2176 9438
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1872 7868 1900 8978
rect 1964 8634 1992 9318
rect 2700 9178 2728 9522
rect 2884 9450 2912 10066
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2792 8634 2820 9318
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2884 8498 2912 8978
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 1952 7880 2004 7886
rect 1872 7840 1952 7868
rect 1952 7822 2004 7828
rect 1964 6866 1992 7822
rect 2884 7546 2912 8298
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2976 7478 3004 9318
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 2332 800 2360 6870
rect 2700 2553 2728 7142
rect 2686 2544 2742 2553
rect 2686 2479 2742 2488
rect 2792 1601 2820 7346
rect 3068 4457 3096 12294
rect 3252 11393 3280 19790
rect 3344 18154 3372 21814
rect 3620 20482 3648 22200
rect 3620 20454 3740 20482
rect 3606 20360 3662 20369
rect 3606 20295 3662 20304
rect 3424 19984 3476 19990
rect 3424 19926 3476 19932
rect 3436 19417 3464 19926
rect 3620 19514 3648 20295
rect 3608 19508 3660 19514
rect 3608 19450 3660 19456
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3436 18578 3464 19343
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 18698 3556 19246
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3436 18550 3556 18578
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3344 16046 3372 16390
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3344 12170 3372 13806
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3238 11384 3294 11393
rect 3238 11319 3294 11328
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10010 3372 10542
rect 3160 9982 3372 10010
rect 3160 9722 3188 9982
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 9178 3188 9386
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3252 9058 3280 9862
rect 3344 9110 3372 9982
rect 3436 9489 3464 18362
rect 3528 12481 3556 18550
rect 3514 12472 3570 12481
rect 3514 12407 3570 12416
rect 3620 11234 3648 18702
rect 3712 18086 3740 20454
rect 3988 19310 4016 22200
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 21146 4108 21247
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 4448 20890 4476 22200
rect 4816 21026 4844 22200
rect 4816 20998 5120 21026
rect 4448 20862 5028 20890
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3804 16130 3832 18906
rect 4080 17785 4108 19654
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4066 17776 4122 17785
rect 4066 17711 4122 17720
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 3988 16590 4016 17002
rect 4172 16776 4200 18158
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4080 16748 4200 16776
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3712 16102 3832 16130
rect 3712 12986 3740 16102
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3712 12442 3740 12922
rect 3804 12850 3832 15982
rect 3896 15978 3924 16526
rect 3988 16250 4016 16526
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12442 3832 12786
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3804 11354 3832 12242
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3620 11206 3740 11234
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3620 10810 3648 11086
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3514 9888 3570 9897
rect 3514 9823 3570 9832
rect 3422 9480 3478 9489
rect 3422 9415 3478 9424
rect 3528 9110 3556 9823
rect 3160 9030 3280 9058
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3160 7410 3188 9030
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8294 3372 8774
rect 3712 8514 3740 11206
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10441 3832 10950
rect 3790 10432 3846 10441
rect 3790 10367 3846 10376
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3620 8486 3740 8514
rect 3792 8492 3844 8498
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3436 8090 3464 8434
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3424 7744 3476 7750
rect 3620 7721 3648 8486
rect 3792 8434 3844 8440
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3424 7686 3476 7692
rect 3606 7712 3662 7721
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3344 4865 3372 6054
rect 3330 4856 3386 4865
rect 3330 4791 3386 4800
rect 3054 4448 3110 4457
rect 3054 4383 3110 4392
rect 3332 2032 3384 2038
rect 3330 2000 3332 2009
rect 3384 2000 3386 2009
rect 3330 1935 3386 1944
rect 2778 1592 2834 1601
rect 2778 1527 2834 1536
rect 1122 232 1178 241
rect 1122 167 1178 176
rect 2318 0 2374 800
rect 3436 649 3464 7686
rect 3606 7647 3662 7656
rect 3712 7546 3740 8366
rect 3804 7954 3832 8434
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3620 7206 3648 7414
rect 3804 7410 3832 7890
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 6662 3648 7142
rect 3896 6730 3924 15914
rect 3988 15026 4016 16186
rect 4080 16028 4108 16748
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16182 4200 16594
rect 4264 16250 4292 17614
rect 4356 16658 4384 19178
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4804 17536 4856 17542
rect 4802 17504 4804 17513
rect 4856 17504 4858 17513
rect 4421 17436 4717 17456
rect 4802 17439 4858 17448
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 4540 17066 4568 17206
rect 4528 17060 4580 17066
rect 4528 17002 4580 17008
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4160 16176 4212 16182
rect 4160 16118 4212 16124
rect 4356 16114 4384 16390
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4816 16114 4844 17002
rect 4908 16794 4936 18090
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4908 16046 4936 16390
rect 5000 16130 5028 20862
rect 5092 16946 5120 20998
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5184 17882 5212 18158
rect 5276 18034 5304 22200
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5460 18290 5488 18770
rect 5736 18426 5764 22200
rect 6000 18624 6052 18630
rect 5998 18592 6000 18601
rect 6052 18592 6054 18601
rect 5998 18527 6054 18536
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5276 18006 5672 18034
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 17134 5212 17614
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5092 16918 5488 16946
rect 5000 16102 5120 16130
rect 4896 16040 4948 16046
rect 4080 16000 4292 16028
rect 4264 15722 4292 16000
rect 4896 15982 4948 15988
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 4264 15694 4384 15722
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 11801 4016 14758
rect 4080 14482 4108 15030
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4172 13530 4200 14418
rect 4264 14074 4292 15506
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4080 12889 4108 12922
rect 4066 12880 4122 12889
rect 4066 12815 4122 12824
rect 4066 11928 4122 11937
rect 4066 11863 4068 11872
rect 4120 11863 4122 11872
rect 4068 11834 4120 11840
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10266 4016 10406
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3974 10024 4030 10033
rect 3974 9959 3976 9968
rect 4028 9959 4030 9968
rect 3976 9930 4028 9936
rect 4080 9874 4108 11290
rect 4172 10742 4200 11562
rect 4264 11014 4292 13398
rect 4356 13394 4384 15694
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4816 14074 4844 15438
rect 5000 15162 5028 15914
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 5092 15042 5120 16102
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15706 5212 15846
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5000 15014 5120 15042
rect 5264 15020 5316 15026
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4632 13530 4660 13806
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4724 13530 4752 13738
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4816 13462 4844 13670
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4356 11558 4384 13126
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4816 12442 4844 12582
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4526 12336 4582 12345
rect 4526 12271 4582 12280
rect 4540 12238 4568 12271
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4528 11688 4580 11694
rect 4816 11676 4844 12174
rect 4580 11648 4844 11676
rect 4528 11630 4580 11636
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11354 4384 11494
rect 4540 11354 4568 11630
rect 4908 11354 4936 12582
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4264 10656 4292 10950
rect 4356 10810 4384 11154
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4344 10668 4396 10674
rect 4264 10628 4344 10656
rect 4160 10192 4212 10198
rect 4158 10160 4160 10169
rect 4212 10160 4214 10169
rect 4158 10095 4214 10104
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3988 9846 4108 9874
rect 3988 8294 4016 9846
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 9081 4108 9454
rect 4172 9450 4200 9998
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4172 8838 4200 9386
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4066 8664 4122 8673
rect 4066 8599 4068 8608
rect 4120 8599 4122 8608
rect 4068 8570 4120 8576
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7177 4016 7754
rect 4080 7342 4108 7822
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3974 6760 4030 6769
rect 3884 6724 3936 6730
rect 3974 6695 4030 6704
rect 3884 6666 3936 6672
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 3505 3648 6598
rect 3988 6458 4016 6695
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 4080 6225 4108 6802
rect 4172 6730 4200 8774
rect 4264 7274 4292 10628
rect 4344 10610 4396 10616
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8566 4384 8978
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4356 7750 4384 8230
rect 4540 8090 4568 8298
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4724 7886 4752 8366
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4816 7410 4844 10066
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8498 4936 8774
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4632 7002 4660 7142
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4816 6934 4844 7346
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4068 5296 4120 5302
rect 4066 5264 4068 5273
rect 4120 5264 4122 5273
rect 4066 5199 4122 5208
rect 4172 3913 4200 6666
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4158 3904 4214 3913
rect 4158 3839 4214 3848
rect 3606 3496 3662 3505
rect 3606 3431 3662 3440
rect 4356 2961 4384 6598
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4342 2952 4398 2961
rect 4342 2887 4398 2896
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 2038 4844 6870
rect 5000 2990 5028 15014
rect 5264 14962 5316 14968
rect 5276 14482 5304 14962
rect 5368 14890 5396 15506
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5460 14770 5488 16918
rect 5552 16250 5580 17750
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 15162 5580 15438
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5368 14742 5488 14770
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 13938 5304 14418
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5276 13326 5304 13874
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11354 5120 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10538 5120 10610
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10062 5120 10474
rect 5184 10470 5212 12854
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5276 12374 5304 12786
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5276 11830 5304 12310
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 5276 11150 5304 11766
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5368 10996 5396 14742
rect 5552 14550 5580 15098
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5538 12472 5594 12481
rect 5538 12407 5594 12416
rect 5552 11286 5580 12407
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5276 10968 5396 10996
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10169 5212 10406
rect 5170 10160 5226 10169
rect 5170 10095 5226 10104
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9586 5120 9998
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5092 8090 5120 9046
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5184 7546 5212 10095
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 6662 5212 7142
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5276 6390 5304 10968
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5368 10266 5396 10746
rect 5460 10674 5488 11086
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10266 5488 10610
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 10198 5580 10406
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5368 7206 5396 7482
rect 5460 7478 5488 7890
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5460 6798 5488 7414
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5644 2990 5672 18006
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 6012 17338 6040 17682
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 6104 17218 6132 22200
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6380 19514 6408 21082
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6196 18329 6224 18566
rect 6182 18320 6238 18329
rect 6182 18255 6238 18264
rect 6472 17626 6500 18770
rect 6564 18290 6592 22200
rect 7024 19394 7052 22200
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7024 19366 7236 19394
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 6642 19136 6698 19145
rect 6642 19071 6698 19080
rect 6656 18834 6684 19071
rect 6840 18902 6868 19246
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6472 17598 6592 17626
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6012 17190 6132 17218
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5736 14278 5764 14894
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5736 14074 5764 14214
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5736 13938 5764 14010
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 9654 5764 10406
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 7546 5764 8230
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5828 5370 5856 16594
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5920 15502 5948 16526
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 13870 5948 14758
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5920 12918 5948 13262
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 6012 12170 6040 17190
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6196 16658 6224 17070
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6196 15706 6224 16594
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6288 15502 6316 16934
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6288 14958 6316 15438
rect 6380 15162 6408 17478
rect 6472 16658 6500 17478
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6472 14822 6500 14894
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6380 12850 6408 13330
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 6104 11898 6132 12650
rect 6288 12102 6316 12650
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10470 6040 11154
rect 6196 11150 6224 11698
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10538 6224 11086
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 9722 6040 10406
rect 6196 10130 6224 10474
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6196 7546 6224 8842
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6288 7954 6316 8434
rect 6380 8362 6408 8910
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6380 8090 6408 8298
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6380 7410 6408 8026
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6730 6132 7142
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 6472 5302 6500 14758
rect 6564 11354 6592 17598
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6656 9994 6684 18634
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6748 17746 6776 18022
rect 6840 17814 6868 18158
rect 6932 17882 6960 18158
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 7024 17066 7052 19246
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 7024 16658 7052 17002
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7116 16250 7144 17682
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6748 12374 6776 15302
rect 7024 14890 7052 15302
rect 7208 14906 7236 19366
rect 7300 18170 7328 20198
rect 7392 18465 7420 22200
rect 7852 20346 7880 22200
rect 7760 20318 7880 20346
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 18902 7604 19178
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7378 18456 7434 18465
rect 7378 18391 7434 18400
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7300 18142 7420 18170
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 17882 7328 18022
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7392 17626 7420 18142
rect 7300 17598 7420 17626
rect 7300 15008 7328 17598
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 16794 7420 17478
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7392 15570 7420 15982
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7392 15434 7420 15506
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7484 15094 7512 18226
rect 7576 17066 7604 18226
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7668 17882 7696 18022
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7576 16794 7604 17002
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7576 16114 7604 16730
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7576 15706 7604 15846
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7300 14980 7420 15008
rect 7012 14884 7064 14890
rect 7208 14878 7328 14906
rect 7012 14826 7064 14832
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14006 6868 14758
rect 7024 14074 7052 14826
rect 7300 14822 7328 14878
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14618 7328 14758
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 7208 13682 7236 14418
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7300 13870 7328 14350
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7392 13734 7420 14980
rect 7380 13728 7432 13734
rect 6932 13530 6960 13670
rect 7208 13654 7328 13682
rect 7380 13670 7432 13676
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11082 6776 11494
rect 6840 11082 6868 12106
rect 7208 11626 7236 13466
rect 7300 13326 7328 13654
rect 7392 13530 7420 13670
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7576 13274 7604 15506
rect 7760 14906 7788 20318
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 8128 18068 8156 18294
rect 8220 18170 8248 22200
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19174 8340 19654
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8298 19000 8354 19009
rect 8298 18935 8300 18944
rect 8352 18935 8354 18944
rect 8300 18906 8352 18912
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8312 18358 8340 18770
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8404 18290 8432 18770
rect 8496 18630 8524 19858
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8482 18320 8538 18329
rect 8392 18284 8444 18290
rect 8482 18255 8484 18264
rect 8392 18226 8444 18232
rect 8536 18255 8538 18264
rect 8484 18226 8536 18232
rect 8220 18142 8616 18170
rect 8392 18080 8444 18086
rect 8128 18040 8248 18068
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8220 17882 8248 18040
rect 8392 18022 8444 18028
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7852 17338 7880 17614
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8220 17066 8248 17818
rect 8404 17338 8432 18022
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8312 16726 8340 17274
rect 8496 17202 8524 17546
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8496 16114 8524 17138
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8220 15638 8248 15846
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8220 15434 8248 15574
rect 8496 15502 8524 16050
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7668 14878 7788 14906
rect 7944 14890 7972 14962
rect 7932 14884 7984 14890
rect 7668 13410 7696 14878
rect 7932 14826 7984 14832
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 13530 7788 14758
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8220 14618 8248 15098
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8404 14618 8432 14758
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8220 13870 8248 14214
rect 8496 14074 8524 14962
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7668 13382 7788 13410
rect 7576 13246 7696 13274
rect 7576 13138 7604 13246
rect 7668 13190 7696 13246
rect 7484 13110 7604 13138
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7300 12306 7328 12650
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6564 9178 6592 9658
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6656 9110 6684 9930
rect 6748 9654 6776 11018
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 9926 6960 10542
rect 7024 10062 7052 10746
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 7024 9586 7052 9862
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8566 6868 8978
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7954 6684 8230
rect 6918 8120 6974 8129
rect 6918 8055 6974 8064
rect 6932 8022 6960 8055
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6552 7880 6604 7886
rect 6550 7848 6552 7857
rect 6604 7848 6606 7857
rect 6550 7783 6606 7792
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 7116 4842 7144 11086
rect 7208 8566 7236 11562
rect 7300 10606 7328 12242
rect 7484 11694 7512 13110
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12374 7604 12650
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7760 11558 7788 13382
rect 8220 13326 8248 13806
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8128 12714 8156 12786
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8496 12374 8524 14010
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 11762 8064 12174
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8496 11694 8524 12038
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 11286 7788 11494
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7300 9994 7328 10542
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7392 9654 7420 11154
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8220 10810 8248 11086
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7576 9450 7604 10066
rect 7748 9988 7800 9994
rect 7668 9948 7748 9976
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7668 9382 7696 9948
rect 7748 9930 7800 9936
rect 8220 9586 8248 10474
rect 8390 10024 8446 10033
rect 8390 9959 8446 9968
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7656 9376 7708 9382
rect 8300 9376 8352 9382
rect 7656 9318 7708 9324
rect 8220 9336 8300 9364
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7208 8362 7236 8502
rect 7300 8498 7328 8774
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 6840 4814 7144 4842
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 6840 2666 6868 4814
rect 6840 2638 6960 2666
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 4080 1057 4108 1158
rect 4066 1048 4122 1057
rect 4066 983 4122 992
rect 6932 800 6960 2638
rect 7208 1222 7236 8298
rect 7760 7410 7788 8774
rect 8220 8430 8248 9336
rect 8300 9318 8352 9324
rect 8404 9178 8432 9959
rect 8588 9178 8616 18142
rect 8680 18086 8708 22200
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8864 18970 8892 20266
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8772 17898 8800 18634
rect 8680 17870 8800 17898
rect 8864 17882 8892 18702
rect 9034 18456 9090 18465
rect 9034 18391 9090 18400
rect 8852 17876 8904 17882
rect 8680 16697 8708 17870
rect 8852 17818 8904 17824
rect 8864 17270 8892 17818
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8760 16992 8812 16998
rect 8864 16980 8892 17206
rect 8812 16952 8892 16980
rect 8760 16934 8812 16940
rect 8666 16688 8722 16697
rect 8666 16623 8722 16632
rect 8680 11014 8708 16623
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8772 13870 8800 16390
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8864 15502 8892 15914
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 9048 15450 9076 18391
rect 9140 15858 9168 22200
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9232 20058 9260 20198
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9324 17882 9352 19654
rect 9416 19514 9444 19790
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9416 19310 9444 19450
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9416 18766 9444 19246
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9324 17338 9352 17818
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9324 16726 9352 17070
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9140 15830 9352 15858
rect 9048 15422 9260 15450
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8956 14074 8984 15030
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 13530 8800 13670
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8772 13297 8800 13466
rect 8758 13288 8814 13297
rect 8758 13223 8814 13232
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8772 12374 8800 12650
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8944 11756 8996 11762
rect 8864 11716 8944 11744
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8864 10266 8892 11716
rect 8944 11698 8996 11704
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8956 10810 8984 11154
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8496 8430 8524 8910
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 8024 7880 8076 7886
rect 8022 7848 8024 7857
rect 8220 7868 8248 8366
rect 8588 7954 8616 8910
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8076 7848 8248 7868
rect 8078 7840 8248 7848
rect 8022 7783 8078 7792
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8312 7274 8340 7482
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 9048 6798 9076 15302
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9140 14074 9168 14418
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9232 13326 9260 15422
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9128 12776 9180 12782
rect 9126 12744 9128 12753
rect 9180 12744 9182 12753
rect 9126 12679 9182 12688
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9140 12102 9168 12378
rect 9232 12306 9260 13262
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9232 11898 9260 12242
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11218 9352 15830
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9220 11144 9272 11150
rect 9126 11112 9182 11121
rect 9220 11086 9272 11092
rect 9126 11047 9182 11056
rect 9140 9994 9168 11047
rect 9232 10606 9260 11086
rect 9324 10742 9352 11154
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9232 10266 9260 10542
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9416 9330 9444 15642
rect 9508 15162 9536 22200
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9692 18834 9720 20470
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 18601 9628 18634
rect 9586 18592 9642 18601
rect 9586 18527 9642 18536
rect 9588 18352 9640 18358
rect 9640 18329 9720 18340
rect 9640 18320 9734 18329
rect 9640 18312 9678 18320
rect 9588 18294 9640 18300
rect 9678 18255 9734 18264
rect 9784 17678 9812 19790
rect 9968 19224 9996 22200
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 10060 19990 10088 20402
rect 10048 19984 10100 19990
rect 10048 19926 10100 19932
rect 10060 19514 10088 19926
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9968 19196 10272 19224
rect 10138 19136 10194 19145
rect 10138 19071 10194 19080
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9968 18358 9996 18702
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 10152 18290 10180 19071
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9772 17672 9824 17678
rect 9678 17640 9734 17649
rect 9772 17614 9824 17620
rect 9678 17575 9734 17584
rect 9692 17542 9720 17575
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17202 9720 17478
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16046 9720 16934
rect 9784 16658 9812 17614
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9876 16998 9904 17138
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9680 15904 9732 15910
rect 9784 15858 9812 16594
rect 9876 16590 9904 16730
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9968 16522 9996 17138
rect 10060 16998 10088 17274
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9876 15910 9904 16118
rect 9732 15852 9812 15858
rect 9680 15846 9812 15852
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9692 15830 9812 15846
rect 9692 15502 9720 15830
rect 9968 15570 9996 16458
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16046 10088 16390
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9508 14482 9536 15098
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9692 13938 9720 15438
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9692 13410 9720 13874
rect 9784 13734 9812 14418
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9784 13530 9812 13670
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9692 13382 9812 13410
rect 9784 12782 9812 13382
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9508 12209 9536 12378
rect 9494 12200 9550 12209
rect 9494 12135 9550 12144
rect 9692 11898 9720 12718
rect 9772 12232 9824 12238
rect 9770 12200 9772 12209
rect 9824 12200 9826 12209
rect 9770 12135 9826 12144
rect 9784 12102 9812 12135
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9586 11792 9642 11801
rect 9642 11750 9720 11778
rect 9586 11727 9642 11736
rect 9494 10024 9550 10033
rect 9494 9959 9550 9968
rect 9508 9926 9536 9959
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9692 9500 9720 11750
rect 9876 10470 9904 15302
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10060 14618 10088 15030
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 14074 10088 14214
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 13462 10088 13738
rect 10048 13456 10100 13462
rect 10046 13424 10048 13433
rect 10100 13424 10102 13433
rect 10046 13359 10102 13368
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9968 12345 9996 12854
rect 9954 12336 10010 12345
rect 9954 12271 10010 12280
rect 10152 12288 10180 18022
rect 10244 15026 10272 19196
rect 10428 18578 10456 22200
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10612 19514 10640 19858
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10612 18970 10640 19110
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10428 18550 10548 18578
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10322 17504 10378 17513
rect 10322 17439 10378 17448
rect 10336 16998 10364 17439
rect 10428 17202 10456 18362
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10324 16992 10376 16998
rect 10322 16960 10324 16969
rect 10376 16960 10378 16969
rect 10322 16895 10378 16904
rect 10336 15366 10364 16895
rect 10416 16584 10468 16590
rect 10414 16552 10416 16561
rect 10468 16552 10470 16561
rect 10414 16487 10470 16496
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10428 15366 10456 15914
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10520 14804 10548 18550
rect 10244 14776 10548 14804
rect 10244 12356 10272 14776
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10336 13938 10364 14350
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10428 13870 10456 14486
rect 10520 13938 10548 14554
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 13530 10456 13806
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10612 13462 10640 18770
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10520 12646 10548 13126
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10508 12368 10560 12374
rect 10244 12328 10508 12356
rect 10508 12310 10560 12316
rect 9968 11898 9996 12271
rect 10152 12260 10364 12288
rect 10048 12096 10100 12102
rect 10232 12096 10284 12102
rect 10100 12056 10180 12084
rect 10048 12038 10100 12044
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10048 11824 10100 11830
rect 10046 11792 10048 11801
rect 10100 11792 10102 11801
rect 10152 11762 10180 12056
rect 10232 12038 10284 12044
rect 10046 11727 10102 11736
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11014 10088 11494
rect 10138 11384 10194 11393
rect 10138 11319 10194 11328
rect 10152 11286 10180 11319
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10152 11150 10180 11222
rect 10244 11150 10272 12038
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10244 10674 10272 11086
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 10060 10130 10088 10610
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10244 10033 10272 10406
rect 10336 10266 10364 12260
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10520 11286 10548 11494
rect 10508 11280 10560 11286
rect 10704 11234 10732 17138
rect 10796 11694 10824 22200
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10888 18086 10916 19246
rect 11256 18986 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11716 19786 11744 22200
rect 12084 19938 12112 22200
rect 12544 20074 12572 22200
rect 11900 19910 12112 19938
rect 12452 20046 12572 20074
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 10980 18958 11284 18986
rect 11336 18964 11388 18970
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10888 17202 10916 17682
rect 10980 17218 11008 18958
rect 11336 18906 11388 18912
rect 11348 18850 11376 18906
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11164 18822 11376 18850
rect 11072 17882 11100 18770
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11060 17332 11112 17338
rect 11164 17320 11192 18822
rect 11336 18760 11388 18766
rect 11256 18720 11336 18748
rect 11256 18222 11284 18720
rect 11336 18702 11388 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11794 18592 11850 18601
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11716 18290 11744 18566
rect 11794 18527 11850 18536
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11244 18216 11296 18222
rect 11808 18193 11836 18527
rect 11244 18158 11296 18164
rect 11794 18184 11850 18193
rect 11256 17610 11284 18158
rect 11704 18148 11756 18154
rect 11794 18119 11850 18128
rect 11704 18090 11756 18096
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11716 17338 11744 18090
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11112 17292 11192 17320
rect 11704 17332 11756 17338
rect 11060 17274 11112 17280
rect 11704 17274 11756 17280
rect 10876 17196 10928 17202
rect 10980 17190 11100 17218
rect 10876 17138 10928 17144
rect 10874 15872 10930 15881
rect 10874 15807 10930 15816
rect 10888 15706 10916 15807
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10966 15056 11022 15065
rect 10966 14991 11022 15000
rect 10980 14958 11008 14991
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10888 13870 10916 14282
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10980 12714 11008 13466
rect 11072 12730 11100 17190
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11428 16992 11480 16998
rect 11256 16952 11428 16980
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11164 15434 11192 16526
rect 11256 16250 11284 16952
rect 11428 16934 11480 16940
rect 11716 16658 11744 17138
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11716 16250 11744 16594
rect 11808 16454 11836 18022
rect 11900 17184 11928 19910
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 11992 18970 12020 19790
rect 12084 19174 12112 19790
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12084 18834 12112 18906
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11992 18154 12020 18702
rect 11980 18148 12032 18154
rect 12032 18108 12112 18136
rect 11980 18090 12032 18096
rect 11980 17672 12032 17678
rect 11978 17640 11980 17649
rect 12032 17640 12034 17649
rect 11978 17575 12034 17584
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 17338 12020 17478
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11900 17156 12020 17184
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11808 16046 11836 16390
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 15502 11652 15846
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11164 15026 11192 15370
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11164 12986 11192 13738
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 10968 12708 11020 12714
rect 11072 12702 11192 12730
rect 10968 12650 11020 12656
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10888 11234 10916 12242
rect 10980 11393 11008 12310
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10966 11384 11022 11393
rect 10966 11319 11022 11328
rect 10508 11222 10560 11228
rect 10612 11206 10732 11234
rect 10796 11218 10916 11234
rect 10784 11212 10916 11218
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10336 10169 10364 10202
rect 10322 10160 10378 10169
rect 10322 10095 10378 10104
rect 10230 10024 10286 10033
rect 10230 9959 10286 9968
rect 9692 9472 9996 9500
rect 9968 9382 9996 9472
rect 9324 9302 9444 9330
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9324 7954 9352 9302
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9416 8430 9444 9114
rect 10336 9042 10364 10095
rect 10520 10062 10548 10406
rect 10612 10130 10640 11206
rect 10836 11206 10916 11212
rect 10784 11154 10836 11160
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10704 10674 10732 11086
rect 11072 10810 11100 11834
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10612 9178 10640 10066
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10704 9110 10732 10610
rect 10874 10160 10930 10169
rect 11164 10146 11192 12702
rect 11256 11830 11284 15438
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11716 15026 11744 15574
rect 11808 15162 11836 15574
rect 11900 15434 11928 17002
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11900 14958 11928 15098
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11716 12986 11744 13262
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11716 12850 11744 12922
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11808 12782 11836 13194
rect 11900 13190 11928 14758
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 12102 11836 12582
rect 11796 12096 11848 12102
rect 11992 12050 12020 17156
rect 12084 16794 12112 18108
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12084 16250 12112 16730
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 14822 12112 15982
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 14346 12112 14758
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 12084 12850 12112 13398
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11796 12038 11848 12044
rect 11900 12022 12020 12050
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11900 11898 11928 12022
rect 11888 11892 11940 11898
rect 12176 11880 12204 19722
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12360 18766 12388 19178
rect 12348 18760 12400 18766
rect 12268 18720 12348 18748
rect 12268 18358 12296 18720
rect 12348 18702 12400 18708
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12268 17066 12296 17274
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12348 16992 12400 16998
rect 12346 16960 12348 16969
rect 12400 16960 12402 16969
rect 12346 16895 12402 16904
rect 12254 15056 12310 15065
rect 12254 14991 12256 15000
rect 12308 14991 12310 15000
rect 12256 14962 12308 14968
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12360 13977 12388 14826
rect 12452 14618 12480 20046
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12544 18698 12572 19926
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12636 19310 12664 19654
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12912 18952 12940 22200
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 20058 13124 20198
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13084 19236 13136 19242
rect 13084 19178 13136 19184
rect 12820 18924 12940 18952
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17270 12756 17478
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12728 16046 12756 16458
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12530 14376 12586 14385
rect 12346 13968 12402 13977
rect 12346 13903 12402 13912
rect 12452 13841 12480 14350
rect 12530 14311 12586 14320
rect 12544 14278 12572 14311
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12820 13954 12848 18924
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12912 18290 12940 18770
rect 13096 18766 13124 19178
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 13004 17785 13032 18702
rect 12990 17776 13046 17785
rect 12990 17711 13046 17720
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 15026 12940 15302
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12820 13938 12940 13954
rect 12820 13932 12952 13938
rect 12820 13926 12900 13932
rect 12716 13864 12768 13870
rect 12254 13832 12310 13841
rect 12254 13767 12310 13776
rect 12438 13832 12494 13841
rect 12820 13852 12848 13926
rect 12900 13874 12952 13880
rect 12768 13824 12848 13852
rect 13004 13852 13032 17614
rect 13188 17202 13216 19654
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16658 13124 16934
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13004 13824 13216 13852
rect 12716 13806 12768 13812
rect 12438 13767 12494 13776
rect 12268 13734 12296 13767
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12360 12186 12388 13262
rect 12452 12345 12480 13330
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12438 12336 12494 12345
rect 12820 12306 12848 12378
rect 12438 12271 12494 12280
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12440 12232 12492 12238
rect 12360 12180 12440 12186
rect 12360 12174 12492 12180
rect 11888 11834 11940 11840
rect 11992 11852 12204 11880
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11796 11824 11848 11830
rect 11848 11772 11928 11778
rect 11796 11766 11928 11772
rect 11808 11750 11928 11766
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11256 11218 11284 11562
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 11257 11560 11494
rect 11518 11248 11574 11257
rect 11244 11212 11296 11218
rect 11518 11183 11574 11192
rect 11244 11154 11296 11160
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11808 10470 11836 10746
rect 11900 10713 11928 11750
rect 11886 10704 11942 10713
rect 11886 10639 11942 10648
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11164 10118 11284 10146
rect 10874 10095 10876 10104
rect 10928 10095 10930 10104
rect 10876 10066 10928 10072
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11058 9616 11114 9625
rect 11058 9551 11114 9560
rect 11072 9450 11100 9551
rect 11164 9450 11192 9998
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9178 11008 9318
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10980 9042 11008 9114
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8498 9812 8774
rect 9876 8634 9904 8842
rect 9968 8634 9996 8910
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 10244 8430 10272 8774
rect 9404 8424 9456 8430
rect 10232 8424 10284 8430
rect 9404 8366 9456 8372
rect 9968 8362 10180 8378
rect 10232 8366 10284 8372
rect 10980 8362 11008 8978
rect 11256 8634 11284 10118
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 8974 11376 9318
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11716 8838 11744 9114
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11716 8634 11744 8774
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11256 8430 11284 8570
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 9956 8356 10192 8362
rect 10008 8350 10140 8356
rect 9956 8298 10008 8304
rect 10140 8298 10192 8304
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9324 7546 9352 7890
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9416 7410 9444 7686
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11900 6458 11928 10639
rect 11992 10452 12020 11852
rect 12268 11830 12296 12174
rect 12360 12158 12480 12174
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12360 11762 12388 12158
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12084 11098 12112 11698
rect 12360 11558 12388 11698
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12176 11354 12204 11494
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12084 11070 12204 11098
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10606 12112 10950
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12176 10470 12204 11070
rect 12164 10464 12216 10470
rect 11992 10424 12112 10452
rect 12084 8634 12112 10424
rect 12164 10406 12216 10412
rect 12176 9654 12204 10406
rect 12256 9920 12308 9926
rect 12254 9888 12256 9897
rect 12308 9888 12310 9897
rect 12254 9823 12310 9832
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12360 9500 12388 11494
rect 12452 10810 12480 11630
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12912 10742 12940 11834
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 13004 11286 13032 11766
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 13188 10606 13216 13824
rect 13280 12209 13308 16390
rect 13372 12306 13400 22200
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13556 19417 13584 19722
rect 13542 19408 13598 19417
rect 13542 19343 13598 19352
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 16726 13492 17478
rect 13556 17338 13584 17546
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13556 16590 13584 17138
rect 13648 17066 13676 17546
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13740 16522 13768 17138
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13832 16454 13860 22200
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13924 18902 13952 19110
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13924 17882 13952 18362
rect 14108 18222 14136 20334
rect 14200 19145 14228 22200
rect 14660 20398 14688 22200
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 15120 20330 15148 22200
rect 14556 20324 14608 20330
rect 14556 20266 14608 20272
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 14568 20058 14596 20266
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15488 20058 15516 22200
rect 15948 20058 15976 22200
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 14384 19938 14412 19994
rect 14384 19910 14596 19938
rect 14568 19786 14596 19910
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14464 19712 14516 19718
rect 14384 19660 14464 19666
rect 14384 19654 14516 19660
rect 14384 19638 14504 19654
rect 14384 19514 14412 19638
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14384 19174 14412 19450
rect 14372 19168 14424 19174
rect 14186 19136 14242 19145
rect 14186 19071 14242 19080
rect 14292 19116 14372 19122
rect 14292 19110 14424 19116
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14292 19094 14412 19110
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14200 18222 14228 18770
rect 14292 18306 14320 19094
rect 14384 19045 14412 19094
rect 14476 18986 14504 19110
rect 14384 18958 14504 18986
rect 14384 18426 14412 18958
rect 14464 18896 14516 18902
rect 14464 18838 14516 18844
rect 14476 18426 14504 18838
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14292 18278 14412 18306
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13924 16998 13952 17818
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13924 16046 13952 16390
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 14292 15978 14320 16526
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 13728 15904 13780 15910
rect 14096 15904 14148 15910
rect 13728 15846 13780 15852
rect 14094 15872 14096 15881
rect 14148 15872 14150 15881
rect 13740 15570 13768 15846
rect 14094 15807 14150 15816
rect 14384 15586 14412 18278
rect 14476 17746 14504 18362
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14476 15706 14504 16934
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 13728 15564 13780 15570
rect 14384 15558 14504 15586
rect 13728 15506 13780 15512
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14482 13584 14962
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13556 14006 13584 14418
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12986 13492 13262
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13556 12986 13584 13126
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13648 12918 13676 14894
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13734 13768 14350
rect 14108 14278 14136 14826
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 13938 14136 14214
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14200 13870 14228 14826
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 13912 13796 13964 13802
rect 13964 13756 14044 13784
rect 13912 13738 13964 13744
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 14016 13462 14044 13756
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 13740 12850 13768 13126
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 12442 13768 12786
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12442 13860 12718
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13266 12200 13322 12209
rect 13266 12135 13322 12144
rect 13280 11354 13308 12135
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13372 11218 13400 12242
rect 13740 11626 13768 12378
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11694 13952 12038
rect 14016 11778 14044 13398
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14108 11898 14136 12582
rect 14200 11898 14228 13466
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14384 12102 14412 13262
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14016 11750 14136 11778
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13832 11150 13860 11494
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 10674 13860 11086
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13188 10266 13216 10542
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12440 10192 12492 10198
rect 12440 10134 12492 10140
rect 12452 10033 12480 10134
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12438 10024 12494 10033
rect 12438 9959 12494 9968
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9625 12480 9862
rect 12438 9616 12494 9625
rect 12438 9551 12494 9560
rect 12440 9512 12492 9518
rect 12360 9472 12440 9500
rect 12440 9454 12492 9460
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12268 8838 12296 9386
rect 12452 9042 12480 9454
rect 12912 9178 12940 10066
rect 13188 9926 13216 10202
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13832 9382 13860 9998
rect 14108 9625 14136 11750
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 9994 14228 10610
rect 14384 10130 14412 11154
rect 14476 11121 14504 15558
rect 14568 11218 14596 19722
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 15198 19408 15254 19417
rect 14936 19242 14964 19382
rect 15198 19343 15254 19352
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 15212 19174 15240 19343
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14646 19000 14702 19009
rect 14817 18992 15113 19012
rect 14646 18935 14702 18944
rect 14660 18834 14688 18935
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14660 14822 14688 16594
rect 14752 16454 14780 18158
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15304 17202 15332 19858
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15396 17882 15424 19110
rect 15580 18426 15608 19790
rect 16132 19514 16160 19858
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15856 18222 15884 18702
rect 16040 18426 16068 19314
rect 16316 19174 16344 22200
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16132 18970 16160 19110
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16118 18728 16174 18737
rect 16118 18663 16174 18672
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16040 18290 16068 18362
rect 16132 18329 16160 18663
rect 16118 18320 16174 18329
rect 16028 18284 16080 18290
rect 16118 18255 16174 18264
rect 16028 18226 16080 18232
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 17882 15792 18022
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15856 17678 15884 18158
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15488 17066 15516 17614
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14752 15502 14780 15914
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15212 15638 15240 16390
rect 15304 16250 15332 17002
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15580 16794 15608 16934
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 15764 15162 15792 15574
rect 15856 15502 15884 16526
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15948 15434 15976 15642
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 12374 14688 14214
rect 14752 14074 14780 14418
rect 15304 14414 15332 14758
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14752 13190 14780 13466
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12850 15148 13126
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14752 11694 14780 12582
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 14936 11898 14964 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14936 11540 14964 11834
rect 15120 11762 15148 12038
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14752 11512 14964 11540
rect 14752 11370 14780 11512
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14660 11342 14780 11370
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14462 11112 14518 11121
rect 14462 11047 14518 11056
rect 14554 10568 14610 10577
rect 14554 10503 14610 10512
rect 14568 10266 14596 10503
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14094 9616 14150 9625
rect 14094 9551 14150 9560
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 14108 9178 14136 9551
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 13280 8634 13308 8910
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 14660 8566 14688 11342
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9450 14780 10406
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15212 10146 15240 13738
rect 15304 13462 15332 14350
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15292 13320 15344 13326
rect 15396 13308 15424 14758
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13870 15700 14214
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15344 13280 15424 13308
rect 15292 13262 15344 13268
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15488 12238 15516 12786
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15476 12232 15528 12238
rect 15672 12209 15700 12242
rect 15476 12174 15528 12180
rect 15658 12200 15714 12209
rect 15658 12135 15714 12144
rect 15672 11898 15700 12135
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11150 15516 11494
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15304 10690 15332 11086
rect 15304 10662 15516 10690
rect 15212 10118 15424 10146
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15212 9178 15240 9930
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14752 6866 14780 8774
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15396 8022 15424 10118
rect 15488 9586 15516 10662
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 10198 15608 10610
rect 15752 10600 15804 10606
rect 15750 10568 15752 10577
rect 15804 10568 15806 10577
rect 15750 10503 15806 10512
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 9382 15608 10134
rect 15672 9654 15700 10406
rect 15856 9722 15884 15030
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 9489 15792 9522
rect 15844 9512 15896 9518
rect 15750 9480 15806 9489
rect 15844 9454 15896 9460
rect 15750 9415 15806 9424
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 9178 15792 9318
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15764 8906 15792 9114
rect 15856 8974 15884 9454
rect 15948 9042 15976 15370
rect 16316 15162 16344 16594
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15638 16436 16050
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 16132 7750 16160 15098
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16316 13938 16344 14350
rect 16500 14346 16528 17206
rect 16592 16726 16620 19858
rect 16776 19242 16804 22200
rect 17132 20392 17184 20398
rect 17132 20334 17184 20340
rect 17144 19378 17172 20334
rect 17236 20262 17264 22200
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17512 19990 17540 20334
rect 17604 20058 17632 22200
rect 18064 20534 18092 22200
rect 18524 20890 18552 22200
rect 18524 20862 18644 20890
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18616 20602 18644 20862
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18052 20528 18104 20534
rect 18052 20470 18104 20476
rect 18892 20058 18920 22200
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 17500 19984 17552 19990
rect 17500 19926 17552 19932
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 18064 19514 18092 19790
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17408 19304 17460 19310
rect 17868 19304 17920 19310
rect 17408 19246 17460 19252
rect 17682 19272 17738 19281
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16684 18154 16712 18702
rect 16776 18630 16804 18770
rect 16764 18624 16816 18630
rect 16816 18584 16896 18612
rect 16764 18566 16816 18572
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16684 16590 16712 18090
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16684 15978 16712 16526
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16684 15314 16712 15914
rect 16764 15360 16816 15366
rect 16684 15308 16764 15314
rect 16684 15302 16816 15308
rect 16684 15286 16804 15302
rect 16684 14958 16712 15286
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16684 14482 16712 14894
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16408 13802 16436 13942
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16224 12102 16252 12242
rect 16408 12102 16436 12378
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16224 11898 16252 12038
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16408 11558 16436 12038
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16224 9654 16252 10202
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16500 9518 16528 14010
rect 16592 13802 16620 14418
rect 16684 13802 16712 14418
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 11694 16620 13262
rect 16684 11801 16712 13398
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16670 11792 16726 11801
rect 16670 11727 16726 11736
rect 16776 11694 16804 12038
rect 16868 11801 16896 18584
rect 17052 17202 17080 19246
rect 17420 18902 17448 19246
rect 17868 19246 17920 19252
rect 17682 19207 17738 19216
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17512 18426 17540 18770
rect 17696 18465 17724 19207
rect 17880 18766 17908 19246
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17682 18456 17738 18465
rect 17500 18420 17552 18426
rect 17682 18391 17738 18400
rect 17500 18362 17552 18368
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17144 16697 17172 18294
rect 17512 18290 17540 18362
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17420 17542 17448 17750
rect 17512 17678 17540 18226
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17696 17814 17724 18022
rect 17972 17882 18000 19178
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18064 18426 18092 19110
rect 18616 18902 18644 19314
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17868 17536 17920 17542
rect 18064 17524 18092 18022
rect 18156 17785 18184 18566
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18142 17776 18198 17785
rect 18142 17711 18198 17720
rect 17920 17496 18092 17524
rect 17868 17478 17920 17484
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 17144 14074 17172 16623
rect 17314 16552 17370 16561
rect 17314 16487 17370 16496
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17236 15026 17264 16118
rect 17328 16046 17356 16487
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16854 11792 16910 11801
rect 16854 11727 16910 11736
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16764 11688 16816 11694
rect 16816 11636 16896 11642
rect 16764 11630 16896 11636
rect 16592 11014 16620 11630
rect 16776 11614 16896 11630
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10130 16620 10950
rect 16776 10742 16804 11086
rect 16868 11082 16896 11614
rect 16960 11354 16988 12242
rect 17144 11626 17172 13670
rect 17420 12345 17448 17478
rect 17880 17270 17908 17478
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18524 16794 18552 17070
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17512 15706 17540 16594
rect 17788 16046 17816 16662
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17512 15008 17540 15642
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17696 15366 17724 15506
rect 17788 15502 17816 15982
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17972 15366 18000 15846
rect 18064 15638 18092 16390
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18708 16250 18736 18362
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17592 15020 17644 15026
rect 17512 14980 17592 15008
rect 17592 14962 17644 14968
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 12850 17540 13330
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17406 12336 17462 12345
rect 17406 12271 17462 12280
rect 17512 12238 17540 12786
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 17052 11014 17080 11222
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16684 10266 16712 10610
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16500 9042 16528 9454
rect 16672 9444 16724 9450
rect 16592 9404 16672 9432
rect 16592 9178 16620 9404
rect 16672 9386 16724 9392
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16684 8090 16712 9114
rect 16762 8936 16818 8945
rect 16762 8871 16764 8880
rect 16816 8871 16818 8880
rect 16764 8842 16816 8848
rect 16868 8820 16896 10066
rect 17144 9382 17172 11562
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17236 10674 17264 11154
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17328 9489 17356 11630
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 11014 17632 11086
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10266 17632 10950
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17696 9489 17724 15302
rect 18064 15178 18092 15574
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 17972 15150 18092 15178
rect 17972 15094 18000 15150
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 18708 14958 18736 15302
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18248 14414 18276 14826
rect 18236 14408 18288 14414
rect 18064 14368 18236 14396
rect 18064 14006 18092 14368
rect 18236 14350 18288 14356
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18142 13832 18198 13841
rect 18142 13767 18144 13776
rect 18196 13767 18198 13776
rect 18144 13738 18196 13744
rect 18800 13569 18828 17750
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18786 13560 18842 13569
rect 18786 13495 18842 13504
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17972 13326 18000 13398
rect 18800 13326 18828 13495
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17788 10470 17816 12718
rect 18064 12646 18092 13194
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11898 17908 12174
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17880 11150 17908 11290
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17972 10810 18000 12242
rect 18064 11354 18092 12242
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 18052 10736 18104 10742
rect 17958 10704 18014 10713
rect 18052 10678 18104 10684
rect 17958 10639 18014 10648
rect 17972 10606 18000 10639
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17776 10464 17828 10470
rect 18064 10441 18092 10678
rect 18156 10674 18184 12650
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18432 12442 18460 12582
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18616 11898 18644 12582
rect 18708 12374 18736 13126
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18800 11762 18828 12922
rect 18892 12646 18920 15914
rect 18984 12986 19012 16934
rect 19076 16590 19104 20334
rect 19352 20074 19380 22200
rect 19720 20602 19748 22200
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19260 20046 19380 20074
rect 19260 19854 19288 20046
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19260 18426 19288 18838
rect 19352 18426 19380 19858
rect 19444 18970 19472 19858
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19536 19174 19564 19790
rect 19984 19304 20036 19310
rect 20180 19258 20208 22200
rect 20640 21434 20668 22200
rect 20718 21720 20774 21729
rect 20718 21655 20774 21664
rect 20456 21406 20668 21434
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 19310 20392 20198
rect 19984 19246 20036 19252
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19444 18204 19472 18702
rect 19260 18193 19472 18204
rect 19246 18184 19472 18193
rect 19302 18176 19472 18184
rect 19246 18119 19302 18128
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16726 19196 17070
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 19076 15502 19104 16526
rect 19260 16266 19288 16594
rect 19352 16454 19380 17002
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19260 16250 19472 16266
rect 19260 16244 19484 16250
rect 19260 16238 19432 16244
rect 19432 16186 19484 16192
rect 19536 16046 19564 19110
rect 19720 18698 19748 19178
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19720 18290 19748 18634
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19996 17814 20024 19246
rect 20088 19230 20208 19258
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20088 18737 20116 19230
rect 20456 18834 20484 21406
rect 20626 21312 20682 21321
rect 20626 21247 20682 21256
rect 20534 20768 20590 20777
rect 20534 20703 20590 20712
rect 20548 19786 20576 20703
rect 20640 20058 20668 21247
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20732 19514 20760 21655
rect 21008 19938 21036 22200
rect 21086 22199 21142 22208
rect 21454 22200 21510 23000
rect 21546 22672 21602 22681
rect 21546 22607 21602 22616
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20916 19910 21036 19938
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20074 18728 20130 18737
rect 20074 18663 20130 18672
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 20180 17542 20208 18770
rect 20732 18630 20760 19246
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 18086 20760 18158
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 19720 16794 19748 17478
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19168 15706 19196 15914
rect 19260 15706 19288 15914
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 15162 19104 15438
rect 19352 15434 19380 15506
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18984 12782 19012 12922
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 17776 10406 17828 10412
rect 18050 10432 18106 10441
rect 18050 10367 18106 10376
rect 17958 9752 18014 9761
rect 17958 9687 18014 9696
rect 18052 9716 18104 9722
rect 17868 9512 17920 9518
rect 17314 9480 17370 9489
rect 17314 9415 17370 9424
rect 17682 9480 17738 9489
rect 17868 9454 17920 9460
rect 17682 9415 17738 9424
rect 17328 9382 17356 9415
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 16948 8832 17000 8838
rect 16868 8792 16948 8820
rect 16948 8774 17000 8780
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16960 7886 16988 8774
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 9600 3126 9628 6326
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 11256 1442 11284 2790
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11256 1414 11560 1442
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 11532 800 11560 1414
rect 16132 800 16160 2926
rect 17144 2553 17172 9318
rect 17130 2544 17186 2553
rect 17130 2479 17186 2488
rect 17328 1601 17356 9318
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17420 8498 17448 8978
rect 17880 8838 17908 9454
rect 17972 9081 18000 9687
rect 18052 9658 18104 9664
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 18064 8922 18092 9658
rect 17972 8894 18092 8922
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17972 7857 18000 8894
rect 18156 8514 18184 10610
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 9178 18276 9318
rect 18524 9178 18552 9386
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18524 8820 18552 9114
rect 18616 8922 18644 11698
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18708 11098 18736 11494
rect 18699 11070 18736 11098
rect 18699 11014 18727 11070
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18786 10840 18842 10849
rect 18892 10810 18920 11494
rect 18984 11354 19012 12174
rect 19076 11393 19104 14894
rect 19168 14618 19196 14894
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19154 14376 19210 14385
rect 19154 14311 19210 14320
rect 19168 13938 19196 14311
rect 19352 13954 19380 15370
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19444 14006 19472 14418
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19536 14074 19564 14350
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19260 13926 19380 13954
rect 19432 14000 19484 14006
rect 19628 13977 19656 14214
rect 19432 13942 19484 13948
rect 19614 13968 19670 13977
rect 19260 13433 19288 13926
rect 19614 13903 19670 13912
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19246 13424 19302 13433
rect 19246 13359 19302 13368
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19260 12986 19288 13262
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19352 12442 19380 13806
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19444 12322 19472 12582
rect 19260 12294 19472 12322
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19168 12102 19196 12174
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11762 19196 12038
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19062 11384 19118 11393
rect 18972 11348 19024 11354
rect 19062 11319 19118 11328
rect 18972 11290 19024 11296
rect 19064 11280 19116 11286
rect 19062 11248 19064 11257
rect 19116 11248 19118 11257
rect 18972 11212 19024 11218
rect 19062 11183 19118 11192
rect 18972 11154 19024 11160
rect 18786 10775 18842 10784
rect 18880 10804 18932 10810
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18708 9110 18736 9998
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18616 8894 18736 8922
rect 18524 8792 18644 8820
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18616 8634 18644 8792
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18156 8486 18276 8514
rect 18248 8430 18276 8486
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 17958 7848 18014 7857
rect 17958 7783 18014 7792
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17972 5817 18000 6734
rect 18064 6225 18092 7890
rect 18050 6216 18106 6225
rect 18050 6151 18106 6160
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 4865 18000 5306
rect 18156 5273 18184 8366
rect 18340 8090 18368 8434
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18432 7818 18460 8230
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18708 6769 18736 8894
rect 18800 8673 18828 10775
rect 18880 10746 18932 10752
rect 18984 10713 19012 11154
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 18970 10704 19026 10713
rect 19076 10674 19104 10950
rect 19168 10826 19196 11698
rect 19260 10962 19288 12294
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19352 11218 19380 11834
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19338 11112 19394 11121
rect 19338 11047 19394 11056
rect 19352 10962 19380 11047
rect 19444 11014 19472 11154
rect 19260 10934 19380 10962
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19338 10840 19394 10849
rect 19168 10798 19338 10826
rect 19338 10775 19394 10784
rect 18970 10639 19026 10648
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 19338 10568 19394 10577
rect 19338 10503 19394 10512
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18892 8945 18920 9930
rect 18984 9382 19012 10406
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18878 8936 18934 8945
rect 18878 8871 18934 8880
rect 18786 8664 18842 8673
rect 18786 8599 18842 8608
rect 18694 6760 18750 6769
rect 18694 6695 18750 6704
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18142 5264 18198 5273
rect 18142 5199 18198 5208
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18892 3505 18920 8871
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 7834 19012 8774
rect 19076 8294 19104 10406
rect 19352 10146 19380 10503
rect 19444 10470 19472 10950
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19260 10118 19380 10146
rect 19536 10130 19564 11290
rect 19628 10554 19656 13903
rect 19720 13258 19748 14418
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 19708 12912 19760 12918
rect 19708 12854 19760 12860
rect 19720 12442 19748 12854
rect 19812 12850 19840 13738
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 12986 19932 13670
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19720 11558 19748 11766
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19812 11286 19840 11766
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19904 11150 19932 11698
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19706 10840 19762 10849
rect 19706 10775 19762 10784
rect 19720 10674 19748 10775
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19904 10606 19932 10950
rect 19892 10600 19944 10606
rect 19628 10526 19840 10554
rect 19892 10542 19944 10548
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19628 10198 19656 10406
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19524 10124 19576 10130
rect 19168 9625 19196 10066
rect 19154 9616 19210 9625
rect 19154 9551 19210 9560
rect 19168 8537 19196 9551
rect 19154 8528 19210 8537
rect 19154 8463 19210 8472
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19168 8004 19196 8366
rect 19260 8129 19288 10118
rect 19524 10066 19576 10072
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19352 8634 19380 9998
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19444 9110 19472 9590
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19720 8634 19748 10066
rect 19812 9586 19840 10526
rect 19996 9636 20024 15982
rect 20180 13297 20208 17478
rect 20272 16028 20300 17682
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20364 16658 20392 17614
rect 20548 17610 20576 18022
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20626 17504 20682 17513
rect 20626 17439 20682 17448
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20364 16182 20392 16594
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20272 16000 20392 16028
rect 20166 13288 20222 13297
rect 20166 13223 20222 13232
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 12442 20116 12582
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20088 11286 20116 11630
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 20168 10668 20220 10674
rect 20272 10656 20300 12378
rect 20364 12209 20392 16000
rect 20548 15910 20576 17002
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20456 15026 20484 15506
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14278 20484 14758
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20442 13560 20498 13569
rect 20442 13495 20444 13504
rect 20496 13495 20498 13504
rect 20444 13466 20496 13472
rect 20444 13320 20496 13326
rect 20548 13297 20576 15846
rect 20640 15706 20668 17439
rect 20732 17270 20760 18022
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14618 20668 14894
rect 20732 14890 20760 17070
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20444 13262 20496 13268
rect 20534 13288 20590 13297
rect 20456 12850 20484 13262
rect 20640 13258 20668 13942
rect 20824 13546 20852 19858
rect 20916 19281 20944 19910
rect 20994 19816 21050 19825
rect 20994 19751 21050 19760
rect 21008 19514 21036 19751
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20902 19272 20958 19281
rect 20902 19207 20958 19216
rect 21100 18970 21128 22199
rect 21468 20482 21496 22200
rect 21284 20454 21496 20482
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 19922 21220 20198
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21178 19408 21234 19417
rect 21178 19343 21234 19352
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20994 18864 21050 18873
rect 20904 18828 20956 18834
rect 20994 18799 21050 18808
rect 20904 18770 20956 18776
rect 20916 18154 20944 18770
rect 21008 18426 21036 18799
rect 21086 18456 21142 18465
rect 20996 18420 21048 18426
rect 21086 18391 21142 18400
rect 20996 18362 21048 18368
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20994 18048 21050 18057
rect 20994 17983 21050 17992
rect 21008 17338 21036 17983
rect 21100 17882 21128 18391
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21100 17218 21128 17478
rect 21008 17190 21128 17218
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16658 20944 16934
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20916 15026 20944 15506
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20824 13518 20944 13546
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20534 13223 20590 13232
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20824 12850 20852 13330
rect 20916 12866 20944 13518
rect 21008 13190 21036 17190
rect 21086 17096 21142 17105
rect 21086 17031 21142 17040
rect 21100 16794 21128 17031
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21100 15609 21128 15642
rect 21086 15600 21142 15609
rect 21086 15535 21142 15544
rect 21086 14648 21142 14657
rect 21192 14618 21220 19343
rect 21284 18329 21312 20454
rect 21362 20360 21418 20369
rect 21362 20295 21418 20304
rect 21376 19514 21404 20295
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21270 18320 21326 18329
rect 21270 18255 21326 18264
rect 21376 17542 21404 18770
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21270 16552 21326 16561
rect 21270 16487 21326 16496
rect 21284 16250 21312 16487
rect 21272 16244 21324 16250
rect 21468 16232 21496 19858
rect 21560 18970 21588 22607
rect 21914 22200 21970 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 21928 19009 21956 22200
rect 22296 19718 22324 22200
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22756 19145 22784 22200
rect 22742 19136 22798 19145
rect 22742 19071 22798 19080
rect 21914 19000 21970 19009
rect 21548 18964 21600 18970
rect 21914 18935 21970 18944
rect 21548 18906 21600 18912
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21468 16204 21588 16232
rect 21272 16186 21324 16192
rect 21454 16144 21510 16153
rect 21454 16079 21510 16088
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21086 14583 21142 14592
rect 21180 14612 21232 14618
rect 21100 14074 21128 14583
rect 21180 14554 21232 14560
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21192 13462 21220 14418
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20812 12844 20864 12850
rect 20916 12838 21128 12866
rect 20812 12786 20864 12792
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20350 12200 20406 12209
rect 20350 12135 20406 12144
rect 20732 11626 20760 12650
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20456 10674 20484 11086
rect 20444 10668 20496 10674
rect 20272 10628 20392 10656
rect 20168 10610 20220 10616
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20088 9722 20116 10406
rect 20180 10062 20208 10610
rect 20260 10532 20312 10538
rect 20260 10474 20312 10480
rect 20272 10130 20300 10474
rect 20364 10470 20392 10628
rect 20444 10610 20496 10616
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20548 10198 20576 11154
rect 20536 10192 20588 10198
rect 20536 10134 20588 10140
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 20180 9654 20208 9998
rect 19904 9608 20024 9636
rect 20168 9648 20220 9654
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19812 9450 19840 9522
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19246 8120 19302 8129
rect 19246 8055 19302 8064
rect 19168 7976 19288 8004
rect 19156 7880 19208 7886
rect 18984 7828 19156 7834
rect 18984 7822 19208 7828
rect 18984 7806 19196 7822
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 18984 7177 19012 7686
rect 18970 7168 19026 7177
rect 18970 7103 19026 7112
rect 18878 3496 18934 3505
rect 18878 3431 18934 3440
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 17314 1592 17370 1601
rect 17314 1527 17370 1536
rect 19076 1057 19104 7686
rect 19168 7410 19196 7806
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19062 1048 19118 1057
rect 19062 983 19118 992
rect 3422 640 3478 649
rect 3422 575 3478 584
rect 6918 0 6974 800
rect 11518 0 11574 800
rect 16118 0 16174 800
rect 19260 241 19288 7976
rect 19904 7342 19932 9608
rect 20168 9590 20220 9596
rect 20640 8906 20668 11494
rect 20732 11354 20760 11562
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 9382 20760 10406
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20364 8430 20392 8774
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20272 7750 20300 7958
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20272 6458 20300 7210
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20364 2009 20392 8366
rect 20456 8294 20484 8842
rect 20824 8634 20852 10542
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20916 10062 20944 10406
rect 20994 10160 21050 10169
rect 20994 10095 21050 10104
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20916 9518 20944 9862
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 21008 9178 21036 10095
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 21008 8362 21036 9114
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 2961 20484 8230
rect 21100 8022 21128 12838
rect 21284 11898 21312 15846
rect 21468 15706 21496 16079
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21362 15192 21418 15201
rect 21362 15127 21364 15136
rect 21416 15127 21418 15136
rect 21364 15098 21416 15104
rect 21362 14240 21418 14249
rect 21362 14175 21418 14184
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21284 11234 21312 11494
rect 21376 11354 21404 14175
rect 21454 13832 21510 13841
rect 21454 13767 21510 13776
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21284 11206 21404 11234
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21284 9586 21312 10542
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21192 8430 21220 8910
rect 21376 8838 21404 11206
rect 21468 10810 21496 13767
rect 21560 11762 21588 16204
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21744 10169 21772 18566
rect 21730 10160 21786 10169
rect 21730 10095 21786 10104
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21560 9382 21588 9862
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20548 7478 20576 7890
rect 20640 7546 20668 7890
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20548 6322 20576 7414
rect 21192 7410 21220 7686
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 6866 20668 7142
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 4457 20576 6054
rect 20534 4448 20590 4457
rect 20534 4383 20590 4392
rect 21560 3913 21588 9318
rect 21546 3904 21602 3913
rect 21546 3839 21602 3848
rect 20442 2952 20498 2961
rect 20442 2887 20498 2896
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20350 2000 20406 2009
rect 20350 1935 20406 1944
rect 20732 800 20760 2858
rect 19246 232 19302 241
rect 19246 167 19302 176
rect 20718 0 20774 800
<< via2 >>
rect 2778 22616 2834 22672
rect 1950 19352 2006 19408
rect 1674 18944 1730 19000
rect 1858 19116 1860 19136
rect 1860 19116 1912 19136
rect 1912 19116 1914 19136
rect 1858 19080 1914 19116
rect 2042 19216 2098 19272
rect 1950 18808 2006 18864
rect 1950 17992 2006 18048
rect 1950 17040 2006 17096
rect 1950 16088 2006 16144
rect 1950 15156 2006 15192
rect 1950 15136 1952 15156
rect 1952 15136 2004 15156
rect 2004 15136 2006 15156
rect 1950 14612 2006 14648
rect 1950 14592 1952 14612
rect 1952 14592 2004 14612
rect 2004 14592 2006 14612
rect 2594 19388 2596 19408
rect 2596 19388 2648 19408
rect 2648 19388 2650 19408
rect 2594 19352 2650 19388
rect 2962 22208 3018 22264
rect 21086 22208 21142 22264
rect 2870 20712 2926 20768
rect 2778 19760 2834 19816
rect 3146 21664 3202 21720
rect 2410 18128 2466 18184
rect 2686 18692 2742 18728
rect 2686 18672 2688 18692
rect 2688 18672 2740 18692
rect 2740 18672 2742 18692
rect 2778 18400 2834 18456
rect 2870 17448 2926 17504
rect 2778 16496 2834 16552
rect 2778 15544 2834 15600
rect 2870 14184 2926 14240
rect 2778 13776 2834 13832
rect 2226 13232 2282 13288
rect 2686 12688 2742 12744
rect 1674 9832 1730 9888
rect 1490 5752 1546 5808
rect 2686 2488 2742 2544
rect 3606 20304 3662 20360
rect 3422 19352 3478 19408
rect 3238 11328 3294 11384
rect 3514 12416 3570 12472
rect 4066 21256 4122 21312
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4066 17720 4122 17776
rect 3514 9832 3570 9888
rect 3422 9424 3478 9480
rect 3790 10376 3846 10432
rect 3330 4800 3386 4856
rect 3054 4392 3110 4448
rect 3330 1980 3332 2000
rect 3332 1980 3384 2000
rect 3384 1980 3386 2000
rect 3330 1944 3386 1980
rect 2778 1536 2834 1592
rect 1122 176 1178 232
rect 3606 7656 3662 7712
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4802 17484 4804 17504
rect 4804 17484 4856 17504
rect 4856 17484 4858 17504
rect 4802 17448 4858 17484
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 5998 18572 6000 18592
rect 6000 18572 6052 18592
rect 6052 18572 6054 18592
rect 5998 18536 6054 18572
rect 4066 12824 4122 12880
rect 4066 11892 4122 11928
rect 4066 11872 4068 11892
rect 4068 11872 4120 11892
rect 4120 11872 4122 11892
rect 3974 11736 4030 11792
rect 3974 9988 4030 10024
rect 3974 9968 3976 9988
rect 3976 9968 4028 9988
rect 4028 9968 4030 9988
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4526 12280 4582 12336
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4158 10140 4160 10160
rect 4160 10140 4212 10160
rect 4212 10140 4214 10160
rect 4158 10104 4214 10140
rect 4066 9016 4122 9072
rect 4066 8628 4122 8664
rect 4066 8608 4068 8628
rect 4068 8608 4120 8628
rect 4120 8608 4122 8628
rect 3974 7112 4030 7168
rect 3974 6704 4030 6760
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4066 6160 4122 6216
rect 4066 5244 4068 5264
rect 4068 5244 4120 5264
rect 4120 5244 4122 5264
rect 4066 5208 4122 5244
rect 4158 3848 4214 3904
rect 3606 3440 3662 3496
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4342 2896 4398 2952
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5538 12416 5594 12472
rect 5170 10104 5226 10160
rect 6182 18264 6238 18320
rect 6642 19080 6698 19136
rect 7378 18400 7434 18456
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 8298 18964 8354 19000
rect 8298 18944 8300 18964
rect 8300 18944 8352 18964
rect 8352 18944 8354 18964
rect 8482 18284 8538 18320
rect 8482 18264 8484 18284
rect 8484 18264 8536 18284
rect 8536 18264 8538 18284
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 6918 8064 6974 8120
rect 6550 7828 6552 7848
rect 6552 7828 6604 7848
rect 6604 7828 6606 7848
rect 6550 7792 6606 7828
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 8390 9968 8446 10024
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 4066 992 4122 1048
rect 9034 18400 9090 18456
rect 8666 16632 8722 16688
rect 8758 13232 8814 13288
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 8022 7828 8024 7848
rect 8024 7828 8076 7848
rect 8076 7828 8078 7848
rect 8022 7792 8078 7828
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 9126 12724 9128 12744
rect 9128 12724 9180 12744
rect 9180 12724 9182 12744
rect 9126 12688 9182 12724
rect 9126 11056 9182 11112
rect 9586 18536 9642 18592
rect 9678 18264 9734 18320
rect 10138 19080 10194 19136
rect 9678 17584 9734 17640
rect 9494 12144 9550 12200
rect 9770 12180 9772 12200
rect 9772 12180 9824 12200
rect 9824 12180 9826 12200
rect 9770 12144 9826 12180
rect 9586 11736 9642 11792
rect 9494 9968 9550 10024
rect 10046 13404 10048 13424
rect 10048 13404 10100 13424
rect 10100 13404 10102 13424
rect 10046 13368 10102 13404
rect 9954 12280 10010 12336
rect 10322 17448 10378 17504
rect 10322 16940 10324 16960
rect 10324 16940 10376 16960
rect 10376 16940 10378 16960
rect 10322 16904 10378 16940
rect 10414 16532 10416 16552
rect 10416 16532 10468 16552
rect 10468 16532 10470 16552
rect 10414 16496 10470 16532
rect 10046 11772 10048 11792
rect 10048 11772 10100 11792
rect 10100 11772 10102 11792
rect 10046 11736 10102 11772
rect 10138 11328 10194 11384
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11794 18536 11850 18592
rect 11794 18128 11850 18184
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 10874 15816 10930 15872
rect 10966 15000 11022 15056
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11978 17620 11980 17640
rect 11980 17620 12032 17640
rect 12032 17620 12034 17640
rect 11978 17584 12034 17620
rect 10966 11328 11022 11384
rect 10322 10104 10378 10160
rect 10230 9968 10286 10024
rect 10874 10124 10930 10160
rect 10874 10104 10876 10124
rect 10876 10104 10928 10124
rect 10928 10104 10930 10124
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 12346 16940 12348 16960
rect 12348 16940 12400 16960
rect 12400 16940 12402 16960
rect 12346 16904 12402 16940
rect 12254 15020 12310 15056
rect 12254 15000 12256 15020
rect 12256 15000 12308 15020
rect 12308 15000 12310 15020
rect 12346 13912 12402 13968
rect 12530 14320 12586 14376
rect 12990 17720 13046 17776
rect 12254 13776 12310 13832
rect 12438 13776 12494 13832
rect 12438 12280 12494 12336
rect 11518 11192 11574 11248
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11886 10648 11942 10704
rect 11058 9560 11114 9616
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 12254 9868 12256 9888
rect 12256 9868 12308 9888
rect 12308 9868 12310 9888
rect 12254 9832 12310 9868
rect 13542 19352 13598 19408
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14186 19080 14242 19136
rect 14094 15852 14096 15872
rect 14096 15852 14148 15872
rect 14148 15852 14150 15872
rect 14094 15816 14150 15852
rect 13266 12144 13322 12200
rect 12438 9968 12494 10024
rect 12438 9560 12494 9616
rect 15198 19352 15254 19408
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14646 18944 14702 19000
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 16118 18672 16174 18728
rect 16118 18264 16174 18320
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14462 11056 14518 11112
rect 14554 10512 14610 10568
rect 14094 9560 14150 9616
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 15658 12144 15714 12200
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 15750 10548 15752 10568
rect 15752 10548 15804 10568
rect 15804 10548 15806 10568
rect 15750 10512 15806 10548
rect 15750 9424 15806 9480
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 16670 11736 16726 11792
rect 17682 19216 17738 19272
rect 17682 18400 17738 18456
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18142 17720 18198 17776
rect 17130 16632 17186 16688
rect 17314 16496 17370 16552
rect 16854 11736 16910 11792
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 17406 12280 17462 12336
rect 16762 8900 16818 8936
rect 16762 8880 16764 8900
rect 16764 8880 16816 8900
rect 16816 8880 16818 8900
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18142 13796 18198 13832
rect 18142 13776 18144 13796
rect 18144 13776 18196 13796
rect 18196 13776 18198 13796
rect 18786 13504 18842 13560
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 17958 10648 18014 10704
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 20718 21664 20774 21720
rect 19246 18128 19302 18184
rect 20626 21256 20682 21312
rect 20534 20712 20590 20768
rect 21546 22616 21602 22672
rect 20074 18672 20130 18728
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18050 10376 18106 10432
rect 17958 9696 18014 9752
rect 17314 9424 17370 9480
rect 17682 9424 17738 9480
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 17130 2488 17186 2544
rect 17958 9016 18014 9072
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18786 10784 18842 10840
rect 19154 14320 19210 14376
rect 19614 13912 19670 13968
rect 19246 13368 19302 13424
rect 19062 11328 19118 11384
rect 19062 11228 19064 11248
rect 19064 11228 19116 11248
rect 19116 11228 19118 11248
rect 19062 11192 19118 11228
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 17958 7792 18014 7848
rect 18050 6160 18106 6216
rect 17958 5752 18014 5808
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18970 10648 19026 10704
rect 19338 11056 19394 11112
rect 19338 10784 19394 10840
rect 19338 10512 19394 10568
rect 18878 8880 18934 8936
rect 18786 8608 18842 8664
rect 18694 6704 18750 6760
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18142 5208 18198 5264
rect 17958 4800 18014 4856
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 19706 10784 19762 10840
rect 19154 9560 19210 9616
rect 19154 8472 19210 8528
rect 20626 17448 20682 17504
rect 20166 13232 20222 13288
rect 20442 13524 20498 13560
rect 20442 13504 20444 13524
rect 20444 13504 20496 13524
rect 20496 13504 20498 13524
rect 20534 13232 20590 13288
rect 20994 19760 21050 19816
rect 20902 19216 20958 19272
rect 21178 19352 21234 19408
rect 20994 18808 21050 18864
rect 21086 18400 21142 18456
rect 20994 17992 21050 18048
rect 21086 17040 21142 17096
rect 21086 15544 21142 15600
rect 21086 14592 21142 14648
rect 21362 20304 21418 20360
rect 21270 18264 21326 18320
rect 21270 16496 21326 16552
rect 22742 19080 22798 19136
rect 21914 18944 21970 19000
rect 21454 16088 21510 16144
rect 20350 12144 20406 12200
rect 19246 8064 19302 8120
rect 18970 7112 19026 7168
rect 18878 3440 18934 3496
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 17314 1536 17370 1592
rect 19062 992 19118 1048
rect 3422 584 3478 640
rect 20994 10104 21050 10160
rect 21362 15156 21418 15192
rect 21362 15136 21364 15156
rect 21364 15136 21416 15156
rect 21416 15136 21418 15156
rect 21362 14184 21418 14240
rect 21454 13776 21510 13832
rect 21730 10104 21786 10160
rect 20534 4392 20590 4448
rect 21546 3848 21602 3904
rect 20442 2896 20498 2952
rect 20350 1944 20406 2000
rect 19246 176 19302 232
<< metal3 >>
rect 0 22674 800 22704
rect 2773 22674 2839 22677
rect 0 22672 2839 22674
rect 0 22616 2778 22672
rect 2834 22616 2839 22672
rect 0 22614 2839 22616
rect 0 22584 800 22614
rect 2773 22611 2839 22614
rect 21541 22674 21607 22677
rect 22200 22674 23000 22704
rect 21541 22672 23000 22674
rect 21541 22616 21546 22672
rect 21602 22616 23000 22672
rect 21541 22614 23000 22616
rect 21541 22611 21607 22614
rect 22200 22584 23000 22614
rect 0 22266 800 22296
rect 2957 22266 3023 22269
rect 0 22264 3023 22266
rect 0 22208 2962 22264
rect 3018 22208 3023 22264
rect 0 22206 3023 22208
rect 0 22176 800 22206
rect 2957 22203 3023 22206
rect 21081 22266 21147 22269
rect 22200 22266 23000 22296
rect 21081 22264 23000 22266
rect 21081 22208 21086 22264
rect 21142 22208 23000 22264
rect 21081 22206 23000 22208
rect 21081 22203 21147 22206
rect 22200 22176 23000 22206
rect 0 21722 800 21752
rect 3141 21722 3207 21725
rect 0 21720 3207 21722
rect 0 21664 3146 21720
rect 3202 21664 3207 21720
rect 0 21662 3207 21664
rect 0 21632 800 21662
rect 3141 21659 3207 21662
rect 20713 21722 20779 21725
rect 22200 21722 23000 21752
rect 20713 21720 23000 21722
rect 20713 21664 20718 21720
rect 20774 21664 23000 21720
rect 20713 21662 23000 21664
rect 20713 21659 20779 21662
rect 22200 21632 23000 21662
rect 0 21314 800 21344
rect 4061 21314 4127 21317
rect 0 21312 4127 21314
rect 0 21256 4066 21312
rect 4122 21256 4127 21312
rect 0 21254 4127 21256
rect 0 21224 800 21254
rect 4061 21251 4127 21254
rect 20621 21314 20687 21317
rect 22200 21314 23000 21344
rect 20621 21312 23000 21314
rect 20621 21256 20626 21312
rect 20682 21256 23000 21312
rect 20621 21254 23000 21256
rect 20621 21251 20687 21254
rect 22200 21224 23000 21254
rect 0 20770 800 20800
rect 2865 20770 2931 20773
rect 0 20768 2931 20770
rect 0 20712 2870 20768
rect 2926 20712 2931 20768
rect 0 20710 2931 20712
rect 0 20680 800 20710
rect 2865 20707 2931 20710
rect 20529 20770 20595 20773
rect 22200 20770 23000 20800
rect 20529 20768 23000 20770
rect 20529 20712 20534 20768
rect 20590 20712 23000 20768
rect 20529 20710 23000 20712
rect 20529 20707 20595 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22200 20680 23000 20710
rect 18270 20639 18590 20640
rect 0 20362 800 20392
rect 3601 20362 3667 20365
rect 0 20360 3667 20362
rect 0 20304 3606 20360
rect 3662 20304 3667 20360
rect 0 20302 3667 20304
rect 0 20272 800 20302
rect 3601 20299 3667 20302
rect 21357 20362 21423 20365
rect 22200 20362 23000 20392
rect 21357 20360 23000 20362
rect 21357 20304 21362 20360
rect 21418 20304 23000 20360
rect 21357 20302 23000 20304
rect 21357 20299 21423 20302
rect 22200 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 2773 19818 2839 19821
rect 0 19816 2839 19818
rect 0 19760 2778 19816
rect 2834 19760 2839 19816
rect 0 19758 2839 19760
rect 0 19728 800 19758
rect 2773 19755 2839 19758
rect 20989 19818 21055 19821
rect 22200 19818 23000 19848
rect 20989 19816 23000 19818
rect 20989 19760 20994 19816
rect 21050 19760 23000 19816
rect 20989 19758 23000 19760
rect 20989 19755 21055 19758
rect 22200 19728 23000 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 1945 19410 2011 19413
rect 0 19408 2011 19410
rect 0 19352 1950 19408
rect 2006 19352 2011 19408
rect 0 19350 2011 19352
rect 0 19320 800 19350
rect 1945 19347 2011 19350
rect 2589 19410 2655 19413
rect 3417 19410 3483 19413
rect 2589 19408 3483 19410
rect 2589 19352 2594 19408
rect 2650 19352 3422 19408
rect 3478 19352 3483 19408
rect 2589 19350 3483 19352
rect 2589 19347 2655 19350
rect 3417 19347 3483 19350
rect 13537 19410 13603 19413
rect 15193 19410 15259 19413
rect 13537 19408 15259 19410
rect 13537 19352 13542 19408
rect 13598 19352 15198 19408
rect 15254 19352 15259 19408
rect 13537 19350 15259 19352
rect 13537 19347 13603 19350
rect 15193 19347 15259 19350
rect 21173 19410 21239 19413
rect 22200 19410 23000 19440
rect 21173 19408 23000 19410
rect 21173 19352 21178 19408
rect 21234 19352 23000 19408
rect 21173 19350 23000 19352
rect 21173 19347 21239 19350
rect 22200 19320 23000 19350
rect 2037 19274 2103 19277
rect 17677 19274 17743 19277
rect 20897 19274 20963 19277
rect 2037 19272 17602 19274
rect 2037 19216 2042 19272
rect 2098 19216 17602 19272
rect 2037 19214 17602 19216
rect 2037 19211 2103 19214
rect 1853 19138 1919 19141
rect 6637 19138 6703 19141
rect 1853 19136 6703 19138
rect 1853 19080 1858 19136
rect 1914 19080 6642 19136
rect 6698 19080 6703 19136
rect 1853 19078 6703 19080
rect 1853 19075 1919 19078
rect 6637 19075 6703 19078
rect 10133 19138 10199 19141
rect 14181 19138 14247 19141
rect 10133 19136 14247 19138
rect 10133 19080 10138 19136
rect 10194 19080 14186 19136
rect 14242 19080 14247 19136
rect 10133 19078 14247 19080
rect 17542 19138 17602 19214
rect 17677 19272 20963 19274
rect 17677 19216 17682 19272
rect 17738 19216 20902 19272
rect 20958 19216 20963 19272
rect 17677 19214 20963 19216
rect 17677 19211 17743 19214
rect 20897 19211 20963 19214
rect 22737 19138 22803 19141
rect 17542 19136 22803 19138
rect 17542 19080 22742 19136
rect 22798 19080 22803 19136
rect 17542 19078 22803 19080
rect 10133 19075 10199 19078
rect 14181 19075 14247 19078
rect 22737 19075 22803 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 1669 19002 1735 19005
rect 8293 19002 8359 19005
rect 14641 19002 14707 19005
rect 21909 19002 21975 19005
rect 1669 19000 2146 19002
rect 1669 18944 1674 19000
rect 1730 18944 2146 19000
rect 1669 18942 2146 18944
rect 1669 18939 1735 18942
rect 0 18866 800 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 2086 18866 2146 18942
rect 8293 19000 14707 19002
rect 8293 18944 8298 19000
rect 8354 18944 14646 19000
rect 14702 18944 14707 19000
rect 8293 18942 14707 18944
rect 8293 18939 8359 18942
rect 14641 18939 14707 18942
rect 17174 19000 21975 19002
rect 17174 18944 21914 19000
rect 21970 18944 21975 19000
rect 17174 18942 21975 18944
rect 17174 18866 17234 18942
rect 21909 18939 21975 18942
rect 2086 18806 17234 18866
rect 20989 18866 21055 18869
rect 22200 18866 23000 18896
rect 20989 18864 23000 18866
rect 20989 18808 20994 18864
rect 21050 18808 23000 18864
rect 20989 18806 23000 18808
rect 0 18776 800 18806
rect 1945 18803 2011 18806
rect 20989 18803 21055 18806
rect 22200 18776 23000 18806
rect 2681 18730 2747 18733
rect 16113 18730 16179 18733
rect 20069 18730 20135 18733
rect 2681 18728 16179 18730
rect 2681 18672 2686 18728
rect 2742 18672 16118 18728
rect 16174 18672 16179 18728
rect 2681 18670 16179 18672
rect 2681 18667 2747 18670
rect 16113 18667 16179 18670
rect 16254 18728 20135 18730
rect 16254 18672 20074 18728
rect 20130 18672 20135 18728
rect 16254 18670 20135 18672
rect 5993 18594 6059 18597
rect 9438 18594 9444 18596
rect 5993 18592 9444 18594
rect 5993 18536 5998 18592
rect 6054 18536 9444 18592
rect 5993 18534 9444 18536
rect 5993 18531 6059 18534
rect 9438 18532 9444 18534
rect 9508 18594 9514 18596
rect 9581 18594 9647 18597
rect 9508 18592 9647 18594
rect 9508 18536 9586 18592
rect 9642 18536 9647 18592
rect 9508 18534 9647 18536
rect 9508 18532 9514 18534
rect 9581 18531 9647 18534
rect 11789 18594 11855 18597
rect 16254 18594 16314 18670
rect 20069 18667 20135 18670
rect 11789 18592 16314 18594
rect 11789 18536 11794 18592
rect 11850 18536 16314 18592
rect 11789 18534 16314 18536
rect 11789 18531 11855 18534
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 2773 18458 2839 18461
rect 0 18456 2839 18458
rect 0 18400 2778 18456
rect 2834 18400 2839 18456
rect 0 18398 2839 18400
rect 0 18368 800 18398
rect 2773 18395 2839 18398
rect 7373 18458 7439 18461
rect 9029 18458 9095 18461
rect 17677 18458 17743 18461
rect 7373 18456 9095 18458
rect 7373 18400 7378 18456
rect 7434 18400 9034 18456
rect 9090 18400 9095 18456
rect 7373 18398 9095 18400
rect 7373 18395 7439 18398
rect 9029 18395 9095 18398
rect 11792 18456 17743 18458
rect 11792 18400 17682 18456
rect 17738 18400 17743 18456
rect 11792 18398 17743 18400
rect 6177 18322 6243 18325
rect 8477 18322 8543 18325
rect 6177 18320 8543 18322
rect 6177 18264 6182 18320
rect 6238 18264 8482 18320
rect 8538 18264 8543 18320
rect 6177 18262 8543 18264
rect 6177 18259 6243 18262
rect 8477 18259 8543 18262
rect 9673 18322 9739 18325
rect 11792 18322 11852 18398
rect 17677 18395 17743 18398
rect 21081 18458 21147 18461
rect 22200 18458 23000 18488
rect 21081 18456 23000 18458
rect 21081 18400 21086 18456
rect 21142 18400 23000 18456
rect 21081 18398 23000 18400
rect 21081 18395 21147 18398
rect 22200 18368 23000 18398
rect 9673 18320 11852 18322
rect 9673 18264 9678 18320
rect 9734 18264 11852 18320
rect 9673 18262 11852 18264
rect 16113 18322 16179 18325
rect 21265 18322 21331 18325
rect 16113 18320 21331 18322
rect 16113 18264 16118 18320
rect 16174 18264 21270 18320
rect 21326 18264 21331 18320
rect 16113 18262 21331 18264
rect 9673 18259 9739 18262
rect 16113 18259 16179 18262
rect 21265 18259 21331 18262
rect 2405 18186 2471 18189
rect 9078 18186 9506 18220
rect 11789 18186 11855 18189
rect 19241 18186 19307 18189
rect 2405 18184 11855 18186
rect 2405 18128 2410 18184
rect 2466 18160 11794 18184
rect 2466 18128 9138 18160
rect 2405 18126 9138 18128
rect 9446 18128 11794 18160
rect 11850 18128 11855 18184
rect 9446 18126 11855 18128
rect 2405 18123 2471 18126
rect 11789 18123 11855 18126
rect 14414 18184 19307 18186
rect 14414 18128 19246 18184
rect 19302 18128 19307 18184
rect 14414 18126 19307 18128
rect 0 18050 800 18080
rect 1945 18050 2011 18053
rect 0 18048 2011 18050
rect 0 17992 1950 18048
rect 2006 17992 2011 18048
rect 0 17990 2011 17992
rect 0 17960 800 17990
rect 1945 17987 2011 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14414 17914 14474 18126
rect 19241 18123 19307 18126
rect 20989 18050 21055 18053
rect 22200 18050 23000 18080
rect 20989 18048 23000 18050
rect 20989 17992 20994 18048
rect 21050 17992 23000 18048
rect 20989 17990 23000 17992
rect 20989 17987 21055 17990
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 8296 17854 14474 17914
rect 4061 17778 4127 17781
rect 8296 17778 8356 17854
rect 4061 17776 8356 17778
rect 4061 17720 4066 17776
rect 4122 17720 8356 17776
rect 4061 17718 8356 17720
rect 12985 17778 13051 17781
rect 18137 17778 18203 17781
rect 12985 17776 18203 17778
rect 12985 17720 12990 17776
rect 13046 17720 18142 17776
rect 18198 17720 18203 17776
rect 12985 17718 18203 17720
rect 4061 17715 4127 17718
rect 12985 17715 13051 17718
rect 18137 17715 18203 17718
rect 9673 17642 9739 17645
rect 11973 17642 12039 17645
rect 9673 17640 12039 17642
rect 9673 17584 9678 17640
rect 9734 17584 11978 17640
rect 12034 17584 12039 17640
rect 9673 17582 12039 17584
rect 9673 17579 9739 17582
rect 11973 17579 12039 17582
rect 0 17506 800 17536
rect 2865 17506 2931 17509
rect 0 17504 2931 17506
rect 0 17448 2870 17504
rect 2926 17448 2931 17504
rect 0 17446 2931 17448
rect 0 17416 800 17446
rect 2865 17443 2931 17446
rect 4797 17506 4863 17509
rect 10317 17506 10383 17509
rect 4797 17504 10383 17506
rect 4797 17448 4802 17504
rect 4858 17448 10322 17504
rect 10378 17448 10383 17504
rect 4797 17446 10383 17448
rect 4797 17443 4863 17446
rect 10317 17443 10383 17446
rect 20621 17506 20687 17509
rect 22200 17506 23000 17536
rect 20621 17504 23000 17506
rect 20621 17448 20626 17504
rect 20682 17448 23000 17504
rect 20621 17446 23000 17448
rect 20621 17443 20687 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22200 17416 23000 17446
rect 18270 17375 18590 17376
rect 0 17098 800 17128
rect 1945 17098 2011 17101
rect 0 17096 2011 17098
rect 0 17040 1950 17096
rect 2006 17040 2011 17096
rect 0 17038 2011 17040
rect 0 17008 800 17038
rect 1945 17035 2011 17038
rect 21081 17098 21147 17101
rect 22200 17098 23000 17128
rect 21081 17096 23000 17098
rect 21081 17040 21086 17096
rect 21142 17040 23000 17096
rect 21081 17038 23000 17040
rect 21081 17035 21147 17038
rect 22200 17008 23000 17038
rect 10317 16962 10383 16965
rect 12341 16962 12407 16965
rect 10317 16960 12407 16962
rect 10317 16904 10322 16960
rect 10378 16904 12346 16960
rect 12402 16904 12407 16960
rect 10317 16902 12407 16904
rect 10317 16899 10383 16902
rect 12341 16899 12407 16902
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 8661 16690 8727 16693
rect 17125 16690 17191 16693
rect 8661 16688 17191 16690
rect 8661 16632 8666 16688
rect 8722 16632 17130 16688
rect 17186 16632 17191 16688
rect 8661 16630 17191 16632
rect 8661 16627 8727 16630
rect 17125 16627 17191 16630
rect 0 16554 800 16584
rect 2773 16554 2839 16557
rect 0 16552 2839 16554
rect 0 16496 2778 16552
rect 2834 16496 2839 16552
rect 0 16494 2839 16496
rect 0 16464 800 16494
rect 2773 16491 2839 16494
rect 10409 16554 10475 16557
rect 17309 16554 17375 16557
rect 10409 16552 17375 16554
rect 10409 16496 10414 16552
rect 10470 16496 17314 16552
rect 17370 16496 17375 16552
rect 10409 16494 17375 16496
rect 10409 16491 10475 16494
rect 17309 16491 17375 16494
rect 21265 16554 21331 16557
rect 22200 16554 23000 16584
rect 21265 16552 23000 16554
rect 21265 16496 21270 16552
rect 21326 16496 23000 16552
rect 21265 16494 23000 16496
rect 21265 16491 21331 16494
rect 22200 16464 23000 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1945 16146 2011 16149
rect 0 16144 2011 16146
rect 0 16088 1950 16144
rect 2006 16088 2011 16144
rect 0 16086 2011 16088
rect 0 16056 800 16086
rect 1945 16083 2011 16086
rect 21449 16146 21515 16149
rect 22200 16146 23000 16176
rect 21449 16144 23000 16146
rect 21449 16088 21454 16144
rect 21510 16088 23000 16144
rect 21449 16086 23000 16088
rect 21449 16083 21515 16086
rect 22200 16056 23000 16086
rect 10869 15874 10935 15877
rect 14089 15874 14155 15877
rect 10869 15872 14155 15874
rect 10869 15816 10874 15872
rect 10930 15816 14094 15872
rect 14150 15816 14155 15872
rect 10869 15814 14155 15816
rect 10869 15811 10935 15814
rect 14089 15811 14155 15814
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 2773 15602 2839 15605
rect 0 15600 2839 15602
rect 0 15544 2778 15600
rect 2834 15544 2839 15600
rect 0 15542 2839 15544
rect 0 15512 800 15542
rect 2773 15539 2839 15542
rect 21081 15602 21147 15605
rect 22200 15602 23000 15632
rect 21081 15600 23000 15602
rect 21081 15544 21086 15600
rect 21142 15544 23000 15600
rect 21081 15542 23000 15544
rect 21081 15539 21147 15542
rect 22200 15512 23000 15542
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 1945 15194 2011 15197
rect 0 15192 2011 15194
rect 0 15136 1950 15192
rect 2006 15136 2011 15192
rect 0 15134 2011 15136
rect 0 15104 800 15134
rect 1945 15131 2011 15134
rect 21357 15194 21423 15197
rect 22200 15194 23000 15224
rect 21357 15192 23000 15194
rect 21357 15136 21362 15192
rect 21418 15136 23000 15192
rect 21357 15134 23000 15136
rect 21357 15131 21423 15134
rect 22200 15104 23000 15134
rect 10961 15058 11027 15061
rect 12249 15058 12315 15061
rect 10961 15056 12315 15058
rect 10961 15000 10966 15056
rect 11022 15000 12254 15056
rect 12310 15000 12315 15056
rect 10961 14998 12315 15000
rect 10961 14995 11027 14998
rect 12249 14995 12315 14998
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1945 14650 2011 14653
rect 0 14648 2011 14650
rect 0 14592 1950 14648
rect 2006 14592 2011 14648
rect 0 14590 2011 14592
rect 0 14560 800 14590
rect 1945 14587 2011 14590
rect 21081 14650 21147 14653
rect 22200 14650 23000 14680
rect 21081 14648 23000 14650
rect 21081 14592 21086 14648
rect 21142 14592 23000 14648
rect 21081 14590 23000 14592
rect 21081 14587 21147 14590
rect 22200 14560 23000 14590
rect 12525 14378 12591 14381
rect 19149 14378 19215 14381
rect 12525 14376 19215 14378
rect 12525 14320 12530 14376
rect 12586 14320 19154 14376
rect 19210 14320 19215 14376
rect 12525 14318 19215 14320
rect 12525 14315 12591 14318
rect 19149 14315 19215 14318
rect 0 14242 800 14272
rect 2865 14242 2931 14245
rect 0 14240 2931 14242
rect 0 14184 2870 14240
rect 2926 14184 2931 14240
rect 0 14182 2931 14184
rect 0 14152 800 14182
rect 2865 14179 2931 14182
rect 21357 14242 21423 14245
rect 22200 14242 23000 14272
rect 21357 14240 23000 14242
rect 21357 14184 21362 14240
rect 21418 14184 23000 14240
rect 21357 14182 23000 14184
rect 21357 14179 21423 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 12341 13970 12407 13973
rect 19609 13970 19675 13973
rect 12341 13968 19675 13970
rect 12341 13912 12346 13968
rect 12402 13912 19614 13968
rect 19670 13912 19675 13968
rect 12341 13910 19675 13912
rect 12341 13907 12407 13910
rect 19609 13907 19675 13910
rect 0 13834 800 13864
rect 2773 13834 2839 13837
rect 0 13832 2839 13834
rect 0 13776 2778 13832
rect 2834 13776 2839 13832
rect 0 13774 2839 13776
rect 0 13744 800 13774
rect 2773 13771 2839 13774
rect 12249 13834 12315 13837
rect 12433 13834 12499 13837
rect 18137 13834 18203 13837
rect 12249 13832 18203 13834
rect 12249 13776 12254 13832
rect 12310 13776 12438 13832
rect 12494 13776 18142 13832
rect 18198 13776 18203 13832
rect 12249 13774 18203 13776
rect 12249 13771 12315 13774
rect 12433 13771 12499 13774
rect 18137 13771 18203 13774
rect 21449 13834 21515 13837
rect 22200 13834 23000 13864
rect 21449 13832 23000 13834
rect 21449 13776 21454 13832
rect 21510 13776 23000 13832
rect 21449 13774 23000 13776
rect 21449 13771 21515 13774
rect 22200 13744 23000 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 18781 13562 18847 13565
rect 20437 13562 20503 13565
rect 18781 13560 20503 13562
rect 18781 13504 18786 13560
rect 18842 13504 20442 13560
rect 20498 13504 20503 13560
rect 18781 13502 20503 13504
rect 18781 13499 18847 13502
rect 20437 13499 20503 13502
rect 10041 13426 10107 13429
rect 19006 13426 19012 13428
rect 10041 13424 19012 13426
rect 10041 13368 10046 13424
rect 10102 13368 19012 13424
rect 10041 13366 19012 13368
rect 10041 13363 10107 13366
rect 19006 13364 19012 13366
rect 19076 13426 19082 13428
rect 19241 13426 19307 13429
rect 19076 13424 19307 13426
rect 19076 13368 19246 13424
rect 19302 13368 19307 13424
rect 19076 13366 19307 13368
rect 19076 13364 19082 13366
rect 19241 13363 19307 13366
rect 0 13290 800 13320
rect 2221 13290 2287 13293
rect 0 13288 2287 13290
rect 0 13232 2226 13288
rect 2282 13232 2287 13288
rect 0 13230 2287 13232
rect 0 13200 800 13230
rect 2221 13227 2287 13230
rect 8753 13290 8819 13293
rect 20161 13290 20227 13293
rect 20529 13290 20595 13293
rect 22200 13290 23000 13320
rect 8753 13288 20408 13290
rect 8753 13232 8758 13288
rect 8814 13232 20166 13288
rect 20222 13232 20408 13288
rect 8753 13230 20408 13232
rect 8753 13227 8819 13230
rect 20161 13227 20227 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 4061 12882 4127 12885
rect 0 12880 4127 12882
rect 0 12824 4066 12880
rect 4122 12824 4127 12880
rect 0 12822 4127 12824
rect 20348 12882 20408 13230
rect 20529 13288 23000 13290
rect 20529 13232 20534 13288
rect 20590 13232 23000 13288
rect 20529 13230 23000 13232
rect 20529 13227 20595 13230
rect 22200 13200 23000 13230
rect 22200 12882 23000 12912
rect 20348 12822 23000 12882
rect 0 12792 800 12822
rect 4061 12819 4127 12822
rect 22200 12792 23000 12822
rect 2681 12746 2747 12749
rect 9121 12746 9187 12749
rect 2681 12744 9187 12746
rect 2681 12688 2686 12744
rect 2742 12688 9126 12744
rect 9182 12688 9187 12744
rect 2681 12686 9187 12688
rect 2681 12683 2747 12686
rect 9121 12683 9187 12686
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 3509 12474 3575 12477
rect 5533 12474 5599 12477
rect 3509 12472 5599 12474
rect 3509 12416 3514 12472
rect 3570 12416 5538 12472
rect 5594 12416 5599 12472
rect 3509 12414 5599 12416
rect 3509 12411 3575 12414
rect 5533 12411 5599 12414
rect 0 12338 800 12368
rect 4521 12338 4587 12341
rect 9949 12338 10015 12341
rect 0 12278 4354 12338
rect 0 12248 800 12278
rect 4294 12202 4354 12278
rect 4521 12336 10015 12338
rect 4521 12280 4526 12336
rect 4582 12280 9954 12336
rect 10010 12280 10015 12336
rect 4521 12278 10015 12280
rect 4521 12275 4587 12278
rect 9949 12275 10015 12278
rect 12433 12338 12499 12341
rect 17401 12338 17467 12341
rect 22200 12338 23000 12368
rect 12433 12336 23000 12338
rect 12433 12280 12438 12336
rect 12494 12280 17406 12336
rect 17462 12280 23000 12336
rect 12433 12278 23000 12280
rect 12433 12275 12499 12278
rect 17401 12275 17467 12278
rect 22200 12248 23000 12278
rect 9489 12202 9555 12205
rect 4294 12200 9555 12202
rect 4294 12144 9494 12200
rect 9550 12144 9555 12200
rect 4294 12142 9555 12144
rect 9489 12139 9555 12142
rect 9765 12202 9831 12205
rect 13261 12202 13327 12205
rect 9765 12200 13327 12202
rect 9765 12144 9770 12200
rect 9826 12144 13266 12200
rect 13322 12144 13327 12200
rect 9765 12142 13327 12144
rect 9765 12139 9831 12142
rect 13261 12139 13327 12142
rect 15653 12202 15719 12205
rect 20345 12202 20411 12205
rect 15653 12200 20411 12202
rect 15653 12144 15658 12200
rect 15714 12144 20350 12200
rect 20406 12144 20411 12200
rect 15653 12142 20411 12144
rect 15653 12139 15719 12142
rect 20345 12139 20411 12142
rect 4409 12000 4729 12001
rect 0 11930 800 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 4061 11930 4127 11933
rect 22200 11930 23000 11960
rect 0 11928 4127 11930
rect 0 11872 4066 11928
rect 4122 11872 4127 11928
rect 0 11870 4127 11872
rect 0 11840 800 11870
rect 4061 11867 4127 11870
rect 18692 11870 23000 11930
rect 3969 11794 4035 11797
rect 9581 11794 9647 11797
rect 3969 11792 9647 11794
rect 3969 11736 3974 11792
rect 4030 11736 9586 11792
rect 9642 11736 9647 11792
rect 3969 11734 9647 11736
rect 3969 11731 4035 11734
rect 9581 11731 9647 11734
rect 10041 11794 10107 11797
rect 16665 11794 16731 11797
rect 10041 11792 16731 11794
rect 10041 11736 10046 11792
rect 10102 11736 16670 11792
rect 16726 11736 16731 11792
rect 10041 11734 16731 11736
rect 10041 11731 10107 11734
rect 16665 11731 16731 11734
rect 16849 11794 16915 11797
rect 18692 11794 18752 11870
rect 22200 11840 23000 11870
rect 16849 11792 18752 11794
rect 16849 11736 16854 11792
rect 16910 11736 18752 11792
rect 16849 11734 18752 11736
rect 16849 11731 16915 11734
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 3233 11386 3299 11389
rect 0 11384 3299 11386
rect 0 11328 3238 11384
rect 3294 11328 3299 11384
rect 0 11326 3299 11328
rect 0 11296 800 11326
rect 3233 11323 3299 11326
rect 10133 11386 10199 11389
rect 10961 11386 11027 11389
rect 10133 11384 11027 11386
rect 10133 11328 10138 11384
rect 10194 11328 10966 11384
rect 11022 11328 11027 11384
rect 10133 11326 11027 11328
rect 10133 11323 10199 11326
rect 10961 11323 11027 11326
rect 19057 11386 19123 11389
rect 22200 11386 23000 11416
rect 19057 11384 23000 11386
rect 19057 11328 19062 11384
rect 19118 11328 23000 11384
rect 19057 11326 23000 11328
rect 19057 11323 19123 11326
rect 22200 11296 23000 11326
rect 11513 11250 11579 11253
rect 19057 11250 19123 11253
rect 11513 11248 19123 11250
rect 11513 11192 11518 11248
rect 11574 11192 19062 11248
rect 19118 11192 19123 11248
rect 11513 11190 19123 11192
rect 11513 11187 11579 11190
rect 19057 11187 19123 11190
rect 9121 11114 9187 11117
rect 4110 11112 9187 11114
rect 4110 11056 9126 11112
rect 9182 11056 9187 11112
rect 4110 11054 9187 11056
rect 0 10978 800 11008
rect 4110 10978 4170 11054
rect 9121 11051 9187 11054
rect 14457 11114 14523 11117
rect 19333 11116 19399 11117
rect 14457 11112 18752 11114
rect 14457 11056 14462 11112
rect 14518 11056 18752 11112
rect 14457 11054 18752 11056
rect 14457 11051 14523 11054
rect 0 10918 4170 10978
rect 18692 10978 18752 11054
rect 19333 11112 19380 11116
rect 19444 11114 19450 11116
rect 19333 11056 19338 11112
rect 19333 11052 19380 11056
rect 19444 11054 19490 11114
rect 19444 11052 19450 11054
rect 19333 11051 19399 11052
rect 22200 10978 23000 11008
rect 18692 10918 23000 10978
rect 0 10888 800 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 22200 10888 23000 10918
rect 18270 10847 18590 10848
rect 18781 10842 18847 10845
rect 19006 10842 19012 10844
rect 18781 10840 19012 10842
rect 18781 10784 18786 10840
rect 18842 10784 19012 10840
rect 18781 10782 19012 10784
rect 18781 10779 18847 10782
rect 19006 10780 19012 10782
rect 19076 10780 19082 10844
rect 19333 10842 19399 10845
rect 19701 10842 19767 10845
rect 19333 10840 19767 10842
rect 19333 10784 19338 10840
rect 19394 10784 19706 10840
rect 19762 10784 19767 10840
rect 19333 10782 19767 10784
rect 19333 10779 19399 10782
rect 19701 10779 19767 10782
rect 11881 10706 11947 10709
rect 17953 10706 18019 10709
rect 18965 10706 19031 10709
rect 11881 10704 19031 10706
rect 11881 10648 11886 10704
rect 11942 10648 17958 10704
rect 18014 10648 18970 10704
rect 19026 10648 19031 10704
rect 11881 10646 19031 10648
rect 11881 10643 11947 10646
rect 17953 10643 18019 10646
rect 18965 10643 19031 10646
rect 14549 10570 14615 10573
rect 15745 10570 15811 10573
rect 14549 10568 15811 10570
rect 14549 10512 14554 10568
rect 14610 10512 15750 10568
rect 15806 10512 15811 10568
rect 14549 10510 15811 10512
rect 14549 10507 14615 10510
rect 15745 10507 15811 10510
rect 19333 10572 19399 10573
rect 19333 10568 19380 10572
rect 19444 10570 19450 10572
rect 19333 10512 19338 10568
rect 19333 10508 19380 10512
rect 19444 10510 19490 10570
rect 19444 10508 19450 10510
rect 19333 10507 19399 10508
rect 0 10434 800 10464
rect 3785 10434 3851 10437
rect 0 10432 3851 10434
rect 0 10376 3790 10432
rect 3846 10376 3851 10432
rect 0 10374 3851 10376
rect 0 10344 800 10374
rect 3785 10371 3851 10374
rect 18045 10434 18111 10437
rect 22200 10434 23000 10464
rect 18045 10432 23000 10434
rect 18045 10376 18050 10432
rect 18106 10376 23000 10432
rect 18045 10374 23000 10376
rect 18045 10371 18111 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 4153 10162 4219 10165
rect 5165 10162 5231 10165
rect 4153 10160 5231 10162
rect 4153 10104 4158 10160
rect 4214 10104 5170 10160
rect 5226 10104 5231 10160
rect 4153 10102 5231 10104
rect 4153 10099 4219 10102
rect 5165 10099 5231 10102
rect 10317 10162 10383 10165
rect 10869 10162 10935 10165
rect 20989 10162 21055 10165
rect 21725 10162 21791 10165
rect 10317 10160 10935 10162
rect 10317 10104 10322 10160
rect 10378 10104 10874 10160
rect 10930 10104 10935 10160
rect 10317 10102 10935 10104
rect 10317 10099 10383 10102
rect 10869 10099 10935 10102
rect 16622 10160 21791 10162
rect 16622 10104 20994 10160
rect 21050 10104 21730 10160
rect 21786 10104 21791 10160
rect 16622 10102 21791 10104
rect 0 10026 800 10056
rect 3969 10026 4035 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 800 9966
rect 3969 9963 4035 9966
rect 8385 10026 8451 10029
rect 9489 10028 9555 10029
rect 9438 10026 9444 10028
rect 8385 10024 9444 10026
rect 9508 10026 9555 10028
rect 10225 10026 10291 10029
rect 12433 10026 12499 10029
rect 16622 10026 16682 10102
rect 20989 10099 21055 10102
rect 21725 10099 21791 10102
rect 22200 10026 23000 10056
rect 9508 10024 9600 10026
rect 8385 9968 8390 10024
rect 8446 9968 9444 10024
rect 9550 9968 9600 10024
rect 8385 9966 9444 9968
rect 8385 9963 8451 9966
rect 9438 9964 9444 9966
rect 9508 9966 9600 9968
rect 10225 10024 11852 10026
rect 10225 9968 10230 10024
rect 10286 9968 11852 10024
rect 10225 9966 11852 9968
rect 9508 9964 9555 9966
rect 9489 9963 9555 9964
rect 10225 9963 10291 9966
rect 1669 9890 1735 9893
rect 3509 9890 3575 9893
rect 1669 9888 3575 9890
rect 1669 9832 1674 9888
rect 1730 9832 3514 9888
rect 3570 9832 3575 9888
rect 1669 9830 3575 9832
rect 1669 9827 1735 9830
rect 3509 9827 3575 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 11792 9754 11852 9966
rect 12433 10024 16682 10026
rect 12433 9968 12438 10024
rect 12494 9968 16682 10024
rect 12433 9966 16682 9968
rect 16806 9966 23000 10026
rect 12433 9963 12499 9966
rect 12249 9890 12315 9893
rect 16806 9890 16866 9966
rect 22200 9936 23000 9966
rect 12249 9888 16866 9890
rect 12249 9832 12254 9888
rect 12310 9832 16866 9888
rect 12249 9830 16866 9832
rect 12249 9827 12315 9830
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 17953 9754 18019 9757
rect 11792 9752 18019 9754
rect 11792 9696 17958 9752
rect 18014 9696 18019 9752
rect 11792 9694 18019 9696
rect 17953 9691 18019 9694
rect 11053 9618 11119 9621
rect 12433 9618 12499 9621
rect 11053 9616 12499 9618
rect 11053 9560 11058 9616
rect 11114 9560 12438 9616
rect 12494 9560 12499 9616
rect 11053 9558 12499 9560
rect 11053 9555 11119 9558
rect 12433 9555 12499 9558
rect 14089 9618 14155 9621
rect 19149 9618 19215 9621
rect 14089 9616 19215 9618
rect 14089 9560 14094 9616
rect 14150 9560 19154 9616
rect 19210 9560 19215 9616
rect 14089 9558 19215 9560
rect 14089 9555 14155 9558
rect 19149 9555 19215 9558
rect 0 9482 800 9512
rect 3417 9482 3483 9485
rect 0 9480 3483 9482
rect 0 9424 3422 9480
rect 3478 9424 3483 9480
rect 0 9422 3483 9424
rect 0 9392 800 9422
rect 3417 9419 3483 9422
rect 15745 9482 15811 9485
rect 17309 9482 17375 9485
rect 15745 9480 17375 9482
rect 15745 9424 15750 9480
rect 15806 9424 17314 9480
rect 17370 9424 17375 9480
rect 15745 9422 17375 9424
rect 15745 9419 15811 9422
rect 17309 9419 17375 9422
rect 17677 9482 17743 9485
rect 22200 9482 23000 9512
rect 17677 9480 23000 9482
rect 17677 9424 17682 9480
rect 17738 9424 23000 9480
rect 17677 9422 23000 9424
rect 17677 9419 17743 9422
rect 22200 9392 23000 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 17953 9074 18019 9077
rect 22200 9074 23000 9104
rect 17953 9072 23000 9074
rect 17953 9016 17958 9072
rect 18014 9016 23000 9072
rect 17953 9014 23000 9016
rect 17953 9011 18019 9014
rect 22200 8984 23000 9014
rect 16757 8938 16823 8941
rect 18873 8938 18939 8941
rect 16757 8936 18939 8938
rect 16757 8880 16762 8936
rect 16818 8880 18878 8936
rect 18934 8880 18939 8936
rect 16757 8878 18939 8880
rect 16757 8875 16823 8878
rect 18873 8875 18939 8878
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 4061 8666 4127 8669
rect 0 8664 4127 8666
rect 0 8608 4066 8664
rect 4122 8608 4127 8664
rect 0 8606 4127 8608
rect 0 8576 800 8606
rect 4061 8603 4127 8606
rect 18781 8666 18847 8669
rect 22200 8666 23000 8696
rect 18781 8664 23000 8666
rect 18781 8608 18786 8664
rect 18842 8608 23000 8664
rect 18781 8606 23000 8608
rect 18781 8603 18847 8606
rect 22200 8576 23000 8606
rect 19149 8532 19215 8533
rect 19149 8530 19196 8532
rect 19104 8528 19196 8530
rect 19104 8472 19154 8528
rect 19104 8470 19196 8472
rect 19149 8468 19196 8470
rect 19260 8468 19266 8532
rect 19149 8467 19215 8468
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 6913 8122 6979 8125
rect 0 8120 6979 8122
rect 0 8064 6918 8120
rect 6974 8064 6979 8120
rect 0 8062 6979 8064
rect 0 8032 800 8062
rect 6913 8059 6979 8062
rect 19241 8122 19307 8125
rect 22200 8122 23000 8152
rect 19241 8120 23000 8122
rect 19241 8064 19246 8120
rect 19302 8064 23000 8120
rect 19241 8062 23000 8064
rect 19241 8059 19307 8062
rect 22200 8032 23000 8062
rect 6545 7850 6611 7853
rect 8017 7850 8083 7853
rect 6545 7848 8083 7850
rect 6545 7792 6550 7848
rect 6606 7792 8022 7848
rect 8078 7792 8083 7848
rect 6545 7790 8083 7792
rect 6545 7787 6611 7790
rect 8017 7787 8083 7790
rect 17953 7850 18019 7853
rect 17953 7848 18890 7850
rect 17953 7792 17958 7848
rect 18014 7792 18890 7848
rect 17953 7790 18890 7792
rect 17953 7787 18019 7790
rect 0 7714 800 7744
rect 3601 7714 3667 7717
rect 0 7712 3667 7714
rect 0 7656 3606 7712
rect 3662 7656 3667 7712
rect 0 7654 3667 7656
rect 18830 7714 18890 7790
rect 22200 7714 23000 7744
rect 18830 7654 23000 7714
rect 0 7624 800 7654
rect 3601 7651 3667 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22200 7624 23000 7654
rect 18270 7583 18590 7584
rect 0 7170 800 7200
rect 3969 7170 4035 7173
rect 0 7168 4035 7170
rect 0 7112 3974 7168
rect 4030 7112 4035 7168
rect 0 7110 4035 7112
rect 0 7080 800 7110
rect 3969 7107 4035 7110
rect 18965 7170 19031 7173
rect 22200 7170 23000 7200
rect 18965 7168 23000 7170
rect 18965 7112 18970 7168
rect 19026 7112 23000 7168
rect 18965 7110 23000 7112
rect 18965 7107 19031 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22200 7080 23000 7110
rect 14805 7039 15125 7040
rect 0 6762 800 6792
rect 3969 6762 4035 6765
rect 0 6760 4035 6762
rect 0 6704 3974 6760
rect 4030 6704 4035 6760
rect 0 6702 4035 6704
rect 0 6672 800 6702
rect 3969 6699 4035 6702
rect 18689 6762 18755 6765
rect 22200 6762 23000 6792
rect 18689 6760 23000 6762
rect 18689 6704 18694 6760
rect 18750 6704 23000 6760
rect 18689 6702 23000 6704
rect 18689 6699 18755 6702
rect 22200 6672 23000 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 18045 6218 18111 6221
rect 22200 6218 23000 6248
rect 18045 6216 23000 6218
rect 18045 6160 18050 6216
rect 18106 6160 23000 6216
rect 18045 6158 23000 6160
rect 18045 6155 18111 6158
rect 22200 6128 23000 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 1485 5810 1551 5813
rect 0 5808 1551 5810
rect 0 5752 1490 5808
rect 1546 5752 1551 5808
rect 0 5750 1551 5752
rect 0 5720 800 5750
rect 1485 5747 1551 5750
rect 17953 5810 18019 5813
rect 22200 5810 23000 5840
rect 17953 5808 23000 5810
rect 17953 5752 17958 5808
rect 18014 5752 23000 5808
rect 17953 5750 23000 5752
rect 17953 5747 18019 5750
rect 22200 5720 23000 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5266 800 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 800 5206
rect 4061 5203 4127 5206
rect 18137 5266 18203 5269
rect 22200 5266 23000 5296
rect 18137 5264 23000 5266
rect 18137 5208 18142 5264
rect 18198 5208 23000 5264
rect 18137 5206 23000 5208
rect 18137 5203 18203 5206
rect 22200 5176 23000 5206
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 3325 4858 3391 4861
rect 0 4856 3391 4858
rect 0 4800 3330 4856
rect 3386 4800 3391 4856
rect 0 4798 3391 4800
rect 0 4768 800 4798
rect 3325 4795 3391 4798
rect 17953 4858 18019 4861
rect 22200 4858 23000 4888
rect 17953 4856 23000 4858
rect 17953 4800 17958 4856
rect 18014 4800 23000 4856
rect 17953 4798 23000 4800
rect 17953 4795 18019 4798
rect 22200 4768 23000 4798
rect 0 4450 800 4480
rect 3049 4450 3115 4453
rect 0 4448 3115 4450
rect 0 4392 3054 4448
rect 3110 4392 3115 4448
rect 0 4390 3115 4392
rect 0 4360 800 4390
rect 3049 4387 3115 4390
rect 20529 4450 20595 4453
rect 22200 4450 23000 4480
rect 20529 4448 23000 4450
rect 20529 4392 20534 4448
rect 20590 4392 23000 4448
rect 20529 4390 23000 4392
rect 20529 4387 20595 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22200 4360 23000 4390
rect 18270 4319 18590 4320
rect 0 3906 800 3936
rect 4153 3906 4219 3909
rect 0 3904 4219 3906
rect 0 3848 4158 3904
rect 4214 3848 4219 3904
rect 0 3846 4219 3848
rect 0 3816 800 3846
rect 4153 3843 4219 3846
rect 21541 3906 21607 3909
rect 22200 3906 23000 3936
rect 21541 3904 23000 3906
rect 21541 3848 21546 3904
rect 21602 3848 23000 3904
rect 21541 3846 23000 3848
rect 21541 3843 21607 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 0 3498 800 3528
rect 3601 3498 3667 3501
rect 0 3496 3667 3498
rect 0 3440 3606 3496
rect 3662 3440 3667 3496
rect 0 3438 3667 3440
rect 0 3408 800 3438
rect 3601 3435 3667 3438
rect 18873 3498 18939 3501
rect 22200 3498 23000 3528
rect 18873 3496 23000 3498
rect 18873 3440 18878 3496
rect 18934 3440 23000 3496
rect 18873 3438 23000 3440
rect 18873 3435 18939 3438
rect 22200 3408 23000 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 0 2954 800 2984
rect 4337 2954 4403 2957
rect 0 2952 4403 2954
rect 0 2896 4342 2952
rect 4398 2896 4403 2952
rect 0 2894 4403 2896
rect 0 2864 800 2894
rect 4337 2891 4403 2894
rect 20437 2954 20503 2957
rect 22200 2954 23000 2984
rect 20437 2952 23000 2954
rect 20437 2896 20442 2952
rect 20498 2896 23000 2952
rect 20437 2894 23000 2896
rect 20437 2891 20503 2894
rect 22200 2864 23000 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 2681 2546 2747 2549
rect 0 2544 2747 2546
rect 0 2488 2686 2544
rect 2742 2488 2747 2544
rect 0 2486 2747 2488
rect 0 2456 800 2486
rect 2681 2483 2747 2486
rect 17125 2546 17191 2549
rect 22200 2546 23000 2576
rect 17125 2544 23000 2546
rect 17125 2488 17130 2544
rect 17186 2488 23000 2544
rect 17125 2486 23000 2488
rect 17125 2483 17191 2486
rect 22200 2456 23000 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 3325 2002 3391 2005
rect 0 2000 3391 2002
rect 0 1944 3330 2000
rect 3386 1944 3391 2000
rect 0 1942 3391 1944
rect 0 1912 800 1942
rect 3325 1939 3391 1942
rect 20345 2002 20411 2005
rect 22200 2002 23000 2032
rect 20345 2000 23000 2002
rect 20345 1944 20350 2000
rect 20406 1944 23000 2000
rect 20345 1942 23000 1944
rect 20345 1939 20411 1942
rect 22200 1912 23000 1942
rect 0 1594 800 1624
rect 2773 1594 2839 1597
rect 0 1592 2839 1594
rect 0 1536 2778 1592
rect 2834 1536 2839 1592
rect 0 1534 2839 1536
rect 0 1504 800 1534
rect 2773 1531 2839 1534
rect 17309 1594 17375 1597
rect 22200 1594 23000 1624
rect 17309 1592 23000 1594
rect 17309 1536 17314 1592
rect 17370 1536 23000 1592
rect 17309 1534 23000 1536
rect 17309 1531 17375 1534
rect 22200 1504 23000 1534
rect 0 1050 800 1080
rect 4061 1050 4127 1053
rect 0 1048 4127 1050
rect 0 992 4066 1048
rect 4122 992 4127 1048
rect 0 990 4127 992
rect 0 960 800 990
rect 4061 987 4127 990
rect 19057 1050 19123 1053
rect 22200 1050 23000 1080
rect 19057 1048 23000 1050
rect 19057 992 19062 1048
rect 19118 992 23000 1048
rect 19057 990 23000 992
rect 19057 987 19123 990
rect 22200 960 23000 990
rect 0 642 800 672
rect 3417 642 3483 645
rect 0 640 3483 642
rect 0 584 3422 640
rect 3478 584 3483 640
rect 0 582 3483 584
rect 0 552 800 582
rect 3417 579 3483 582
rect 19190 580 19196 644
rect 19260 642 19266 644
rect 22200 642 23000 672
rect 19260 582 23000 642
rect 19260 580 19266 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 1117 234 1183 237
rect 0 232 1183 234
rect 0 176 1122 232
rect 1178 176 1183 232
rect 0 174 1183 176
rect 0 144 800 174
rect 1117 171 1183 174
rect 19241 234 19307 237
rect 22200 234 23000 264
rect 19241 232 23000 234
rect 19241 176 19246 232
rect 19302 176 23000 232
rect 19241 174 23000 176
rect 19241 171 19307 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 9444 18532 9508 18596
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 19012 13364 19076 13428
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 19380 11112 19444 11116
rect 19380 11056 19394 11112
rect 19394 11056 19444 11112
rect 19380 11052 19444 11056
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 19012 10780 19076 10844
rect 19380 10568 19444 10572
rect 19380 10512 19394 10568
rect 19394 10512 19444 10568
rect 19380 10508 19444 10512
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 9444 10024 9508 10028
rect 9444 9968 9494 10024
rect 9494 9968 9508 10024
rect 9444 9964 9508 9968
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 19196 8528 19260 8532
rect 19196 8472 19210 8528
rect 19210 8472 19260 8528
rect 19196 8468 19260 8472
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
rect 19196 580 19260 644
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 9443 18596 9509 18597
rect 9443 18532 9444 18596
rect 9508 18532 9509 18596
rect 9443 18531 9509 18532
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 9446 10029 9506 18531
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 9443 10028 9509 10029
rect 9443 9964 9444 10028
rect 9508 9964 9509 10028
rect 9443 9963 9509 9964
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 19011 13428 19077 13429
rect 19011 13364 19012 13428
rect 19076 13364 19077 13428
rect 19011 13363 19077 13364
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 19014 10845 19074 13363
rect 19379 11116 19445 11117
rect 19379 11052 19380 11116
rect 19444 11052 19445 11116
rect 19379 11051 19445 11052
rect 19011 10844 19077 10845
rect 19011 10780 19012 10844
rect 19076 10780 19077 10844
rect 19011 10779 19077 10780
rect 19382 10573 19442 11051
rect 19379 10572 19445 10573
rect 19379 10508 19380 10572
rect 19444 10508 19445 10572
rect 19379 10507 19445 10508
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 19195 8532 19261 8533
rect 19195 8468 19196 8532
rect 19260 8468 19261 8532
rect 19195 8467 19261 8468
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
rect 19198 645 19258 8467
rect 19195 644 19261 645
rect 19195 580 19196 644
rect 19260 580 19261 644
rect 19195 579 19261 580
use sky130_fd_sc_hd__decap_12  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4692 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608910539
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4784 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1608910539
transform 1 0 5520 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1608910539
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1608910539
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_N_FTB01_A
timestamp 1608910539
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1608910539
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1608910539
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608910539
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1608910539
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608910539
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_164
timestamp 1608910539
transform 1 0 16192 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp 1608910539
transform 1 0 15364 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608910539
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_N_FTB01_A
timestamp 1608910539
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1608910539
transform 1 0 15456 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1608910539
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1608910539
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1608910539
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1608910539
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1608910539
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1608910539
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1608910539
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp 1608910539
transform 1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1608910539
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1608910539
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608910539
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608910539
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608910539
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608910539
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608910539
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1608910539
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1608910539
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608910539
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1608910539
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1608910539
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1608910539
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1608910539
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608910539
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608910539
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608910539
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1608910539
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608910539
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1608910539
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1608910539
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1608910539
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1608910539
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1608910539
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1608910539
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1608910539
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1608910539
transform 1 0 21344 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608910539
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608910539
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608910539
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608910539
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608910539
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1608910539
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1608910539
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1608910539
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1608910539
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1608910539
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1608910539
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1608910539
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1608910539
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608910539
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1608910539
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1608910539
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1608910539
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1608910539
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1608910539
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1608910539
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1608910539
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1608910539
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1608910539
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1608910539
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1608910539
transform 1 0 21344 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608910539
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608910539
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1608910539
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608910539
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1608910539
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1608910539
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1608910539
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1608910539
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1608910539
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1608910539
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1608910539
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1608910539
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1608910539
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1608910539
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1608910539
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1608910539
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1608910539
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1608910539
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1608910539
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1608910539
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1608910539
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1608910539
transform 1 0 19136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1608910539
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1608910539
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1608910539
transform 1 0 21252 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1932 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1608910539
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4784 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_61
timestamp 1608910539
transform 1 0 6716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_49
timestamp 1608910539
transform 1 0 5612 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_73
timestamp 1608910539
transform 1 0 7820 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1608910539
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1608910539
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1608910539
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1608910539
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1608910539
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1608910539
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1608910539
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1608910539
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_202
timestamp 1608910539
transform 1 0 19688 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1608910539
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1608910539
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20424 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2852 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_37
timestamp 1608910539
transform 1 0 4508 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608910539
transform 1 0 4600 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_78
timestamp 1608910539
transform 1 0 8280 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1608910539
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7268 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_102
timestamp 1608910539
transform 1 0 10488 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_90
timestamp 1608910539
transform 1 0 9384 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1608910539
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1608910539
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1608910539
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1608910539
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1608910539
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19136 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1608910539
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1608910539
transform 1 0 20608 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1608910539
transform 1 0 1932 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2024 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1608910539
transform 1 0 4600 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4692 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608910539
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1608910539
transform 1 0 6164 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6532 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8004 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1608910539
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1608910539
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1608910539
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1608910539
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1608910539
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_166
timestamp 1608910539
transform 1 0 16376 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16928 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1608910539
transform 1 0 19228 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_194
timestamp 1608910539
transform 1 0 18952 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_188
timestamp 1608910539
transform 1 0 18400 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19320 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1608910539
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 1932 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2760 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4416 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5244 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_73
timestamp 1608910539
transform 1 0 7820 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8372 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_104
timestamp 1608910539
transform 1 0 10672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_123
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_116
timestamp 1608910539
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_145
timestamp 1608910539
transform 1 0 14444 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_133
timestamp 1608910539
transform 1 0 13340 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_157
timestamp 1608910539
transform 1 0 15548 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1608910539
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1608910539
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16652 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_204
timestamp 1608910539
transform 1 0 19872 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 19964 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18860 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 20792 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1748 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_36
timestamp 1608910539
transform 1 0 4416 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1608910539
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1608910539
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_60
timestamp 1608910539
transform 1 0 6624 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_48
timestamp 1608910539
transform 1 0 5520 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 6716 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_72
timestamp 1608910539
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10580 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9752 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1608910539
transform 1 0 11776 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11868 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_144
timestamp 1608910539
transform 1 0 14352 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_150
timestamp 1608910539
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608910539
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1608910539
transform 1 0 16744 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17112 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_206
timestamp 1608910539
transform 1 0 20056 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 18584 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1608910539
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_210
timestamp 1608910539
transform 1 0 20424 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608910539
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 1472 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _057_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1656 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1608910539
transform 1 0 2852 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2852 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1608910539
transform 1 0 3220 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_35
timestamp 1608910539
transform 1 0 4324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1608910539
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1608910539
transform 1 0 4600 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1608910539
transform 1 0 4508 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608910539
transform 1 0 4232 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_46
timestamp 1608910539
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_47
timestamp 1608910539
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5520 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_83
timestamp 1608910539
transform 1 0 8740 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_64
timestamp 1608910539
transform 1 0 6992 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8464 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7360 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1608910539
transform 1 0 6992 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7820 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608910539
transform 1 0 8188 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1608910539
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1608910539
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_95
timestamp 1608910539
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9936 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_123
timestamp 1608910539
transform 1 0 12420 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1608910539
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608910539
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1608910539
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12512 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_143
timestamp 1608910539
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1608910539
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13892 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1608910539
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 16284 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_186
timestamp 1608910539
transform 1 0 18216 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1608910539
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1608910539
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16744 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1608910539
transform 1 0 20148 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_200
timestamp 1608910539
transform 1 0 19504 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 18492 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 19320 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 20056 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1608910539
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1608910539
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608910539
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1608910539
transform 1 0 3128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3496 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1608910539
transform 1 0 4324 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_55
timestamp 1608910539
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_83
timestamp 1608910539
transform 1 0 8740 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_64
timestamp 1608910539
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7268 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_103
timestamp 1608910539
transform 1 0 10580 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_87
timestamp 1608910539
transform 1 0 9108 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9384 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10856 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1608910539
transform 1 0 13524 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608910539
transform 1 0 13248 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1608910539
transform 1 0 14536 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15732 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_186
timestamp 1608910539
transform 1 0 18216 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_180
timestamp 1608910539
transform 1 0 17664 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1608910539
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_168
timestamp 1608910539
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1608910539
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1608910539
transform 1 0 20424 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608910539
transform 1 0 21252 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1564 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_35
timestamp 1608910539
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_21
timestamp 1608910539
transform 1 0 3036 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1608910539
transform 1 0 4140 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 4508 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_60
timestamp 1608910539
transform 1 0 6624 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1608910539
transform 1 0 8004 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7176 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10672 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12144 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_143
timestamp 1608910539
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_129
timestamp 1608910539
transform 1 0 12972 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13064 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1608910539
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15456 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1608910539
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1608910539
transform 1 0 18216 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1608910539
transform 1 0 17940 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1608910539
transform 1 0 19872 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 19044 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1608910539
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_17
timestamp 1608910539
transform 1 0 2668 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1608910539
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_29
timestamp 1608910539
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3864 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1608910539
transform 1 0 5336 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_65
timestamp 1608910539
transform 1 0 7084 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7452 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_130
timestamp 1608910539
transform 1 0 13064 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1608910539
transform 1 0 12696 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13156 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1608910539
transform 1 0 15732 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 15456 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16468 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_188
timestamp 1608910539
transform 1 0 18400 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 18492 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1608910539
transform 1 0 19320 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1608910539
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20332 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1564 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608910539
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3036 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4876 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_57
timestamp 1608910539
transform 1 0 6348 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1608910539
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7268 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8096 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_95
timestamp 1608910539
transform 1 0 9844 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9936 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1608910539
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12144 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11960 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11592 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10764 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12512 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13984 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1608910539
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 1608910539
transform 1 0 16468 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16560 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_188
timestamp 1608910539
transform 1 0 18400 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 19320 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 18492 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1608910539
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1608910539
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1608910539
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1608910539
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_29
timestamp 1608910539
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_21
timestamp 1608910539
transform 1 0 3036 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_35
timestamp 1608910539
transform 1 0 4324 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_34
timestamp 1608910539
transform 1 0 4232 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 4140 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4600 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_52
timestamp 1608910539
transform 1 0 5888 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1608910539
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608910539
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1608910539
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_53
timestamp 1608910539
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1608910539
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1608910539
transform 1 0 6808 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608910539
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7636 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8464 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1608910539
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1608910539
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_100
timestamp 1608910539
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_95
timestamp 1608910539
transform 1 0 9844 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10488 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9936 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_125
timestamp 1608910539
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1608910539
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11408 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12328 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1608910539
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13800 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13432 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1608910539
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_161
timestamp 1608910539
transform 1 0 15916 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_146
timestamp 1608910539
transform 1 0 14536 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1608910539
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608910539
transform 1 0 15640 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_187
timestamp 1608910539
transform 1 0 18308 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1608910539
transform 1 0 16744 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1608910539
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_173
timestamp 1608910539
transform 1 0 17020 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 16836 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_193
timestamp 1608910539
transform 1 0 18860 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1608910539
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 19136 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 19964 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 19228 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 20056 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1608910539
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1608910539
transform 1 0 21528 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1608910539
transform 1 0 20884 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_17
timestamp 1608910539
transform 1 0 2668 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_25
timestamp 1608910539
transform 1 0 3404 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3496 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1608910539
transform 1 0 4324 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1608910539
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_64
timestamp 1608910539
transform 1 0 6992 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7360 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_96
timestamp 1608910539
transform 1 0 9936 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_84
timestamp 1608910539
transform 1 0 8832 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10856 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13616 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12788 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_147
timestamp 1608910539
transform 1 0 14628 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14904 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15732 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1608910539
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_173
timestamp 1608910539
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608910539
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 19504 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1608910539
transform 1 0 21252 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20332 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608910539
transform 1 0 20884 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608910539
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1608910539
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1608910539
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608910539
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5520 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_64
timestamp 1608910539
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_102
timestamp 1608910539
transform 1 0 10488 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_114
timestamp 1608910539
transform 1 0 11592 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11868 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12696 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1608910539
transform 1 0 15640 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_187
timestamp 1608910539
transform 1 0 18308 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1608910539
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16652 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 19872 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 18400 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1608910539
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1608910539
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1608910539
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1608910539
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1608910539
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1608910539
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3036 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4232 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5888 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7636 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1608910539
transform 1 0 9660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_88
timestamp 1608910539
transform 1 0 9200 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1608910539
transform 1 0 8832 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_105
timestamp 1608910539
transform 1 0 10764 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10856 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608910539
transform 1 0 11684 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_134
timestamp 1608910539
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 13524 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13800 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_158
timestamp 1608910539
transform 1 0 15640 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_154
timestamp 1608910539
transform 1 0 15272 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 15916 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16192 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1608910539
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17020 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_205
timestamp 1608910539
transform 1 0 19964 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_197
timestamp 1608910539
transform 1 0 19228 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20056 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1608910539
transform 1 0 21528 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20608 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608910539
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_19
timestamp 1608910539
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1608910539
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1608910539
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1608910539
transform 1 0 2116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1608910539
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_60
timestamp 1608910539
transform 1 0 6624 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1608910539
transform 1 0 6256 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 5980 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5152 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_73
timestamp 1608910539
transform 1 0 7820 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_65
timestamp 1608910539
transform 1 0 7084 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 7360 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608910539
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608910539
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11960 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1608910539
transform 1 0 11132 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1608910539
transform 1 0 14076 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1608910539
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14168 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608910539
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16100 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17756 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1608910539
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608910539
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608910539
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1608910539
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2576 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1608910539
transform 1 0 2116 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1608910539
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4232 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1608910539
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_52
timestamp 1608910539
transform 1 0 5888 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5060 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_80
timestamp 1608910539
transform 1 0 8464 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 8556 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1608910539
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_88
timestamp 1608910539
transform 1 0 9200 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1608910539
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9292 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10120 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_116
timestamp 1608910539
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13892 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15364 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16836 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608910539
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_188
timestamp 1608910539
transform 1 0 18400 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 20240 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18768 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1608910539
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608910539
transform 1 0 21068 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608910539
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_13
timestamp 1608910539
transform 1 0 2300 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1608910539
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1608910539
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1608910539
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608910539
transform 1 0 2116 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_19
timestamp 1608910539
transform 1 0 2852 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1608910539
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4876 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3036 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4600 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3128 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_62
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1608910539
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_54
timestamp 1608910539
transform 1 0 6072 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_54
timestamp 1608910539
transform 1 0 6072 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6164 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_75
timestamp 1608910539
transform 1 0 8004 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_71
timestamp 1608910539
transform 1 0 7636 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8096 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6900 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_88
timestamp 1608910539
transform 1 0 9200 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9476 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10028 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_106
timestamp 1608910539
transform 1 0 10856 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12512 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11132 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11408 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1608910539
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14076 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13708 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13064 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12880 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1608910539
transform 1 0 14812 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14904 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608910539
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1608910539
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16284 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_158
timestamp 1608910539
transform 1 0 15640 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608910539
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_174
timestamp 1608910539
transform 1 0 17112 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_170
timestamp 1608910539
transform 1 0 16744 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_187
timestamp 1608910539
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17204 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16836 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1608910539
transform 1 0 18492 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19136 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 19320 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1608910539
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1608910539
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608910539
transform 1 0 20792 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1608910539
transform 1 0 21528 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_222
timestamp 1608910539
transform 1 0 21528 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1608910539
transform 1 0 21252 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_19
timestamp 1608910539
transform 1 0 2852 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1608910539
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2300 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4324 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_60
timestamp 1608910539
transform 1 0 6624 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 6716 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5152 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7544 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1608910539
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9752 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_124
timestamp 1608910539
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11224 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1608910539
transform 1 0 12052 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_142
timestamp 1608910539
transform 1 0 14168 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_130
timestamp 1608910539
transform 1 0 13064 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_166
timestamp 1608910539
transform 1 0 16376 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_150
timestamp 1608910539
transform 1 0 14904 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608910539
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_186
timestamp 1608910539
transform 1 0 18216 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_181
timestamp 1608910539
transform 1 0 17756 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17848 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16928 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_198
timestamp 1608910539
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 19504 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1608910539
transform 1 0 19688 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_211
timestamp 1608910539
transform 1 0 20516 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1608910539
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1608910539
transform 1 0 21252 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_17
timestamp 1608910539
transform 1 0 2668 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 1608910539
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1608910539
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1608910539
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608910539
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_41
timestamp 1608910539
transform 1 0 4876 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_29
timestamp 1608910539
transform 1 0 3772 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1608910539
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_50
timestamp 1608910539
transform 1 0 5704 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 5152 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1608910539
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_66
timestamp 1608910539
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8096 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_102
timestamp 1608910539
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_94
timestamp 1608910539
transform 1 0 9752 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10672 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_144
timestamp 1608910539
transform 1 0 14352 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_140
timestamp 1608910539
transform 1 0 13984 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_126
timestamp 1608910539
transform 1 0 12696 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16100 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14628 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1608910539
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608910539
transform 1 0 17572 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_193
timestamp 1608910539
transform 1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 19136 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 19504 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1608910539
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1608910539
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1608910539
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1608910539
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608910539
transform 1 0 20792 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608910539
transform 1 0 20332 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1608910539
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1608910539
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608910539
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608910539
transform 1 0 2116 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608910539
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_26
timestamp 1608910539
transform 1 0 3496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_23
timestamp 1608910539
transform 1 0 3220 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1608910539
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1608910539
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1608910539
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_57
timestamp 1608910539
transform 1 0 6348 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_52
timestamp 1608910539
transform 1 0 5888 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_44
timestamp 1608910539
transform 1 0 5152 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6532 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608910539
transform 1 0 5980 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1608910539
transform 1 0 7084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8740 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608910539
transform 1 0 8372 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 1608910539
transform 1 0 10580 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1608910539
transform 1 0 10212 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10672 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12512 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11684 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_135
timestamp 1608910539
transform 1 0 13524 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13616 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1608910539
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16100 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18308 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16836 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1608910539
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608910539
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608910539
transform 1 0 1472 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608910539
transform 1 0 2944 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608910539
transform 1 0 2576 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608910539
transform 1 0 2208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1608910539
transform 1 0 1840 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_29
timestamp 1608910539
transform 1 0 3772 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_24
timestamp 1608910539
transform 1 0 3312 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3864 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608910539
transform 1 0 3404 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_62
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608910539
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_52
timestamp 1608910539
transform 1 0 5888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_44
timestamp 1608910539
transform 1 0 5152 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608910539
transform 1 0 6164 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_70
timestamp 1608910539
transform 1 0 7544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7636 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9108 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608910539
transform 1 0 10580 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12512 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10856 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14812 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1608910539
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16468 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608910539
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608910539
transform 1 0 17020 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_193
timestamp 1608910539
transform 1 0 18860 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18952 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1608910539
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608910539
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608910539
transform 1 0 21160 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608910539
transform 1 0 20792 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1608910539
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608910539
transform 1 0 1472 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608910539
transform 1 0 2576 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608910539
transform 1 0 2208 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608910539
transform 1 0 1840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1608910539
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_24
timestamp 1608910539
transform 1 0 3312 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1608910539
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1608910539
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608910539
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_80
timestamp 1608910539
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1608910539
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9844 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_111
timestamp 1608910539
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12328 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_132
timestamp 1608910539
transform 1 0 13248 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13524 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608910539
transform 1 0 12880 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608910539
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1608910539
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1608910539
transform 1 0 15640 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16100 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608910539
transform 1 0 14720 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1608910539
transform 1 0 18124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1608910539
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17572 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608910539
transform 1 0 18216 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608910539
transform 1 0 17020 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608910539
transform 1 0 16652 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19780 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18952 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608910539
transform 1 0 18584 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 1608910539
transform 1 0 20332 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608910539
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608910539
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_14
timestamp 1608910539
transform 1 0 2392 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_9
timestamp 1608910539
transform 1 0 1932 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_5
timestamp 1608910539
transform 1 0 1564 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1608910539
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1608910539
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_30
timestamp 1608910539
transform 1 0 3864 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_26
timestamp 1608910539
transform 1 0 3496 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1608910539
transform 1 0 6256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1608910539
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_75
timestamp 1608910539
transform 1 0 8004 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8740 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_92
timestamp 1608910539
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_182
timestamp 1608910539
transform 1 0 17848 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608910539
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608910539
transform 1 0 17112 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_207
timestamp 1608910539
transform 1 0 20148 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_201
timestamp 1608910539
transform 1 0 19596 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1608910539
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1608910539
transform 1 0 20240 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608910539
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1608910539
transform 1 0 21528 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1608910539
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_210
timestamp 1608910539
transform 1 0 20424 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1608910539
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
<< labels >>
rlabel metal2 s 202 22200 258 23000 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 SC_OUT_TOP
port 1 nsew signal tristate
rlabel metal2 s 4434 22200 4490 23000 6 Test_en_N_out
port 2 nsew signal tristate
rlabel metal2 s 20718 0 20774 800 6 Test_en_S_in
port 3 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 ccff_head
port 4 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 ccff_tail
port 5 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[0]
port 6 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 7 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 8 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 9 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 10 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[14]
port 11 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 12 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 13 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 14 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[18]
port 15 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 16 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 17 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 18 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 19 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 20 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 21 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 22 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[7]
port 23 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 24 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 25 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 26 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[10]
port 27 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 28 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[12]
port 29 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 30 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[14]
port 31 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 32 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[16]
port 33 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 34 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[18]
port 35 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 36 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 37 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 38 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[3]
port 39 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 40 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[5]
port 41 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 42 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[7]
port 43 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[8]
port 44 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[9]
port 45 nsew signal tristate
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[0]
port 46 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[10]
port 47 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[11]
port 48 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[12]
port 49 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[13]
port 50 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[14]
port 51 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[15]
port 52 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[16]
port 53 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[17]
port 54 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[18]
port 55 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_in[19]
port 56 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[1]
port 57 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[2]
port 58 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[3]
port 59 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[4]
port 60 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[5]
port 61 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[6]
port 62 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[7]
port 63 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[8]
port 64 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[9]
port 65 nsew signal input
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[0]
port 66 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[10]
port 67 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[11]
port 68 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[12]
port 69 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[13]
port 70 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[14]
port 71 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[15]
port 72 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[16]
port 73 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[17]
port 74 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[18]
port 75 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 chanx_right_out[19]
port 76 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[1]
port 77 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[2]
port 78 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[3]
port 79 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[4]
port 80 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[5]
port 81 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[6]
port 82 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[7]
port 83 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[8]
port 84 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[9]
port 85 nsew signal tristate
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[0]
port 86 nsew signal input
rlabel metal2 s 9954 22200 10010 23000 6 chany_top_in[10]
port 87 nsew signal input
rlabel metal2 s 10414 22200 10470 23000 6 chany_top_in[11]
port 88 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[12]
port 89 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[13]
port 90 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[14]
port 91 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_in[15]
port 92 nsew signal input
rlabel metal2 s 12530 22200 12586 23000 6 chany_top_in[16]
port 93 nsew signal input
rlabel metal2 s 12898 22200 12954 23000 6 chany_top_in[17]
port 94 nsew signal input
rlabel metal2 s 13358 22200 13414 23000 6 chany_top_in[18]
port 95 nsew signal input
rlabel metal2 s 13818 22200 13874 23000 6 chany_top_in[19]
port 96 nsew signal input
rlabel metal2 s 6090 22200 6146 23000 6 chany_top_in[1]
port 97 nsew signal input
rlabel metal2 s 6550 22200 6606 23000 6 chany_top_in[2]
port 98 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[3]
port 99 nsew signal input
rlabel metal2 s 7378 22200 7434 23000 6 chany_top_in[4]
port 100 nsew signal input
rlabel metal2 s 7838 22200 7894 23000 6 chany_top_in[5]
port 101 nsew signal input
rlabel metal2 s 8206 22200 8262 23000 6 chany_top_in[6]
port 102 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[7]
port 103 nsew signal input
rlabel metal2 s 9126 22200 9182 23000 6 chany_top_in[8]
port 104 nsew signal input
rlabel metal2 s 9494 22200 9550 23000 6 chany_top_in[9]
port 105 nsew signal input
rlabel metal2 s 14186 22200 14242 23000 6 chany_top_out[0]
port 106 nsew signal tristate
rlabel metal2 s 18510 22200 18566 23000 6 chany_top_out[10]
port 107 nsew signal tristate
rlabel metal2 s 18878 22200 18934 23000 6 chany_top_out[11]
port 108 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[12]
port 109 nsew signal tristate
rlabel metal2 s 19706 22200 19762 23000 6 chany_top_out[13]
port 110 nsew signal tristate
rlabel metal2 s 20166 22200 20222 23000 6 chany_top_out[14]
port 111 nsew signal tristate
rlabel metal2 s 20626 22200 20682 23000 6 chany_top_out[15]
port 112 nsew signal tristate
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 113 nsew signal tristate
rlabel metal2 s 21454 22200 21510 23000 6 chany_top_out[17]
port 114 nsew signal tristate
rlabel metal2 s 21914 22200 21970 23000 6 chany_top_out[18]
port 115 nsew signal tristate
rlabel metal2 s 22282 22200 22338 23000 6 chany_top_out[19]
port 116 nsew signal tristate
rlabel metal2 s 14646 22200 14702 23000 6 chany_top_out[1]
port 117 nsew signal tristate
rlabel metal2 s 15106 22200 15162 23000 6 chany_top_out[2]
port 118 nsew signal tristate
rlabel metal2 s 15474 22200 15530 23000 6 chany_top_out[3]
port 119 nsew signal tristate
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[4]
port 120 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[5]
port 121 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[6]
port 122 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[7]
port 123 nsew signal tristate
rlabel metal2 s 17590 22200 17646 23000 6 chany_top_out[8]
port 124 nsew signal tristate
rlabel metal2 s 18050 22200 18106 23000 6 chany_top_out[9]
port 125 nsew signal tristate
rlabel metal2 s 4802 22200 4858 23000 6 clk_3_N_out
port 126 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 clk_3_S_in
port 127 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 128 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 129 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 130 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 131 nsew signal input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 132 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 133 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 134 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 135 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 136 nsew signal input
rlabel metal2 s 3974 22200 4030 23000 6 prog_clk_0_N_in
port 137 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 prog_clk_3_N_out
port 138 nsew signal tristate
rlabel metal2 s 11518 0 11574 800 6 prog_clk_3_S_in
port 139 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_11_
port 140 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_13_
port 141 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_15_
port 142 nsew signal input
rlabel metal3 s 22200 3816 23000 3936 6 right_bottom_grid_pin_17_
port 143 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_1_
port 144 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_3_
port 145 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_5_
port 146 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_7_
port 147 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_9_
port 148 nsew signal input
rlabel metal2 s 570 22200 626 23000 6 top_left_grid_pin_42_
port 149 nsew signal input
rlabel metal2 s 1030 22200 1086 23000 6 top_left_grid_pin_43_
port 150 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 top_left_grid_pin_44_
port 151 nsew signal input
rlabel metal2 s 1858 22200 1914 23000 6 top_left_grid_pin_45_
port 152 nsew signal input
rlabel metal2 s 2318 22200 2374 23000 6 top_left_grid_pin_46_
port 153 nsew signal input
rlabel metal2 s 2686 22200 2742 23000 6 top_left_grid_pin_47_
port 154 nsew signal input
rlabel metal2 s 3146 22200 3202 23000 6 top_left_grid_pin_48_
port 155 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 top_left_grid_pin_49_
port 156 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 157 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 158 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 159 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 160 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 161 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
