magic
tech sky130A
magscale 1 2
timestamp 1605198840
<< locali >>
rect 11805 19771 11839 19941
rect 2513 19295 2547 19397
rect 12265 19295 12299 19465
rect 2789 18683 2823 18785
rect 6653 18615 6687 18717
rect 12265 18071 12299 18309
rect 4353 17187 4387 17289
rect 19349 17051 19383 17153
rect 22017 16779 22051 17833
rect 3065 15895 3099 16201
rect 2697 15419 2731 15521
rect 8585 15419 8619 15589
rect 11161 15419 11195 15657
rect 16497 15351 16531 15521
rect 18153 15351 18187 15453
rect 20085 15351 20119 15521
rect 18095 15317 18187 15351
rect 6653 14399 6687 14501
rect 4997 12699 5031 12869
rect 11989 12155 12023 12325
rect 15393 12087 15427 12189
rect 7665 11203 7699 11305
rect 9413 10999 9447 11237
rect 14565 11203 14599 11305
rect 9413 9027 9447 9061
rect 9689 9027 9723 9129
rect 9413 8993 9723 9027
rect 18889 8823 18923 8993
rect 9965 8347 9999 8517
rect 10517 7191 10551 7429
rect 12173 7191 12207 7361
rect 16957 6715 16991 6953
rect 16865 5559 16899 5729
rect 12173 5015 12207 5185
rect 14105 5083 14139 5253
rect 17417 4607 17451 4777
rect 10333 3927 10367 4165
rect 17785 3927 17819 4029
rect 2881 3451 2915 3621
rect 17877 2941 17969 2975
rect 17877 2839 17911 2941
<< viali >>
rect 1961 20553 1995 20587
rect 2513 20553 2547 20587
rect 5825 20553 5859 20587
rect 15025 20553 15059 20587
rect 15945 20553 15979 20587
rect 16681 20553 16715 20587
rect 19533 20553 19567 20587
rect 20729 20553 20763 20587
rect 10333 20485 10367 20519
rect 12633 20485 12667 20519
rect 20177 20485 20211 20519
rect 6377 20417 6411 20451
rect 8033 20417 8067 20451
rect 9045 20417 9079 20451
rect 10793 20417 10827 20451
rect 10977 20417 11011 20451
rect 11897 20417 11931 20451
rect 13277 20417 13311 20451
rect 1777 20349 1811 20383
rect 2329 20349 2363 20383
rect 4077 20349 4111 20383
rect 4344 20349 4378 20383
rect 11713 20349 11747 20383
rect 13645 20349 13679 20383
rect 14841 20349 14875 20383
rect 15761 20349 15795 20383
rect 16497 20349 16531 20383
rect 19349 20349 19383 20383
rect 19993 20349 20027 20383
rect 20545 20349 20579 20383
rect 7757 20281 7791 20315
rect 8769 20281 8803 20315
rect 13093 20281 13127 20315
rect 13921 20281 13955 20315
rect 5457 20213 5491 20247
rect 6193 20213 6227 20247
rect 6285 20213 6319 20247
rect 7389 20213 7423 20247
rect 7849 20213 7883 20247
rect 8401 20213 8435 20247
rect 8861 20213 8895 20247
rect 10701 20213 10735 20247
rect 11345 20213 11379 20247
rect 11805 20213 11839 20247
rect 13001 20213 13035 20247
rect 1961 20009 1995 20043
rect 3065 20009 3099 20043
rect 7389 20009 7423 20043
rect 9045 20009 9079 20043
rect 9873 20009 9907 20043
rect 14841 20009 14875 20043
rect 16497 20009 16531 20043
rect 17785 20009 17819 20043
rect 18797 20009 18831 20043
rect 19901 20009 19935 20043
rect 20453 20009 20487 20043
rect 21097 20009 21131 20043
rect 4620 19941 4654 19975
rect 6276 19941 6310 19975
rect 7932 19941 7966 19975
rect 10600 19941 10634 19975
rect 11805 19941 11839 19975
rect 12256 19941 12290 19975
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 2881 19873 2915 19907
rect 6009 19873 6043 19907
rect 9689 19873 9723 19907
rect 10333 19873 10367 19907
rect 4353 19805 4387 19839
rect 7665 19805 7699 19839
rect 14013 19873 14047 19907
rect 14657 19873 14691 19907
rect 15577 19873 15611 19907
rect 15853 19873 15887 19907
rect 16313 19873 16347 19907
rect 16865 19873 16899 19907
rect 17601 19873 17635 19907
rect 18613 19873 18647 19907
rect 19165 19873 19199 19907
rect 19717 19873 19751 19907
rect 20269 19873 20303 19907
rect 20913 19873 20947 19907
rect 21281 19873 21315 19907
rect 11989 19805 12023 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 11713 19737 11747 19771
rect 11805 19737 11839 19771
rect 13645 19737 13679 19771
rect 17049 19737 17083 19771
rect 19349 19737 19383 19771
rect 2513 19669 2547 19703
rect 5733 19669 5767 19703
rect 13369 19669 13403 19703
rect 5733 19465 5767 19499
rect 8493 19465 8527 19499
rect 10977 19465 11011 19499
rect 12265 19465 12299 19499
rect 13829 19465 13863 19499
rect 21005 19465 21039 19499
rect 2513 19397 2547 19431
rect 3249 19329 3283 19363
rect 4169 19329 4203 19363
rect 5273 19329 5307 19363
rect 6377 19329 6411 19363
rect 9137 19329 9171 19363
rect 11805 19329 11839 19363
rect 11989 19329 12023 19363
rect 14657 19329 14691 19363
rect 1777 19261 1811 19295
rect 2513 19261 2547 19295
rect 5089 19261 5123 19295
rect 6837 19261 6871 19295
rect 8953 19261 8987 19295
rect 9597 19261 9631 19295
rect 12265 19261 12299 19295
rect 12449 19261 12483 19295
rect 12705 19261 12739 19295
rect 14473 19261 14507 19295
rect 15117 19261 15151 19295
rect 15393 19261 15427 19295
rect 15945 19261 15979 19295
rect 16221 19261 16255 19295
rect 16681 19261 16715 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 19165 19261 19199 19295
rect 19717 19261 19751 19295
rect 20269 19261 20303 19295
rect 20821 19261 20855 19295
rect 3065 19193 3099 19227
rect 4997 19193 5031 19227
rect 6193 19193 6227 19227
rect 7104 19193 7138 19227
rect 9864 19193 9898 19227
rect 14565 19193 14599 19227
rect 1961 19125 1995 19159
rect 2605 19125 2639 19159
rect 2973 19125 3007 19159
rect 3617 19125 3651 19159
rect 3985 19125 4019 19159
rect 4077 19125 4111 19159
rect 4629 19125 4663 19159
rect 6101 19125 6135 19159
rect 8217 19125 8251 19159
rect 8861 19125 8895 19159
rect 11345 19125 11379 19159
rect 11713 19125 11747 19159
rect 14105 19125 14139 19159
rect 16865 19125 16899 19159
rect 17601 19125 17635 19159
rect 18245 19125 18279 19159
rect 19349 19125 19383 19159
rect 19901 19125 19935 19159
rect 20453 19125 20487 19159
rect 1869 18921 1903 18955
rect 2973 18921 3007 18955
rect 3341 18921 3375 18955
rect 4537 18921 4571 18955
rect 5733 18921 5767 18955
rect 6193 18921 6227 18955
rect 6929 18921 6963 18955
rect 9689 18921 9723 18955
rect 11161 18921 11195 18955
rect 14381 18921 14415 18955
rect 18521 18921 18555 18955
rect 21097 18921 21131 18955
rect 2513 18853 2547 18887
rect 4445 18853 4479 18887
rect 12532 18853 12566 18887
rect 1685 18785 1719 18819
rect 2237 18785 2271 18819
rect 2789 18785 2823 18819
rect 5089 18785 5123 18819
rect 6101 18785 6135 18819
rect 7297 18785 7331 18819
rect 8769 18785 8803 18819
rect 10057 18785 10091 18819
rect 11069 18785 11103 18819
rect 11713 18785 11747 18819
rect 14289 18785 14323 18819
rect 17233 18785 17267 18819
rect 17509 18785 17543 18819
rect 18337 18785 18371 18819
rect 19717 18785 19751 18819
rect 20269 18785 20303 18819
rect 20913 18785 20947 18819
rect 3433 18717 3467 18751
rect 3617 18717 3651 18751
rect 4629 18717 4663 18751
rect 5365 18717 5399 18751
rect 6377 18717 6411 18751
rect 6653 18717 6687 18751
rect 7389 18717 7423 18751
rect 7573 18717 7607 18751
rect 7941 18717 7975 18751
rect 8861 18717 8895 18751
rect 9045 18717 9079 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 11253 18717 11287 18751
rect 12265 18717 12299 18751
rect 14473 18717 14507 18751
rect 2789 18649 2823 18683
rect 10701 18649 10735 18683
rect 13645 18649 13679 18683
rect 13921 18649 13955 18683
rect 19901 18649 19935 18683
rect 4077 18581 4111 18615
rect 6653 18581 6687 18615
rect 6745 18581 6779 18615
rect 8401 18581 8435 18615
rect 11897 18581 11931 18615
rect 20453 18581 20487 18615
rect 1961 18377 1995 18411
rect 2513 18377 2547 18411
rect 2881 18377 2915 18411
rect 5549 18377 5583 18411
rect 6837 18377 6871 18411
rect 7941 18377 7975 18411
rect 9045 18377 9079 18411
rect 11069 18377 11103 18411
rect 12541 18377 12575 18411
rect 13553 18377 13587 18411
rect 14749 18377 14783 18411
rect 21281 18377 21315 18411
rect 5273 18309 5307 18343
rect 12265 18309 12299 18343
rect 3341 18241 3375 18275
rect 3525 18241 3559 18275
rect 6101 18241 6135 18275
rect 7481 18241 7515 18275
rect 8493 18241 8527 18275
rect 9689 18241 9723 18275
rect 10701 18241 10735 18275
rect 11621 18241 11655 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 3893 18173 3927 18207
rect 7205 18173 7239 18207
rect 8309 18173 8343 18207
rect 4160 18105 4194 18139
rect 6009 18105 6043 18139
rect 9413 18105 9447 18139
rect 11437 18105 11471 18139
rect 13185 18241 13219 18275
rect 14013 18241 14047 18275
rect 14197 18241 14231 18275
rect 16865 18241 16899 18275
rect 18889 18241 18923 18275
rect 19073 18241 19107 18275
rect 19809 18241 19843 18275
rect 20637 18241 20671 18275
rect 14565 18173 14599 18207
rect 18797 18173 18831 18207
rect 19625 18173 19659 18207
rect 20361 18173 20395 18207
rect 21097 18173 21131 18207
rect 13001 18105 13035 18139
rect 15117 18105 15151 18139
rect 16681 18105 16715 18139
rect 3249 18037 3283 18071
rect 5917 18037 5951 18071
rect 7297 18037 7331 18071
rect 7665 18037 7699 18071
rect 8401 18037 8435 18071
rect 9505 18037 9539 18071
rect 10057 18037 10091 18071
rect 10425 18037 10459 18071
rect 10517 18037 10551 18071
rect 11529 18037 11563 18071
rect 12265 18037 12299 18071
rect 12909 18037 12943 18071
rect 13921 18037 13955 18071
rect 16313 18037 16347 18071
rect 16773 18037 16807 18071
rect 18429 18037 18463 18071
rect 1593 17833 1627 17867
rect 2973 17833 3007 17867
rect 3433 17833 3467 17867
rect 4537 17833 4571 17867
rect 7481 17833 7515 17867
rect 7849 17833 7883 17867
rect 11069 17833 11103 17867
rect 11345 17833 11379 17867
rect 11713 17833 11747 17867
rect 12449 17833 12483 17867
rect 13461 17833 13495 17867
rect 13829 17833 13863 17867
rect 16313 17833 16347 17867
rect 17877 17833 17911 17867
rect 21097 17833 21131 17867
rect 22017 17833 22051 17867
rect 2237 17765 2271 17799
rect 4445 17765 4479 17799
rect 5632 17765 5666 17799
rect 12909 17765 12943 17799
rect 17969 17765 18003 17799
rect 18981 17765 19015 17799
rect 20177 17765 20211 17799
rect 1409 17697 1443 17731
rect 1950 17697 1984 17731
rect 3341 17697 3375 17731
rect 8861 17697 8895 17731
rect 8953 17697 8987 17731
rect 9945 17697 9979 17731
rect 12817 17697 12851 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 16681 17697 16715 17731
rect 16773 17697 16807 17731
rect 18889 17697 18923 17731
rect 20913 17697 20947 17731
rect 3525 17629 3559 17663
rect 4629 17629 4663 17663
rect 5365 17629 5399 17663
rect 7941 17629 7975 17663
rect 8125 17629 8159 17663
rect 9137 17629 9171 17663
rect 9689 17629 9723 17663
rect 11805 17629 11839 17663
rect 11897 17629 11931 17663
rect 13093 17629 13127 17663
rect 13921 17629 13955 17663
rect 14013 17629 14047 17663
rect 15853 17629 15887 17663
rect 16957 17629 16991 17663
rect 18061 17629 18095 17663
rect 19073 17629 19107 17663
rect 20269 17629 20303 17663
rect 20453 17629 20487 17663
rect 4077 17561 4111 17595
rect 15301 17561 15335 17595
rect 18521 17561 18555 17595
rect 6745 17493 6779 17527
rect 8493 17493 8527 17527
rect 17509 17493 17543 17527
rect 19809 17493 19843 17527
rect 1961 17289 1995 17323
rect 4169 17289 4203 17323
rect 4353 17289 4387 17323
rect 4445 17289 4479 17323
rect 5733 17289 5767 17323
rect 7021 17289 7055 17323
rect 9413 17289 9447 17323
rect 10701 17289 10735 17323
rect 15577 17289 15611 17323
rect 16865 17289 16899 17323
rect 18429 17289 18463 17323
rect 2789 17153 2823 17187
rect 4353 17153 4387 17187
rect 4997 17153 5031 17187
rect 6193 17153 6227 17187
rect 6377 17153 6411 17187
rect 7573 17153 7607 17187
rect 8033 17153 8067 17187
rect 10149 17153 10183 17187
rect 10241 17153 10275 17187
rect 11345 17153 11379 17187
rect 11713 17153 11747 17187
rect 16405 17153 16439 17187
rect 17325 17153 17359 17187
rect 17417 17153 17451 17187
rect 18889 17153 18923 17187
rect 18981 17153 19015 17187
rect 19349 17153 19383 17187
rect 19901 17153 19935 17187
rect 19993 17153 20027 17187
rect 21005 17153 21039 17187
rect 1777 17085 1811 17119
rect 3056 17085 3090 17119
rect 11069 17085 11103 17119
rect 12449 17085 12483 17119
rect 12716 17085 12750 17119
rect 14197 17085 14231 17119
rect 16221 17085 16255 17119
rect 20913 17085 20947 17119
rect 6101 17017 6135 17051
rect 7481 17017 7515 17051
rect 8300 17017 8334 17051
rect 14464 17017 14498 17051
rect 16313 17017 16347 17051
rect 17233 17017 17267 17051
rect 19349 17017 19383 17051
rect 4813 16949 4847 16983
rect 4905 16949 4939 16983
rect 7389 16949 7423 16983
rect 9689 16949 9723 16983
rect 10057 16949 10091 16983
rect 11161 16949 11195 16983
rect 13829 16949 13863 16983
rect 15853 16949 15887 16983
rect 18797 16949 18831 16983
rect 19441 16949 19475 16983
rect 19809 16949 19843 16983
rect 20453 16949 20487 16983
rect 20821 16949 20855 16983
rect 1593 16745 1627 16779
rect 2329 16745 2363 16779
rect 2973 16745 3007 16779
rect 4353 16745 4387 16779
rect 6653 16745 6687 16779
rect 10885 16745 10919 16779
rect 11897 16745 11931 16779
rect 15301 16745 15335 16779
rect 15669 16745 15703 16779
rect 15761 16745 15795 16779
rect 16313 16745 16347 16779
rect 16773 16745 16807 16779
rect 17325 16745 17359 16779
rect 17693 16745 17727 16779
rect 18337 16745 18371 16779
rect 19349 16745 19383 16779
rect 21097 16745 21131 16779
rect 22017 16745 22051 16779
rect 2421 16677 2455 16711
rect 4813 16677 4847 16711
rect 6561 16677 6595 16711
rect 8024 16677 8058 16711
rect 10333 16677 10367 16711
rect 11345 16677 11379 16711
rect 12265 16677 12299 16711
rect 17785 16677 17819 16711
rect 18705 16677 18739 16711
rect 18797 16677 18831 16711
rect 19809 16677 19843 16711
rect 1409 16609 1443 16643
rect 3341 16609 3375 16643
rect 4721 16609 4755 16643
rect 7757 16609 7791 16643
rect 10241 16609 10275 16643
rect 11253 16609 11287 16643
rect 13360 16609 13394 16643
rect 14749 16609 14783 16643
rect 16681 16609 16715 16643
rect 19717 16609 19751 16643
rect 20913 16609 20947 16643
rect 2605 16541 2639 16575
rect 3433 16541 3467 16575
rect 3617 16541 3651 16575
rect 4905 16541 4939 16575
rect 6745 16541 6779 16575
rect 10517 16541 10551 16575
rect 11437 16541 11471 16575
rect 12357 16541 12391 16575
rect 12449 16541 12483 16575
rect 13093 16541 13127 16575
rect 15853 16541 15887 16575
rect 16865 16541 16899 16575
rect 17877 16541 17911 16575
rect 18889 16541 18923 16575
rect 19901 16541 19935 16575
rect 14473 16473 14507 16507
rect 1961 16405 1995 16439
rect 6193 16405 6227 16439
rect 9137 16405 9171 16439
rect 9873 16405 9907 16439
rect 16129 16405 16163 16439
rect 3065 16201 3099 16235
rect 4537 16201 4571 16235
rect 5733 16201 5767 16235
rect 8769 16201 8803 16235
rect 13829 16201 13863 16235
rect 14105 16201 14139 16235
rect 16865 16201 16899 16235
rect 20361 16201 20395 16235
rect 1593 16133 1627 16167
rect 2145 16133 2179 16167
rect 2789 16065 2823 16099
rect 1409 15997 1443 16031
rect 2053 15929 2087 15963
rect 2605 15929 2639 15963
rect 8309 16133 8343 16167
rect 19349 16133 19383 16167
rect 6377 16065 6411 16099
rect 6929 16065 6963 16099
rect 9321 16065 9355 16099
rect 10333 16065 10367 16099
rect 11437 16065 11471 16099
rect 14565 16065 14599 16099
rect 14749 16065 14783 16099
rect 17417 16065 17451 16099
rect 18613 16065 18647 16099
rect 19993 16065 20027 16099
rect 20821 16065 20855 16099
rect 20913 16065 20947 16099
rect 3157 15997 3191 16031
rect 6101 15997 6135 16031
rect 7196 15997 7230 16031
rect 9137 15997 9171 16031
rect 11161 15997 11195 16031
rect 12449 15997 12483 16031
rect 14473 15997 14507 16031
rect 15209 15997 15243 16031
rect 15476 15997 15510 16031
rect 17233 15997 17267 16031
rect 18429 15997 18463 16031
rect 20729 15997 20763 16031
rect 3424 15929 3458 15963
rect 10149 15929 10183 15963
rect 12716 15929 12750 15963
rect 18521 15929 18555 15963
rect 2513 15861 2547 15895
rect 3065 15861 3099 15895
rect 4813 15861 4847 15895
rect 6193 15861 6227 15895
rect 8677 15861 8711 15895
rect 9229 15861 9263 15895
rect 9781 15861 9815 15895
rect 10241 15861 10275 15895
rect 10793 15861 10827 15895
rect 11253 15861 11287 15895
rect 16589 15861 16623 15895
rect 17325 15861 17359 15895
rect 18061 15861 18095 15895
rect 19717 15861 19751 15895
rect 19809 15861 19843 15895
rect 1685 15657 1719 15691
rect 2881 15657 2915 15691
rect 2973 15657 3007 15691
rect 3433 15657 3467 15691
rect 4077 15657 4111 15691
rect 4445 15657 4479 15691
rect 8493 15657 8527 15691
rect 10241 15657 10275 15691
rect 10609 15657 10643 15691
rect 10701 15657 10735 15691
rect 11161 15657 11195 15691
rect 12909 15657 12943 15691
rect 14381 15657 14415 15691
rect 15301 15657 15335 15691
rect 18705 15657 18739 15691
rect 20453 15657 20487 15691
rect 2329 15589 2363 15623
rect 8585 15589 8619 15623
rect 9045 15589 9079 15623
rect 1501 15521 1535 15555
rect 2053 15521 2087 15555
rect 2697 15521 2731 15555
rect 3341 15521 3375 15555
rect 4537 15521 4571 15555
rect 5713 15521 5747 15555
rect 7113 15521 7147 15555
rect 7380 15521 7414 15555
rect 3525 15453 3559 15487
rect 4629 15453 4663 15487
rect 5457 15453 5491 15487
rect 8769 15521 8803 15555
rect 10793 15453 10827 15487
rect 2697 15385 2731 15419
rect 6837 15385 6871 15419
rect 8585 15385 8619 15419
rect 13369 15589 13403 15623
rect 14289 15589 14323 15623
rect 15669 15589 15703 15623
rect 16856 15589 16890 15623
rect 19717 15589 19751 15623
rect 11253 15521 11287 15555
rect 11520 15521 11554 15555
rect 13277 15521 13311 15555
rect 16497 15521 16531 15555
rect 16589 15521 16623 15555
rect 18613 15521 18647 15555
rect 19625 15521 19659 15555
rect 20085 15521 20119 15555
rect 20269 15521 20303 15555
rect 20913 15521 20947 15555
rect 13461 15453 13495 15487
rect 14473 15453 14507 15487
rect 15761 15453 15795 15487
rect 15945 15453 15979 15487
rect 11161 15385 11195 15419
rect 13921 15385 13955 15419
rect 18153 15453 18187 15487
rect 18797 15453 18831 15487
rect 19901 15453 19935 15487
rect 18245 15385 18279 15419
rect 21097 15453 21131 15487
rect 12633 15317 12667 15351
rect 16497 15317 16531 15351
rect 17969 15317 18003 15351
rect 18061 15317 18095 15351
rect 19257 15317 19291 15351
rect 20085 15317 20119 15351
rect 1869 15113 1903 15147
rect 3249 15113 3283 15147
rect 7941 15113 7975 15147
rect 11897 15113 11931 15147
rect 12449 15113 12483 15147
rect 13461 15113 13495 15147
rect 14105 15113 14139 15147
rect 15485 15113 15519 15147
rect 19441 15113 19475 15147
rect 21005 15113 21039 15147
rect 4261 15045 4295 15079
rect 10149 15045 10183 15079
rect 3801 14977 3835 15011
rect 4905 14977 4939 15011
rect 5733 14977 5767 15011
rect 5917 14977 5951 15011
rect 7389 14977 7423 15011
rect 8493 14977 8527 15011
rect 9689 14977 9723 15011
rect 13001 14977 13035 15011
rect 14657 14977 14691 15011
rect 20361 14977 20395 15011
rect 1685 14909 1719 14943
rect 2237 14909 2271 14943
rect 6469 14909 6503 14943
rect 7205 14909 7239 14943
rect 8309 14909 8343 14943
rect 8401 14909 8435 14943
rect 10333 14909 10367 14943
rect 10517 14909 10551 14943
rect 10784 14909 10818 14943
rect 12817 14909 12851 14943
rect 13645 14909 13679 14943
rect 15301 14909 15335 14943
rect 15853 14909 15887 14943
rect 16120 14909 16154 14943
rect 18061 14909 18095 14943
rect 20177 14909 20211 14943
rect 20821 14909 20855 14943
rect 2513 14841 2547 14875
rect 3157 14841 3191 14875
rect 5641 14841 5675 14875
rect 9045 14841 9079 14875
rect 9597 14841 9631 14875
rect 18328 14841 18362 14875
rect 20085 14841 20119 14875
rect 3617 14773 3651 14807
rect 3709 14773 3743 14807
rect 4629 14773 4663 14807
rect 4721 14773 4755 14807
rect 5273 14773 5307 14807
rect 6285 14773 6319 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 9137 14773 9171 14807
rect 9505 14773 9539 14807
rect 12909 14773 12943 14807
rect 14473 14773 14507 14807
rect 14565 14773 14599 14807
rect 17233 14773 17267 14807
rect 17509 14773 17543 14807
rect 19717 14773 19751 14807
rect 1961 14569 1995 14603
rect 3525 14569 3559 14603
rect 7205 14569 7239 14603
rect 8953 14569 8987 14603
rect 11805 14569 11839 14603
rect 15301 14569 15335 14603
rect 16773 14569 16807 14603
rect 18797 14569 18831 14603
rect 19257 14569 19291 14603
rect 19809 14569 19843 14603
rect 21097 14569 21131 14603
rect 2789 14501 2823 14535
rect 4344 14501 4378 14535
rect 6653 14501 6687 14535
rect 8309 14501 8343 14535
rect 10416 14501 10450 14535
rect 14473 14501 14507 14535
rect 15669 14501 15703 14535
rect 15761 14501 15795 14535
rect 18245 14501 18279 14535
rect 19165 14501 19199 14535
rect 1777 14433 1811 14467
rect 2697 14433 2731 14467
rect 3341 14433 3375 14467
rect 6101 14433 6135 14467
rect 7113 14433 7147 14467
rect 8401 14433 8435 14467
rect 10149 14433 10183 14467
rect 12173 14433 12207 14467
rect 13369 14433 13403 14467
rect 14381 14433 14415 14467
rect 16681 14433 16715 14467
rect 18153 14433 18187 14467
rect 20177 14433 20211 14467
rect 20913 14433 20947 14467
rect 2973 14365 3007 14399
rect 4077 14365 4111 14399
rect 6193 14365 6227 14399
rect 6377 14365 6411 14399
rect 6653 14365 6687 14399
rect 7297 14365 7331 14399
rect 8493 14365 8527 14399
rect 12265 14365 12299 14399
rect 12449 14365 12483 14399
rect 13461 14365 13495 14399
rect 13553 14365 13587 14399
rect 14565 14365 14599 14399
rect 15853 14365 15887 14399
rect 16865 14365 16899 14399
rect 18429 14365 18463 14399
rect 19349 14365 19383 14399
rect 20269 14365 20303 14399
rect 20361 14365 20395 14399
rect 11529 14297 11563 14331
rect 2329 14229 2363 14263
rect 5457 14229 5491 14263
rect 5733 14229 5767 14263
rect 6745 14229 6779 14263
rect 7941 14229 7975 14263
rect 13001 14229 13035 14263
rect 14013 14229 14047 14263
rect 16313 14229 16347 14263
rect 17785 14229 17819 14263
rect 1593 14025 1627 14059
rect 4445 14025 4479 14059
rect 6101 14025 6135 14059
rect 6469 14025 6503 14059
rect 11161 14025 11195 14059
rect 13093 14025 13127 14059
rect 16589 14025 16623 14059
rect 16865 14025 16899 14059
rect 20085 14025 20119 14059
rect 8493 13957 8527 13991
rect 9137 13957 9171 13991
rect 10149 13957 10183 13991
rect 14749 13957 14783 13991
rect 19809 13957 19843 13991
rect 2605 13889 2639 13923
rect 3065 13889 3099 13923
rect 9689 13889 9723 13923
rect 10793 13889 10827 13923
rect 11713 13889 11747 13923
rect 12449 13889 12483 13923
rect 17417 13889 17451 13923
rect 18429 13889 18463 13923
rect 20637 13889 20671 13923
rect 1409 13821 1443 13855
rect 2421 13821 2455 13855
rect 4721 13821 4755 13855
rect 4988 13821 5022 13855
rect 6653 13821 6687 13855
rect 7113 13821 7147 13855
rect 7369 13821 7403 13855
rect 10609 13821 10643 13855
rect 11621 13821 11655 13855
rect 13277 13821 13311 13855
rect 13369 13821 13403 13855
rect 13636 13821 13670 13855
rect 15209 13821 15243 13855
rect 15476 13821 15510 13855
rect 20545 13821 20579 13855
rect 21097 13821 21131 13855
rect 3332 13753 3366 13787
rect 9505 13753 9539 13787
rect 10517 13753 10551 13787
rect 11529 13753 11563 13787
rect 17325 13753 17359 13787
rect 18674 13753 18708 13787
rect 1961 13685 1995 13719
rect 2329 13685 2363 13719
rect 9597 13685 9631 13719
rect 17233 13685 17267 13719
rect 20453 13685 20487 13719
rect 21281 13685 21315 13719
rect 4353 13481 4387 13515
rect 5181 13481 5215 13515
rect 5549 13481 5583 13515
rect 6377 13481 6411 13515
rect 7389 13481 7423 13515
rect 7757 13481 7791 13515
rect 8401 13481 8435 13515
rect 8861 13481 8895 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 11069 13481 11103 13515
rect 12173 13481 12207 13515
rect 12541 13481 12575 13515
rect 15301 13481 15335 13515
rect 16313 13481 16347 13515
rect 18245 13481 18279 13515
rect 18797 13481 18831 13515
rect 19809 13481 19843 13515
rect 5641 13413 5675 13447
rect 6285 13413 6319 13447
rect 6745 13413 6779 13447
rect 8769 13413 8803 13447
rect 11437 13413 11471 13447
rect 11529 13413 11563 13447
rect 13636 13413 13670 13447
rect 18153 13413 18187 13447
rect 19165 13413 19199 13447
rect 20269 13413 20303 13447
rect 1593 13345 1627 13379
rect 2329 13345 2363 13379
rect 2596 13345 2630 13379
rect 4721 13345 4755 13379
rect 10057 13345 10091 13379
rect 12633 13345 12667 13379
rect 15669 13345 15703 13379
rect 16681 13345 16715 13379
rect 20177 13345 20211 13379
rect 20913 13345 20947 13379
rect 1777 13277 1811 13311
rect 4813 13277 4847 13311
rect 4997 13277 5031 13311
rect 5733 13277 5767 13311
rect 6837 13277 6871 13311
rect 7021 13277 7055 13311
rect 7849 13277 7883 13311
rect 7941 13277 7975 13311
rect 8953 13277 8987 13311
rect 10333 13277 10367 13311
rect 11713 13277 11747 13311
rect 12725 13277 12759 13311
rect 13369 13277 13403 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 16773 13277 16807 13311
rect 16957 13277 16991 13311
rect 18429 13277 18463 13311
rect 19257 13277 19291 13311
rect 19349 13277 19383 13311
rect 20453 13277 20487 13311
rect 21097 13277 21131 13311
rect 3709 13209 3743 13243
rect 14749 13209 14783 13243
rect 17785 13209 17819 13243
rect 2973 12937 3007 12971
rect 4169 12937 4203 12971
rect 5181 12937 5215 12971
rect 8217 12937 8251 12971
rect 10149 12937 10183 12971
rect 11161 12937 11195 12971
rect 13737 12937 13771 12971
rect 15301 12937 15335 12971
rect 17693 12937 17727 12971
rect 19717 12937 19751 12971
rect 4997 12869 5031 12903
rect 13461 12869 13495 12903
rect 18429 12869 18463 12903
rect 3433 12801 3467 12835
rect 4813 12801 4847 12835
rect 1593 12733 1627 12767
rect 3249 12733 3283 12767
rect 5733 12801 5767 12835
rect 6193 12801 6227 12835
rect 10701 12801 10735 12835
rect 11713 12801 11747 12835
rect 13001 12801 13035 12835
rect 14197 12801 14231 12835
rect 14381 12801 14415 12835
rect 15761 12801 15795 12835
rect 15945 12801 15979 12835
rect 16313 12801 16347 12835
rect 19073 12801 19107 12835
rect 20361 12801 20395 12835
rect 5641 12733 5675 12767
rect 6837 12733 6871 12767
rect 8493 12733 8527 12767
rect 13645 12733 13679 12767
rect 14105 12733 14139 12767
rect 20177 12733 20211 12767
rect 20729 12733 20763 12767
rect 1860 12665 1894 12699
rect 4537 12665 4571 12699
rect 4997 12665 5031 12699
rect 5549 12665 5583 12699
rect 7104 12665 7138 12699
rect 8760 12665 8794 12699
rect 11529 12665 11563 12699
rect 12817 12665 12851 12699
rect 14749 12665 14783 12699
rect 16580 12665 16614 12699
rect 18797 12665 18831 12699
rect 19625 12665 19659 12699
rect 20085 12665 20119 12699
rect 21005 12665 21039 12699
rect 4629 12597 4663 12631
rect 9873 12597 9907 12631
rect 10517 12597 10551 12631
rect 10609 12597 10643 12631
rect 11621 12597 11655 12631
rect 12449 12597 12483 12631
rect 12909 12597 12943 12631
rect 15669 12597 15703 12631
rect 18889 12597 18923 12631
rect 3617 12393 3651 12427
rect 4077 12393 4111 12427
rect 5089 12393 5123 12427
rect 8217 12393 8251 12427
rect 13737 12393 13771 12427
rect 17509 12393 17543 12427
rect 19441 12393 19475 12427
rect 19533 12393 19567 12427
rect 2044 12325 2078 12359
rect 7104 12325 7138 12359
rect 11989 12325 12023 12359
rect 12326 12325 12360 12359
rect 14197 12325 14231 12359
rect 18306 12325 18340 12359
rect 19993 12325 20027 12359
rect 1777 12257 1811 12291
rect 3433 12257 3467 12291
rect 4445 12257 4479 12291
rect 4537 12257 4571 12291
rect 5457 12257 5491 12291
rect 6837 12257 6871 12291
rect 8953 12257 8987 12291
rect 10692 12257 10726 12291
rect 4629 12189 4663 12223
rect 5549 12189 5583 12223
rect 5641 12189 5675 12223
rect 9045 12189 9079 12223
rect 9229 12189 9263 12223
rect 10425 12189 10459 12223
rect 12081 12257 12115 12291
rect 14105 12257 14139 12291
rect 15669 12257 15703 12291
rect 16396 12257 16430 12291
rect 17785 12257 17819 12291
rect 19901 12257 19935 12291
rect 20913 12257 20947 12291
rect 14381 12189 14415 12223
rect 15393 12189 15427 12223
rect 16129 12189 16163 12223
rect 18061 12189 18095 12223
rect 20085 12189 20119 12223
rect 21097 12189 21131 12223
rect 3157 12121 3191 12155
rect 11805 12121 11839 12155
rect 11989 12121 12023 12155
rect 8585 12053 8619 12087
rect 13461 12053 13495 12087
rect 15393 12053 15427 12087
rect 15485 12053 15519 12087
rect 1409 11849 1443 11883
rect 6837 11849 6871 11883
rect 16957 11849 16991 11883
rect 21281 11849 21315 11883
rect 3801 11781 3835 11815
rect 5273 11781 5307 11815
rect 9229 11781 9263 11815
rect 10701 11781 10735 11815
rect 13829 11781 13863 11815
rect 19073 11781 19107 11815
rect 2053 11713 2087 11747
rect 4905 11713 4939 11747
rect 5825 11713 5859 11747
rect 7481 11713 7515 11747
rect 7849 11713 7883 11747
rect 10149 11713 10183 11747
rect 11253 11713 11287 11747
rect 12081 11713 12115 11747
rect 12449 11713 12483 11747
rect 14289 11713 14323 11747
rect 16497 11713 16531 11747
rect 17417 11713 17451 11747
rect 17601 11713 17635 11747
rect 18613 11713 18647 11747
rect 19625 11713 19659 11747
rect 20545 11713 20579 11747
rect 20637 11713 20671 11747
rect 2421 11645 2455 11679
rect 4721 11645 4755 11679
rect 5733 11645 5767 11679
rect 11069 11645 11103 11679
rect 11897 11645 11931 11679
rect 11989 11645 12023 11679
rect 12716 11645 12750 11679
rect 14556 11645 14590 11679
rect 16313 11645 16347 11679
rect 16405 11645 16439 11679
rect 19441 11645 19475 11679
rect 19533 11645 19567 11679
rect 21097 11645 21131 11679
rect 2688 11577 2722 11611
rect 5641 11577 5675 11611
rect 8116 11577 8150 11611
rect 9965 11577 9999 11611
rect 17325 11577 17359 11611
rect 18521 11577 18555 11611
rect 18889 11577 18923 11611
rect 1777 11509 1811 11543
rect 1869 11509 1903 11543
rect 4261 11509 4295 11543
rect 4629 11509 4663 11543
rect 6285 11509 6319 11543
rect 7205 11509 7239 11543
rect 7297 11509 7331 11543
rect 9505 11509 9539 11543
rect 9873 11509 9907 11543
rect 11161 11509 11195 11543
rect 11529 11509 11563 11543
rect 15669 11509 15703 11543
rect 15945 11509 15979 11543
rect 18061 11509 18095 11543
rect 18429 11509 18463 11543
rect 20085 11509 20119 11543
rect 20453 11509 20487 11543
rect 1961 11305 1995 11339
rect 2329 11305 2363 11339
rect 2973 11305 3007 11339
rect 4077 11305 4111 11339
rect 4445 11305 4479 11339
rect 5825 11305 5859 11339
rect 6837 11305 6871 11339
rect 7297 11305 7331 11339
rect 7665 11305 7699 11339
rect 12541 11305 12575 11339
rect 14565 11305 14599 11339
rect 14657 11305 14691 11339
rect 18981 11305 19015 11339
rect 19717 11305 19751 11339
rect 20453 11305 20487 11339
rect 2421 11237 2455 11271
rect 6285 11237 6319 11271
rect 8953 11237 8987 11271
rect 9413 11237 9447 11271
rect 1409 11169 1443 11203
rect 3341 11169 3375 11203
rect 6193 11169 6227 11203
rect 7205 11169 7239 11203
rect 7665 11169 7699 11203
rect 8033 11169 8067 11203
rect 9045 11169 9079 11203
rect 2513 11101 2547 11135
rect 3433 11101 3467 11135
rect 3617 11101 3651 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 6377 11101 6411 11135
rect 7481 11101 7515 11135
rect 9229 11101 9263 11135
rect 1593 11033 1627 11067
rect 7849 11033 7883 11067
rect 15669 11237 15703 11271
rect 17846 11237 17880 11271
rect 21189 11237 21223 11271
rect 10333 11169 10367 11203
rect 13001 11169 13035 11203
rect 13268 11169 13302 11203
rect 14565 11169 14599 11203
rect 15761 11169 15795 11203
rect 16681 11169 16715 11203
rect 19625 11169 19659 11203
rect 20269 11169 20303 11203
rect 20913 11169 20947 11203
rect 12633 11101 12667 11135
rect 12725 11101 12759 11135
rect 15853 11101 15887 11135
rect 16773 11101 16807 11135
rect 16865 11101 16899 11135
rect 17601 11101 17635 11135
rect 19809 11101 19843 11135
rect 11621 11033 11655 11067
rect 14381 11033 14415 11067
rect 15301 11033 15335 11067
rect 8585 10965 8619 10999
rect 9413 10965 9447 10999
rect 12173 10965 12207 10999
rect 16313 10965 16347 10999
rect 19257 10965 19291 10999
rect 1961 10761 1995 10795
rect 5549 10761 5583 10795
rect 6837 10761 6871 10795
rect 9689 10761 9723 10795
rect 16773 10761 16807 10795
rect 21189 10761 21223 10795
rect 18061 10693 18095 10727
rect 2513 10625 2547 10659
rect 3617 10625 3651 10659
rect 7389 10625 7423 10659
rect 8217 10625 8251 10659
rect 10333 10625 10367 10659
rect 11437 10625 11471 10659
rect 11713 10625 11747 10659
rect 12817 10625 12851 10659
rect 15025 10625 15059 10659
rect 16221 10625 16255 10659
rect 17417 10625 17451 10659
rect 18613 10625 18647 10659
rect 19349 10625 19383 10659
rect 3341 10557 3375 10591
rect 3433 10557 3467 10591
rect 4169 10557 4203 10591
rect 8033 10557 8067 10591
rect 8484 10557 8518 10591
rect 11345 10557 11379 10591
rect 13084 10557 13118 10591
rect 14933 10557 14967 10591
rect 16037 10557 16071 10591
rect 18429 10557 18463 10591
rect 18521 10557 18555 10591
rect 19616 10557 19650 10591
rect 21005 10557 21039 10591
rect 4436 10489 4470 10523
rect 7297 10489 7331 10523
rect 10057 10489 10091 10523
rect 10149 10489 10183 10523
rect 14841 10489 14875 10523
rect 17233 10489 17267 10523
rect 2329 10421 2363 10455
rect 2421 10421 2455 10455
rect 2973 10421 3007 10455
rect 6285 10421 6319 10455
rect 7205 10421 7239 10455
rect 7849 10421 7883 10455
rect 9597 10421 9631 10455
rect 10885 10421 10919 10455
rect 11253 10421 11287 10455
rect 14197 10421 14231 10455
rect 14473 10421 14507 10455
rect 15669 10421 15703 10455
rect 16129 10421 16163 10455
rect 16865 10421 16899 10455
rect 17325 10421 17359 10455
rect 20729 10421 20763 10455
rect 2237 10217 2271 10251
rect 6285 10217 6319 10251
rect 7941 10217 7975 10251
rect 8217 10217 8251 10251
rect 8585 10217 8619 10251
rect 8677 10217 8711 10251
rect 9781 10217 9815 10251
rect 10241 10217 10275 10251
rect 11989 10217 12023 10251
rect 13277 10217 13311 10251
rect 13645 10217 13679 10251
rect 17417 10217 17451 10251
rect 20269 10217 20303 10251
rect 5172 10149 5206 10183
rect 10876 10149 10910 10183
rect 12725 10149 12759 10183
rect 19156 10149 19190 10183
rect 2605 10081 2639 10115
rect 3249 10081 3283 10115
rect 4905 10081 4939 10115
rect 6817 10081 6851 10115
rect 10149 10081 10183 10115
rect 10609 10081 10643 10115
rect 12633 10081 12667 10115
rect 13737 10081 13771 10115
rect 15301 10081 15335 10115
rect 15568 10081 15602 10115
rect 17325 10081 17359 10115
rect 18889 10081 18923 10115
rect 2697 10013 2731 10047
rect 2881 10013 2915 10047
rect 6561 10013 6595 10047
rect 8769 10013 8803 10047
rect 10333 10013 10367 10047
rect 12817 10013 12851 10047
rect 13829 10013 13863 10047
rect 17601 10013 17635 10047
rect 12265 9877 12299 9911
rect 16681 9877 16715 9911
rect 16957 9877 16991 9911
rect 2053 9673 2087 9707
rect 5733 9605 5767 9639
rect 6837 9605 6871 9639
rect 7849 9605 7883 9639
rect 8953 9605 8987 9639
rect 12449 9605 12483 9639
rect 19441 9605 19475 9639
rect 2605 9537 2639 9571
rect 6377 9537 6411 9571
rect 7389 9537 7423 9571
rect 8401 9537 8435 9571
rect 9505 9537 9539 9571
rect 10517 9537 10551 9571
rect 11529 9537 11563 9571
rect 13093 9537 13127 9571
rect 14105 9537 14139 9571
rect 14841 9537 14875 9571
rect 17049 9537 17083 9571
rect 17509 9537 17543 9571
rect 21005 9537 21039 9571
rect 3249 9469 3283 9503
rect 6101 9469 6135 9503
rect 7205 9469 7239 9503
rect 9413 9469 9447 9503
rect 10333 9469 10367 9503
rect 11437 9469 11471 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 13921 9469 13955 9503
rect 14657 9469 14691 9503
rect 15108 9469 15142 9503
rect 16865 9469 16899 9503
rect 18061 9469 18095 9503
rect 20821 9469 20855 9503
rect 3494 9401 3528 9435
rect 11345 9401 11379 9435
rect 18328 9401 18362 9435
rect 2421 9333 2455 9367
rect 2513 9333 2547 9367
rect 4629 9333 4663 9367
rect 6193 9333 6227 9367
rect 7297 9333 7331 9367
rect 8217 9333 8251 9367
rect 8309 9333 8343 9367
rect 9321 9333 9355 9367
rect 9965 9333 9999 9367
rect 10425 9333 10459 9367
rect 10977 9333 11011 9367
rect 13461 9333 13495 9367
rect 13829 9333 13863 9367
rect 14473 9333 14507 9367
rect 16221 9333 16255 9367
rect 16497 9333 16531 9367
rect 16957 9333 16991 9367
rect 20453 9333 20487 9367
rect 20913 9333 20947 9367
rect 3249 9129 3283 9163
rect 4077 9129 4111 9163
rect 4537 9129 4571 9163
rect 5089 9129 5123 9163
rect 5457 9129 5491 9163
rect 6101 9129 6135 9163
rect 6469 9129 6503 9163
rect 8953 9129 8987 9163
rect 9045 9129 9079 9163
rect 9689 9129 9723 9163
rect 14657 9129 14691 9163
rect 15761 9129 15795 9163
rect 19533 9129 19567 9163
rect 20913 9129 20947 9163
rect 7573 9061 7607 9095
rect 9413 9061 9447 9095
rect 12624 9061 12658 9095
rect 1869 8993 1903 9027
rect 2136 8993 2170 9027
rect 4445 8993 4479 9027
rect 7481 8993 7515 9027
rect 10129 8993 10163 9027
rect 14565 8993 14599 9027
rect 15669 8993 15703 9027
rect 16681 8993 16715 9027
rect 17684 8993 17718 9027
rect 18889 8993 18923 9027
rect 19441 8993 19475 9027
rect 4629 8925 4663 8959
rect 5549 8925 5583 8959
rect 5641 8925 5675 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 7665 8925 7699 8959
rect 8125 8925 8159 8959
rect 9137 8925 9171 8959
rect 9873 8925 9907 8959
rect 12357 8925 12391 8959
rect 14841 8925 14875 8959
rect 15853 8925 15887 8959
rect 16773 8925 16807 8959
rect 16865 8925 16899 8959
rect 17417 8925 17451 8959
rect 7113 8857 7147 8891
rect 8585 8857 8619 8891
rect 11253 8857 11287 8891
rect 13737 8857 13771 8891
rect 15301 8857 15335 8891
rect 18797 8857 18831 8891
rect 19625 8925 19659 8959
rect 14197 8789 14231 8823
rect 16313 8789 16347 8823
rect 18889 8789 18923 8823
rect 19073 8789 19107 8823
rect 3249 8585 3283 8619
rect 5273 8585 5307 8619
rect 11529 8585 11563 8619
rect 12449 8585 12483 8619
rect 4997 8517 5031 8551
rect 6285 8517 6319 8551
rect 8217 8517 8251 8551
rect 9873 8517 9907 8551
rect 9965 8517 9999 8551
rect 13645 8517 13679 8551
rect 18245 8517 18279 8551
rect 18889 8517 18923 8551
rect 5825 8449 5859 8483
rect 6837 8449 6871 8483
rect 8493 8449 8527 8483
rect 1869 8381 1903 8415
rect 3617 8381 3651 8415
rect 6469 8381 6503 8415
rect 7104 8381 7138 8415
rect 8760 8381 8794 8415
rect 10149 8449 10183 8483
rect 13001 8449 13035 8483
rect 14197 8449 14231 8483
rect 15761 8449 15795 8483
rect 15945 8449 15979 8483
rect 16865 8449 16899 8483
rect 19349 8449 19383 8483
rect 19533 8449 19567 8483
rect 20637 8449 20671 8483
rect 15209 8381 15243 8415
rect 15669 8381 15703 8415
rect 18061 8381 18095 8415
rect 2136 8313 2170 8347
rect 3884 8313 3918 8347
rect 5733 8313 5767 8347
rect 9965 8313 9999 8347
rect 10394 8313 10428 8347
rect 12817 8313 12851 8347
rect 13277 8313 13311 8347
rect 14013 8313 14047 8347
rect 16773 8313 16807 8347
rect 19257 8313 19291 8347
rect 5641 8245 5675 8279
rect 12909 8245 12943 8279
rect 14105 8245 14139 8279
rect 15025 8245 15059 8279
rect 15301 8245 15335 8279
rect 16313 8245 16347 8279
rect 16681 8245 16715 8279
rect 20085 8245 20119 8279
rect 20453 8245 20487 8279
rect 20545 8245 20579 8279
rect 2145 8041 2179 8075
rect 4997 8041 5031 8075
rect 6285 8041 6319 8075
rect 7757 8041 7791 8075
rect 8309 8041 8343 8075
rect 8953 8041 8987 8075
rect 9965 8041 9999 8075
rect 11345 8041 11379 8075
rect 11437 8041 11471 8075
rect 16957 8041 16991 8075
rect 17325 8041 17359 8075
rect 17417 8041 17451 8075
rect 18429 8041 18463 8075
rect 2605 7973 2639 8007
rect 6653 7973 6687 8007
rect 10425 7973 10459 8007
rect 19318 7973 19352 8007
rect 2513 7905 2547 7939
rect 3157 7905 3191 7939
rect 5365 7905 5399 7939
rect 5457 7905 5491 7939
rect 6745 7905 6779 7939
rect 7665 7905 7699 7939
rect 8493 7905 8527 7939
rect 10333 7905 10367 7939
rect 11989 7905 12023 7939
rect 12633 7905 12667 7939
rect 12992 7905 13026 7939
rect 14381 7905 14415 7939
rect 15301 7905 15335 7939
rect 15568 7905 15602 7939
rect 18337 7905 18371 7939
rect 2697 7837 2731 7871
rect 5549 7837 5583 7871
rect 6837 7837 6871 7871
rect 7849 7837 7883 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 10609 7837 10643 7871
rect 11621 7837 11655 7871
rect 12725 7837 12759 7871
rect 17509 7837 17543 7871
rect 18521 7837 18555 7871
rect 19073 7837 19107 7871
rect 7297 7769 7331 7803
rect 8585 7701 8619 7735
rect 10977 7701 11011 7735
rect 12449 7701 12483 7735
rect 14105 7701 14139 7735
rect 14565 7701 14599 7735
rect 16681 7701 16715 7735
rect 17969 7701 18003 7735
rect 20453 7701 20487 7735
rect 2329 7497 2363 7531
rect 6193 7497 6227 7531
rect 7481 7497 7515 7531
rect 20085 7497 20119 7531
rect 20361 7497 20395 7531
rect 10517 7429 10551 7463
rect 15577 7429 15611 7463
rect 2881 7361 2915 7395
rect 3893 7361 3927 7395
rect 4813 7361 4847 7395
rect 8125 7361 8159 7395
rect 9321 7361 9355 7395
rect 10241 7361 10275 7395
rect 1593 7293 1627 7327
rect 3709 7293 3743 7327
rect 10057 7293 10091 7327
rect 1869 7225 1903 7259
rect 5058 7225 5092 7259
rect 7941 7225 7975 7259
rect 8585 7225 8619 7259
rect 9045 7225 9079 7259
rect 10149 7225 10183 7259
rect 12173 7361 12207 7395
rect 13001 7361 13035 7395
rect 16405 7361 16439 7395
rect 16497 7361 16531 7395
rect 17601 7361 17635 7395
rect 20913 7361 20947 7395
rect 10701 7293 10735 7327
rect 10968 7225 11002 7259
rect 13461 7293 13495 7327
rect 13728 7293 13762 7327
rect 15393 7293 15427 7327
rect 17325 7293 17359 7327
rect 18061 7293 18095 7327
rect 18705 7293 18739 7327
rect 20821 7293 20855 7327
rect 16313 7225 16347 7259
rect 18972 7225 19006 7259
rect 20729 7225 20763 7259
rect 2697 7157 2731 7191
rect 2789 7157 2823 7191
rect 3341 7157 3375 7191
rect 3801 7157 3835 7191
rect 4353 7157 4387 7191
rect 7849 7157 7883 7191
rect 8677 7157 8711 7191
rect 9137 7157 9171 7191
rect 9689 7157 9723 7191
rect 10517 7157 10551 7191
rect 12081 7157 12115 7191
rect 12173 7157 12207 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 12909 7157 12943 7191
rect 14841 7157 14875 7191
rect 15945 7157 15979 7191
rect 16957 7157 16991 7191
rect 17417 7157 17451 7191
rect 18245 7157 18279 7191
rect 3341 6953 3375 6987
rect 6193 6953 6227 6987
rect 7481 6953 7515 6987
rect 7849 6953 7883 6987
rect 8861 6953 8895 6987
rect 10057 6953 10091 6987
rect 14565 6953 14599 6987
rect 16589 6953 16623 6987
rect 16957 6953 16991 6987
rect 4445 6885 4479 6919
rect 5641 6885 5675 6919
rect 6101 6885 6135 6919
rect 12725 6885 12759 6919
rect 14657 6885 14691 6919
rect 16497 6885 16531 6919
rect 1961 6817 1995 6851
rect 2228 6817 2262 6851
rect 10149 6817 10183 6851
rect 10968 6817 11002 6851
rect 13645 6817 13679 6851
rect 15602 6817 15636 6851
rect 4537 6749 4571 6783
rect 4629 6749 4663 6783
rect 6285 6749 6319 6783
rect 7941 6749 7975 6783
rect 8125 6749 8159 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 10241 6749 10275 6783
rect 10701 6749 10735 6783
rect 12817 6749 12851 6783
rect 12909 6749 12943 6783
rect 14841 6749 14875 6783
rect 16681 6749 16715 6783
rect 17509 6885 17543 6919
rect 17601 6817 17635 6851
rect 18521 6817 18555 6851
rect 18788 6817 18822 6851
rect 20177 6817 20211 6851
rect 17693 6749 17727 6783
rect 20913 6749 20947 6783
rect 8493 6681 8527 6715
rect 14197 6681 14231 6715
rect 16129 6681 16163 6715
rect 16957 6681 16991 6715
rect 17141 6681 17175 6715
rect 19901 6681 19935 6715
rect 4077 6613 4111 6647
rect 5733 6613 5767 6647
rect 9689 6613 9723 6647
rect 12081 6613 12115 6647
rect 12357 6613 12391 6647
rect 13829 6613 13863 6647
rect 15761 6613 15795 6647
rect 20361 6613 20395 6647
rect 2789 6409 2823 6443
rect 3065 6409 3099 6443
rect 9597 6409 9631 6443
rect 11069 6409 11103 6443
rect 16037 6409 16071 6443
rect 19073 6409 19107 6443
rect 20085 6409 20119 6443
rect 5457 6341 5491 6375
rect 9321 6341 9355 6375
rect 14289 6341 14323 6375
rect 18061 6341 18095 6375
rect 3525 6273 3559 6307
rect 3617 6273 3651 6307
rect 6101 6273 6135 6307
rect 7389 6273 7423 6307
rect 10149 6273 10183 6307
rect 11621 6273 11655 6307
rect 15669 6273 15703 6307
rect 16589 6273 16623 6307
rect 18705 6273 18739 6307
rect 19533 6273 19567 6307
rect 19717 6273 19751 6307
rect 20729 6273 20763 6307
rect 1409 6205 1443 6239
rect 4077 6205 4111 6239
rect 6009 6205 6043 6239
rect 7205 6205 7239 6239
rect 7941 6205 7975 6239
rect 11437 6205 11471 6239
rect 11529 6205 11563 6239
rect 12909 6205 12943 6239
rect 13176 6205 13210 6239
rect 15485 6205 15519 6239
rect 16405 6205 16439 6239
rect 17417 6205 17451 6239
rect 20453 6205 20487 6239
rect 20545 6205 20579 6239
rect 21097 6205 21131 6239
rect 1676 6137 1710 6171
rect 4322 6137 4356 6171
rect 7297 6137 7331 6171
rect 8208 6137 8242 6171
rect 18429 6137 18463 6171
rect 3433 6069 3467 6103
rect 5549 6069 5583 6103
rect 5917 6069 5951 6103
rect 6377 6069 6411 6103
rect 6837 6069 6871 6103
rect 9965 6069 9999 6103
rect 10057 6069 10091 6103
rect 10609 6069 10643 6103
rect 15025 6069 15059 6103
rect 15393 6069 15427 6103
rect 16497 6069 16531 6103
rect 17601 6069 17635 6103
rect 18521 6069 18555 6103
rect 19441 6069 19475 6103
rect 21281 6069 21315 6103
rect 3249 5865 3283 5899
rect 4077 5865 4111 5899
rect 4445 5865 4479 5899
rect 5641 5865 5675 5899
rect 6469 5865 6503 5899
rect 6561 5865 6595 5899
rect 7665 5865 7699 5899
rect 8585 5865 8619 5899
rect 17049 5865 17083 5899
rect 19901 5865 19935 5899
rect 4537 5797 4571 5831
rect 8953 5797 8987 5831
rect 10232 5797 10266 5831
rect 14197 5797 14231 5831
rect 15660 5797 15694 5831
rect 18788 5797 18822 5831
rect 1869 5729 1903 5763
rect 2136 5729 2170 5763
rect 5549 5729 5583 5763
rect 7757 5729 7791 5763
rect 9045 5729 9079 5763
rect 9965 5729 9999 5763
rect 12081 5729 12115 5763
rect 12173 5729 12207 5763
rect 13093 5729 13127 5763
rect 14105 5729 14139 5763
rect 16865 5729 16899 5763
rect 17417 5729 17451 5763
rect 18061 5729 18095 5763
rect 18521 5729 18555 5763
rect 20269 5729 20303 5763
rect 20913 5729 20947 5763
rect 4629 5661 4663 5695
rect 5825 5661 5859 5695
rect 6745 5661 6779 5695
rect 7849 5661 7883 5695
rect 9137 5661 9171 5695
rect 12357 5661 12391 5695
rect 13185 5661 13219 5695
rect 13369 5661 13403 5695
rect 14289 5661 14323 5695
rect 14749 5661 14783 5695
rect 15393 5661 15427 5695
rect 11713 5593 11747 5627
rect 12725 5593 12759 5627
rect 17509 5661 17543 5695
rect 17601 5661 17635 5695
rect 20453 5593 20487 5627
rect 5181 5525 5215 5559
rect 6101 5525 6135 5559
rect 7205 5525 7239 5559
rect 7297 5525 7331 5559
rect 11345 5525 11379 5559
rect 13737 5525 13771 5559
rect 16773 5525 16807 5559
rect 16865 5525 16899 5559
rect 21097 5525 21131 5559
rect 1961 5321 1995 5355
rect 8217 5321 8251 5355
rect 11989 5321 12023 5355
rect 17049 5321 17083 5355
rect 19165 5321 19199 5355
rect 20177 5321 20211 5355
rect 8493 5253 8527 5287
rect 14105 5253 14139 5287
rect 14289 5253 14323 5287
rect 17601 5253 17635 5287
rect 2513 5185 2547 5219
rect 3157 5185 3191 5219
rect 6285 5185 6319 5219
rect 9137 5185 9171 5219
rect 10241 5185 10275 5219
rect 11161 5185 11195 5219
rect 11345 5185 11379 5219
rect 12173 5185 12207 5219
rect 13829 5185 13863 5219
rect 3424 5117 3458 5151
rect 6101 5117 6135 5151
rect 6193 5117 6227 5151
rect 6837 5117 6871 5151
rect 8861 5117 8895 5151
rect 11805 5117 11839 5151
rect 2329 5049 2363 5083
rect 7104 5049 7138 5083
rect 10057 5049 10091 5083
rect 12725 5117 12759 5151
rect 13737 5117 13771 5151
rect 14933 5185 14967 5219
rect 18797 5185 18831 5219
rect 19717 5185 19751 5219
rect 20821 5185 20855 5219
rect 21005 5185 21039 5219
rect 14657 5117 14691 5151
rect 15669 5117 15703 5151
rect 15936 5117 15970 5151
rect 17417 5117 17451 5151
rect 18521 5117 18555 5151
rect 20729 5117 20763 5151
rect 13645 5049 13679 5083
rect 14105 5049 14139 5083
rect 18613 5049 18647 5083
rect 19533 5049 19567 5083
rect 2421 4981 2455 5015
rect 4537 4981 4571 5015
rect 5733 4981 5767 5015
rect 8953 4981 8987 5015
rect 9689 4981 9723 5015
rect 10149 4981 10183 5015
rect 10701 4981 10735 5015
rect 11069 4981 11103 5015
rect 12173 4981 12207 5015
rect 12909 4981 12943 5015
rect 13277 4981 13311 5015
rect 14749 4981 14783 5015
rect 18153 4981 18187 5015
rect 19625 4981 19659 5015
rect 20361 4981 20395 5015
rect 2145 4777 2179 4811
rect 4353 4777 4387 4811
rect 4813 4777 4847 4811
rect 7573 4777 7607 4811
rect 7665 4777 7699 4811
rect 9689 4777 9723 4811
rect 11161 4777 11195 4811
rect 17417 4777 17451 4811
rect 19441 4777 19475 4811
rect 2605 4709 2639 4743
rect 4721 4709 4755 4743
rect 10057 4709 10091 4743
rect 14565 4709 14599 4743
rect 16120 4709 16154 4743
rect 2513 4641 2547 4675
rect 3157 4641 3191 4675
rect 5805 4641 5839 4675
rect 8585 4641 8619 4675
rect 10149 4641 10183 4675
rect 11069 4641 11103 4675
rect 12081 4641 12115 4675
rect 12900 4641 12934 4675
rect 14289 4641 14323 4675
rect 15301 4641 15335 4675
rect 15853 4641 15887 4675
rect 19901 4709 19935 4743
rect 17776 4641 17810 4675
rect 19809 4641 19843 4675
rect 20913 4641 20947 4675
rect 2697 4573 2731 4607
rect 4905 4573 4939 4607
rect 5549 4573 5583 4607
rect 7757 4573 7791 4607
rect 8677 4573 8711 4607
rect 8861 4573 8895 4607
rect 10241 4573 10275 4607
rect 11253 4573 11287 4607
rect 12633 4573 12667 4607
rect 17417 4573 17451 4607
rect 17509 4573 17543 4607
rect 20085 4573 20119 4607
rect 6929 4505 6963 4539
rect 17233 4505 17267 4539
rect 18889 4505 18923 4539
rect 7205 4437 7239 4471
rect 8217 4437 8251 4471
rect 10701 4437 10735 4471
rect 12265 4437 12299 4471
rect 14013 4437 14047 4471
rect 15485 4437 15519 4471
rect 21097 4437 21131 4471
rect 2421 4233 2455 4267
rect 9505 4233 9539 4267
rect 15761 4233 15795 4267
rect 9229 4165 9263 4199
rect 10333 4165 10367 4199
rect 2973 4097 3007 4131
rect 3893 4097 3927 4131
rect 4077 4097 4111 4131
rect 7297 4097 7331 4131
rect 7389 4097 7423 4131
rect 10057 4097 10091 4131
rect 2789 4029 2823 4063
rect 4997 4029 5031 4063
rect 5264 4029 5298 4063
rect 7849 4029 7883 4063
rect 9965 4029 9999 4063
rect 3801 3961 3835 3995
rect 8116 3961 8150 3995
rect 11161 4097 11195 4131
rect 11805 4097 11839 4131
rect 13277 4097 13311 4131
rect 14197 4097 14231 4131
rect 14289 4097 14323 4131
rect 15117 4097 15151 4131
rect 16313 4097 16347 4131
rect 17509 4097 17543 4131
rect 18981 4097 19015 4131
rect 20085 4097 20119 4131
rect 20913 4097 20947 4131
rect 21005 4097 21039 4131
rect 11621 4029 11655 4063
rect 13093 4029 13127 4063
rect 17785 4029 17819 4063
rect 19809 4029 19843 4063
rect 14933 3961 14967 3995
rect 15025 3961 15059 3995
rect 15577 3961 15611 3995
rect 16129 3961 16163 3995
rect 18797 3961 18831 3995
rect 2881 3893 2915 3927
rect 3433 3893 3467 3927
rect 6377 3893 6411 3927
rect 6837 3893 6871 3927
rect 7205 3893 7239 3927
rect 9873 3893 9907 3927
rect 10333 3893 10367 3927
rect 10517 3893 10551 3927
rect 10885 3893 10919 3927
rect 10977 3893 11011 3927
rect 12725 3893 12759 3927
rect 13185 3893 13219 3927
rect 13737 3893 13771 3927
rect 14105 3893 14139 3927
rect 14565 3893 14599 3927
rect 16221 3893 16255 3927
rect 16957 3893 16991 3927
rect 17325 3893 17359 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 18429 3893 18463 3927
rect 18889 3893 18923 3927
rect 19441 3893 19475 3927
rect 19901 3893 19935 3927
rect 20453 3893 20487 3927
rect 20821 3893 20855 3927
rect 5181 3689 5215 3723
rect 11437 3689 11471 3723
rect 11897 3689 11931 3723
rect 14197 3689 14231 3723
rect 15301 3689 15335 3723
rect 15669 3689 15703 3723
rect 17049 3689 17083 3723
rect 18521 3689 18555 3723
rect 18889 3689 18923 3723
rect 19533 3689 19567 3723
rect 2329 3621 2363 3655
rect 2881 3621 2915 3655
rect 16957 3621 16991 3655
rect 17877 3621 17911 3655
rect 19993 3621 20027 3655
rect 21189 3621 21223 3655
rect 2421 3553 2455 3587
rect 2605 3485 2639 3519
rect 3341 3553 3375 3587
rect 5825 3553 5859 3587
rect 6081 3553 6115 3587
rect 8197 3553 8231 3587
rect 10048 3553 10082 3587
rect 11805 3553 11839 3587
rect 13084 3553 13118 3587
rect 14473 3553 14507 3587
rect 17601 3553 17635 3587
rect 19901 3553 19935 3587
rect 20913 3553 20947 3587
rect 3433 3485 3467 3519
rect 3525 3485 3559 3519
rect 5273 3485 5307 3519
rect 5457 3485 5491 3519
rect 7941 3485 7975 3519
rect 9781 3485 9815 3519
rect 12081 3485 12115 3519
rect 12817 3485 12851 3519
rect 14657 3485 14691 3519
rect 15761 3485 15795 3519
rect 15945 3485 15979 3519
rect 17233 3485 17267 3519
rect 18981 3485 19015 3519
rect 19073 3485 19107 3519
rect 20177 3485 20211 3519
rect 1961 3417 1995 3451
rect 2881 3417 2915 3451
rect 9321 3417 9355 3451
rect 16589 3417 16623 3451
rect 2973 3349 3007 3383
rect 4813 3349 4847 3383
rect 7205 3349 7239 3383
rect 11161 3349 11195 3383
rect 2973 3145 3007 3179
rect 5641 3145 5675 3179
rect 7205 3145 7239 3179
rect 10057 3145 10091 3179
rect 11897 3145 11931 3179
rect 15301 3145 15335 3179
rect 16497 3145 16531 3179
rect 20453 3145 20487 3179
rect 14473 3077 14507 3111
rect 16313 3077 16347 3111
rect 18889 3077 18923 3111
rect 19441 3077 19475 3111
rect 3617 3009 3651 3043
rect 6193 3009 6227 3043
rect 7665 3009 7699 3043
rect 7757 3009 7791 3043
rect 8677 3009 8711 3043
rect 15117 3009 15151 3043
rect 15945 3009 15979 3043
rect 17049 3009 17083 3043
rect 18613 3009 18647 3043
rect 19901 3009 19935 3043
rect 19993 3009 20027 3043
rect 21097 3009 21131 3043
rect 3433 2941 3467 2975
rect 3985 2941 4019 2975
rect 10517 2941 10551 2975
rect 12817 2941 12851 2975
rect 14841 2941 14875 2975
rect 15669 2941 15703 2975
rect 16865 2941 16899 2975
rect 17969 2941 18003 2975
rect 19809 2941 19843 2975
rect 4252 2873 4286 2907
rect 6101 2873 6135 2907
rect 7573 2873 7607 2907
rect 8944 2873 8978 2907
rect 10784 2873 10818 2907
rect 13084 2873 13118 2907
rect 15761 2873 15795 2907
rect 18429 2873 18463 2907
rect 18521 2873 18555 2907
rect 20821 2873 20855 2907
rect 3341 2805 3375 2839
rect 5365 2805 5399 2839
rect 6009 2805 6043 2839
rect 14197 2805 14231 2839
rect 14933 2805 14967 2839
rect 16957 2805 16991 2839
rect 17877 2805 17911 2839
rect 18061 2805 18095 2839
rect 20913 2805 20947 2839
rect 4813 2601 4847 2635
rect 5825 2601 5859 2635
rect 6285 2601 6319 2635
rect 7389 2601 7423 2635
rect 7941 2601 7975 2635
rect 10885 2601 10919 2635
rect 11437 2601 11471 2635
rect 11897 2601 11931 2635
rect 13001 2601 13035 2635
rect 13645 2601 13679 2635
rect 14013 2601 14047 2635
rect 15485 2601 15519 2635
rect 16497 2601 16531 2635
rect 18337 2601 18371 2635
rect 18705 2601 18739 2635
rect 18797 2601 18831 2635
rect 19717 2601 19751 2635
rect 7297 2533 7331 2567
rect 10793 2533 10827 2567
rect 14933 2533 14967 2567
rect 15853 2533 15887 2567
rect 17785 2533 17819 2567
rect 19809 2533 19843 2567
rect 5181 2465 5215 2499
rect 6193 2465 6227 2499
rect 8309 2465 8343 2499
rect 9137 2465 9171 2499
rect 9873 2465 9907 2499
rect 11805 2465 11839 2499
rect 14105 2465 14139 2499
rect 14657 2465 14691 2499
rect 15945 2465 15979 2499
rect 16865 2465 16899 2499
rect 16957 2465 16991 2499
rect 17509 2465 17543 2499
rect 20545 2465 20579 2499
rect 5273 2397 5307 2431
rect 5457 2397 5491 2431
rect 6469 2397 6503 2431
rect 7481 2397 7515 2431
rect 8401 2397 8435 2431
rect 8585 2397 8619 2431
rect 11069 2397 11103 2431
rect 12081 2397 12115 2431
rect 13093 2397 13127 2431
rect 13185 2397 13219 2431
rect 14197 2397 14231 2431
rect 16037 2397 16071 2431
rect 17049 2397 17083 2431
rect 18889 2397 18923 2431
rect 19901 2397 19935 2431
rect 9321 2329 9355 2363
rect 12633 2329 12667 2363
rect 19349 2329 19383 2363
rect 6929 2261 6963 2295
rect 10057 2261 10091 2295
rect 10425 2261 10459 2295
rect 20729 2261 20763 2295
<< metal1 >>
rect 9858 20748 9864 20800
rect 9916 20788 9922 20800
rect 13538 20788 13544 20800
rect 9916 20760 13544 20788
rect 9916 20748 9922 20760
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 2501 20587 2559 20593
rect 2501 20553 2513 20587
rect 2547 20584 2559 20587
rect 2774 20584 2780 20596
rect 2547 20556 2780 20584
rect 2547 20553 2559 20556
rect 2501 20547 2559 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 3694 20544 3700 20596
rect 3752 20584 3758 20596
rect 5813 20587 5871 20593
rect 3752 20556 5764 20584
rect 3752 20544 3758 20556
rect 5736 20516 5764 20556
rect 5813 20553 5825 20587
rect 5859 20584 5871 20587
rect 15010 20584 15016 20596
rect 5859 20556 12020 20584
rect 14971 20556 15016 20584
rect 5859 20553 5871 20556
rect 5813 20547 5871 20553
rect 9950 20516 9956 20528
rect 5736 20488 9956 20516
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 10321 20519 10379 20525
rect 10321 20485 10333 20519
rect 10367 20485 10379 20519
rect 10321 20479 10379 20485
rect 6365 20451 6423 20457
rect 6365 20417 6377 20451
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 8021 20451 8079 20457
rect 8021 20417 8033 20451
rect 8067 20448 8079 20451
rect 8202 20448 8208 20460
rect 8067 20420 8208 20448
rect 8067 20417 8079 20420
rect 8021 20411 8079 20417
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20380 2375 20383
rect 3326 20380 3332 20392
rect 2363 20352 3332 20380
rect 2363 20349 2375 20352
rect 2317 20343 2375 20349
rect 3326 20340 3332 20352
rect 3384 20340 3390 20392
rect 3786 20340 3792 20392
rect 3844 20380 3850 20392
rect 4065 20383 4123 20389
rect 4065 20380 4077 20383
rect 3844 20352 4077 20380
rect 3844 20340 3850 20352
rect 4065 20349 4077 20352
rect 4111 20349 4123 20383
rect 4065 20343 4123 20349
rect 4332 20383 4390 20389
rect 4332 20349 4344 20383
rect 4378 20380 4390 20383
rect 6380 20380 6408 20411
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 9033 20451 9091 20457
rect 9033 20417 9045 20451
rect 9079 20448 9091 20451
rect 9306 20448 9312 20460
rect 9079 20420 9312 20448
rect 9079 20417 9091 20420
rect 9033 20411 9091 20417
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 7374 20380 7380 20392
rect 4378 20352 7380 20380
rect 4378 20349 4390 20352
rect 4332 20343 4390 20349
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 10336 20380 10364 20479
rect 10594 20476 10600 20528
rect 10652 20516 10658 20528
rect 11054 20516 11060 20528
rect 10652 20488 11060 20516
rect 10652 20476 10658 20488
rect 11054 20476 11060 20488
rect 11112 20516 11118 20528
rect 11112 20488 11928 20516
rect 11112 20476 11118 20488
rect 10410 20408 10416 20460
rect 10468 20448 10474 20460
rect 10781 20451 10839 20457
rect 10781 20448 10793 20451
rect 10468 20420 10793 20448
rect 10468 20408 10474 20420
rect 10781 20417 10793 20420
rect 10827 20417 10839 20451
rect 10962 20448 10968 20460
rect 10923 20420 10968 20448
rect 10781 20411 10839 20417
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 11900 20457 11928 20488
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20417 11943 20451
rect 11992 20448 12020 20556
rect 15010 20544 15016 20556
rect 15068 20544 15074 20596
rect 15930 20584 15936 20596
rect 15891 20556 15936 20584
rect 15930 20544 15936 20556
rect 15988 20544 15994 20596
rect 16669 20587 16727 20593
rect 16669 20553 16681 20587
rect 16715 20584 16727 20587
rect 16942 20584 16948 20596
rect 16715 20556 16948 20584
rect 16715 20553 16727 20556
rect 16669 20547 16727 20553
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 19521 20587 19579 20593
rect 19521 20553 19533 20587
rect 19567 20584 19579 20587
rect 20254 20584 20260 20596
rect 19567 20556 20260 20584
rect 19567 20553 19579 20556
rect 19521 20547 19579 20553
rect 20254 20544 20260 20556
rect 20312 20544 20318 20596
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 20717 20587 20775 20593
rect 20717 20584 20729 20587
rect 20680 20556 20729 20584
rect 20680 20544 20686 20556
rect 20717 20553 20729 20556
rect 20763 20553 20775 20587
rect 20717 20547 20775 20553
rect 12621 20519 12679 20525
rect 12621 20485 12633 20519
rect 12667 20516 12679 20519
rect 14274 20516 14280 20528
rect 12667 20488 14280 20516
rect 12667 20485 12679 20488
rect 12621 20479 12679 20485
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 20165 20519 20223 20525
rect 20165 20485 20177 20519
rect 20211 20516 20223 20519
rect 22186 20516 22192 20528
rect 20211 20488 22192 20516
rect 20211 20485 20223 20488
rect 20165 20479 20223 20485
rect 22186 20476 22192 20488
rect 22244 20476 22250 20528
rect 13265 20451 13323 20457
rect 11992 20420 13032 20448
rect 11885 20411 11943 20417
rect 10336 20352 10640 20380
rect 2774 20272 2780 20324
rect 2832 20312 2838 20324
rect 7190 20312 7196 20324
rect 2832 20284 7196 20312
rect 2832 20272 2838 20284
rect 7190 20272 7196 20284
rect 7248 20272 7254 20324
rect 7745 20315 7803 20321
rect 7745 20281 7757 20315
rect 7791 20312 7803 20315
rect 8757 20315 8815 20321
rect 7791 20284 8432 20312
rect 7791 20281 7803 20284
rect 7745 20275 7803 20281
rect 5258 20204 5264 20256
rect 5316 20244 5322 20256
rect 5445 20247 5503 20253
rect 5445 20244 5457 20247
rect 5316 20216 5457 20244
rect 5316 20204 5322 20216
rect 5445 20213 5457 20216
rect 5491 20213 5503 20247
rect 5445 20207 5503 20213
rect 5994 20204 6000 20256
rect 6052 20244 6058 20256
rect 6181 20247 6239 20253
rect 6181 20244 6193 20247
rect 6052 20216 6193 20244
rect 6052 20204 6058 20216
rect 6181 20213 6193 20216
rect 6227 20213 6239 20247
rect 6181 20207 6239 20213
rect 6270 20204 6276 20256
rect 6328 20244 6334 20256
rect 6328 20216 6373 20244
rect 6328 20204 6334 20216
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7377 20247 7435 20253
rect 7377 20244 7389 20247
rect 6972 20216 7389 20244
rect 6972 20204 6978 20216
rect 7377 20213 7389 20216
rect 7423 20213 7435 20247
rect 7377 20207 7435 20213
rect 7837 20247 7895 20253
rect 7837 20213 7849 20247
rect 7883 20244 7895 20247
rect 8294 20244 8300 20256
rect 7883 20216 8300 20244
rect 7883 20213 7895 20216
rect 7837 20207 7895 20213
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 8404 20253 8432 20284
rect 8757 20281 8769 20315
rect 8803 20312 8815 20315
rect 9398 20312 9404 20324
rect 8803 20284 9404 20312
rect 8803 20281 8815 20284
rect 8757 20275 8815 20281
rect 9398 20272 9404 20284
rect 9456 20272 9462 20324
rect 10612 20312 10640 20352
rect 10686 20340 10692 20392
rect 10744 20380 10750 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 10744 20352 11713 20380
rect 10744 20340 10750 20352
rect 11701 20349 11713 20352
rect 11747 20349 11759 20383
rect 13004 20380 13032 20420
rect 13265 20417 13277 20451
rect 13311 20448 13323 20451
rect 13354 20448 13360 20460
rect 13311 20420 13360 20448
rect 13311 20417 13323 20420
rect 13265 20411 13323 20417
rect 13354 20408 13360 20420
rect 13412 20408 13418 20460
rect 13633 20383 13691 20389
rect 13633 20380 13645 20383
rect 13004 20352 13645 20380
rect 11701 20343 11759 20349
rect 13633 20349 13645 20352
rect 13679 20349 13691 20383
rect 13633 20343 13691 20349
rect 14642 20340 14648 20392
rect 14700 20380 14706 20392
rect 14829 20383 14887 20389
rect 14829 20380 14841 20383
rect 14700 20352 14841 20380
rect 14700 20340 14706 20352
rect 14829 20349 14841 20352
rect 14875 20349 14887 20383
rect 14829 20343 14887 20349
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15749 20383 15807 20389
rect 15749 20380 15761 20383
rect 15252 20352 15761 20380
rect 15252 20340 15258 20352
rect 15749 20349 15761 20352
rect 15795 20349 15807 20383
rect 15749 20343 15807 20349
rect 16390 20340 16396 20392
rect 16448 20380 16454 20392
rect 16485 20383 16543 20389
rect 16485 20380 16497 20383
rect 16448 20352 16497 20380
rect 16448 20340 16454 20352
rect 16485 20349 16497 20352
rect 16531 20349 16543 20383
rect 16485 20343 16543 20349
rect 19337 20383 19395 20389
rect 19337 20349 19349 20383
rect 19383 20380 19395 20383
rect 19518 20380 19524 20392
rect 19383 20352 19524 20380
rect 19383 20349 19395 20352
rect 19337 20343 19395 20349
rect 19518 20340 19524 20352
rect 19576 20340 19582 20392
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20070 20380 20076 20392
rect 20027 20352 20076 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 20533 20383 20591 20389
rect 20533 20380 20545 20383
rect 20220 20352 20545 20380
rect 20220 20340 20226 20352
rect 20533 20349 20545 20352
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 13081 20315 13139 20321
rect 13081 20312 13093 20315
rect 10612 20284 13093 20312
rect 13081 20281 13093 20284
rect 13127 20281 13139 20315
rect 13906 20312 13912 20324
rect 13867 20284 13912 20312
rect 13081 20275 13139 20281
rect 13906 20272 13912 20284
rect 13964 20272 13970 20324
rect 8389 20247 8447 20253
rect 8389 20213 8401 20247
rect 8435 20213 8447 20247
rect 8846 20244 8852 20256
rect 8759 20216 8852 20244
rect 8389 20207 8447 20213
rect 8846 20204 8852 20216
rect 8904 20244 8910 20256
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 8904 20216 10701 20244
rect 8904 20204 8910 20216
rect 10689 20213 10701 20216
rect 10735 20213 10747 20247
rect 11330 20244 11336 20256
rect 11291 20216 11336 20244
rect 10689 20207 10747 20213
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 11698 20204 11704 20256
rect 11756 20244 11762 20256
rect 11793 20247 11851 20253
rect 11793 20244 11805 20247
rect 11756 20216 11805 20244
rect 11756 20204 11762 20216
rect 11793 20213 11805 20216
rect 11839 20213 11851 20247
rect 12986 20244 12992 20256
rect 12947 20216 12992 20244
rect 11793 20207 11851 20213
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1854 20000 1860 20052
rect 1912 20040 1918 20052
rect 1949 20043 2007 20049
rect 1949 20040 1961 20043
rect 1912 20012 1961 20040
rect 1912 20000 1918 20012
rect 1949 20009 1961 20012
rect 1995 20009 2007 20043
rect 3050 20040 3056 20052
rect 3011 20012 3056 20040
rect 1949 20003 2007 20009
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3786 20000 3792 20052
rect 3844 20040 3850 20052
rect 7374 20040 7380 20052
rect 3844 20012 5948 20040
rect 7335 20012 7380 20040
rect 3844 20000 3850 20012
rect 4608 19975 4666 19981
rect 4608 19941 4620 19975
rect 4654 19972 4666 19975
rect 5258 19972 5264 19984
rect 4654 19944 5264 19972
rect 4654 19941 4666 19944
rect 4608 19935 4666 19941
rect 5258 19932 5264 19944
rect 5316 19932 5322 19984
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 1765 19867 1823 19873
rect 1780 19836 1808 19867
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 2869 19907 2927 19913
rect 2869 19904 2881 19907
rect 2832 19876 2881 19904
rect 2832 19864 2838 19876
rect 2869 19873 2881 19876
rect 2915 19873 2927 19907
rect 5920 19904 5948 20012
rect 7374 20000 7380 20012
rect 7432 20000 7438 20052
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 9033 20043 9091 20049
rect 9033 20040 9045 20043
rect 8260 20012 9045 20040
rect 8260 20000 8266 20012
rect 9033 20009 9045 20012
rect 9079 20009 9091 20043
rect 9858 20040 9864 20052
rect 9819 20012 9864 20040
rect 9033 20003 9091 20009
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 14734 20040 14740 20052
rect 11388 20012 14740 20040
rect 11388 20000 11394 20012
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 14829 20043 14887 20049
rect 14829 20009 14841 20043
rect 14875 20040 14887 20043
rect 15470 20040 15476 20052
rect 14875 20012 15476 20040
rect 14875 20009 14887 20012
rect 14829 20003 14887 20009
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 17402 20040 17408 20052
rect 16531 20012 17408 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 17773 20043 17831 20049
rect 17773 20009 17785 20043
rect 17819 20040 17831 20043
rect 17862 20040 17868 20052
rect 17819 20012 17868 20040
rect 17819 20009 17831 20012
rect 17773 20003 17831 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 18785 20043 18843 20049
rect 18785 20009 18797 20043
rect 18831 20040 18843 20043
rect 19794 20040 19800 20052
rect 18831 20012 19800 20040
rect 18831 20009 18843 20012
rect 18785 20003 18843 20009
rect 19794 20000 19800 20012
rect 19852 20000 19858 20052
rect 19886 20000 19892 20052
rect 19944 20040 19950 20052
rect 20438 20040 20444 20052
rect 19944 20012 19989 20040
rect 20399 20012 20444 20040
rect 19944 20000 19950 20012
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 21082 20040 21088 20052
rect 21043 20012 21088 20040
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 6264 19975 6322 19981
rect 6264 19941 6276 19975
rect 6310 19972 6322 19975
rect 6362 19972 6368 19984
rect 6310 19944 6368 19972
rect 6310 19941 6322 19944
rect 6264 19935 6322 19941
rect 6362 19932 6368 19944
rect 6420 19932 6426 19984
rect 7920 19975 7978 19981
rect 7920 19941 7932 19975
rect 7966 19972 7978 19975
rect 9306 19972 9312 19984
rect 7966 19944 9312 19972
rect 7966 19941 7978 19944
rect 7920 19935 7978 19941
rect 9306 19932 9312 19944
rect 9364 19932 9370 19984
rect 10594 19981 10600 19984
rect 10588 19972 10600 19981
rect 10555 19944 10600 19972
rect 10588 19935 10600 19944
rect 10594 19932 10600 19935
rect 10652 19932 10658 19984
rect 10962 19932 10968 19984
rect 11020 19972 11026 19984
rect 11793 19975 11851 19981
rect 11793 19972 11805 19975
rect 11020 19944 11805 19972
rect 11020 19932 11026 19944
rect 11793 19941 11805 19944
rect 11839 19972 11851 19975
rect 12244 19975 12302 19981
rect 12244 19972 12256 19975
rect 11839 19944 12256 19972
rect 11839 19941 11851 19944
rect 11793 19935 11851 19941
rect 12244 19941 12256 19944
rect 12290 19972 12302 19975
rect 14182 19972 14188 19984
rect 12290 19944 14188 19972
rect 12290 19941 12302 19944
rect 12244 19935 12302 19941
rect 14182 19932 14188 19944
rect 14240 19972 14246 19984
rect 14240 19944 14320 19972
rect 14240 19932 14246 19944
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5920 19876 6009 19904
rect 2869 19867 2927 19873
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 5997 19867 6055 19873
rect 6638 19864 6644 19916
rect 6696 19904 6702 19916
rect 6696 19876 7696 19904
rect 6696 19864 6702 19876
rect 7668 19848 7696 19876
rect 9030 19864 9036 19916
rect 9088 19904 9094 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9088 19876 9689 19904
rect 9088 19864 9094 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 10321 19907 10379 19913
rect 10321 19873 10333 19907
rect 10367 19904 10379 19907
rect 14001 19907 14059 19913
rect 10367 19876 11560 19904
rect 10367 19873 10379 19876
rect 10321 19867 10379 19873
rect 3694 19836 3700 19848
rect 1780 19808 3700 19836
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 3786 19796 3792 19848
rect 3844 19836 3850 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 3844 19808 4353 19836
rect 3844 19796 3850 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 7650 19836 7656 19848
rect 7611 19808 7656 19836
rect 4341 19799 4399 19805
rect 7650 19796 7656 19808
rect 7708 19796 7714 19848
rect 11532 19836 11560 19876
rect 14001 19873 14013 19907
rect 14047 19873 14059 19907
rect 14001 19867 14059 19873
rect 11974 19836 11980 19848
rect 11532 19808 11980 19836
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 11701 19771 11759 19777
rect 11701 19737 11713 19771
rect 11747 19768 11759 19771
rect 11793 19771 11851 19777
rect 11793 19768 11805 19771
rect 11747 19740 11805 19768
rect 11747 19737 11759 19740
rect 11701 19731 11759 19737
rect 11793 19737 11805 19740
rect 11839 19737 11851 19771
rect 13633 19771 13691 19777
rect 13633 19768 13645 19771
rect 11793 19731 11851 19737
rect 13004 19740 13645 19768
rect 2501 19703 2559 19709
rect 2501 19669 2513 19703
rect 2547 19700 2559 19703
rect 2866 19700 2872 19712
rect 2547 19672 2872 19700
rect 2547 19669 2559 19672
rect 2501 19663 2559 19669
rect 2866 19660 2872 19672
rect 2924 19660 2930 19712
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 5721 19703 5779 19709
rect 5721 19700 5733 19703
rect 4120 19672 5733 19700
rect 4120 19660 4126 19672
rect 5721 19669 5733 19672
rect 5767 19669 5779 19703
rect 5721 19663 5779 19669
rect 5810 19660 5816 19712
rect 5868 19700 5874 19712
rect 12250 19700 12256 19712
rect 5868 19672 12256 19700
rect 5868 19660 5874 19672
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12342 19660 12348 19712
rect 12400 19700 12406 19712
rect 13004 19700 13032 19740
rect 13633 19737 13645 19740
rect 13679 19737 13691 19771
rect 13633 19731 13691 19737
rect 14016 19712 14044 19867
rect 14292 19845 14320 19944
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 17092 19944 18644 19972
rect 17092 19932 17098 19944
rect 14645 19907 14703 19913
rect 14645 19873 14657 19907
rect 14691 19904 14703 19907
rect 15378 19904 15384 19916
rect 14691 19876 15384 19904
rect 14691 19873 14703 19876
rect 14645 19867 14703 19873
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 15562 19904 15568 19916
rect 15523 19876 15568 19904
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15841 19907 15899 19913
rect 15841 19873 15853 19907
rect 15887 19904 15899 19907
rect 16301 19907 16359 19913
rect 16301 19904 16313 19907
rect 15887 19876 16313 19904
rect 15887 19873 15899 19876
rect 15841 19867 15899 19873
rect 16301 19873 16313 19876
rect 16347 19873 16359 19907
rect 16301 19867 16359 19873
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 18616 19913 18644 19944
rect 16853 19907 16911 19913
rect 16853 19904 16865 19907
rect 16632 19876 16865 19904
rect 16632 19864 16638 19876
rect 16853 19873 16865 19876
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19873 17647 19907
rect 17589 19867 17647 19873
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19873 18659 19907
rect 19150 19904 19156 19916
rect 19111 19876 19156 19904
rect 18601 19867 18659 19873
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 17604 19836 17632 19867
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19873 19763 19907
rect 20254 19904 20260 19916
rect 20215 19876 20260 19904
rect 19705 19867 19763 19873
rect 14277 19799 14335 19805
rect 14568 19808 17632 19836
rect 19720 19836 19748 19867
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19904 20959 19907
rect 21269 19907 21327 19913
rect 21269 19904 21281 19907
rect 20947 19876 21281 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 21269 19873 21281 19876
rect 21315 19873 21327 19907
rect 21269 19867 21327 19873
rect 20438 19836 20444 19848
rect 19720 19808 20444 19836
rect 14108 19768 14136 19799
rect 14458 19768 14464 19780
rect 14108 19740 14464 19768
rect 14458 19728 14464 19740
rect 14516 19728 14522 19780
rect 13354 19700 13360 19712
rect 12400 19672 13032 19700
rect 13315 19672 13360 19700
rect 12400 19660 12406 19672
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13998 19700 14004 19712
rect 13911 19672 14004 19700
rect 13998 19660 14004 19672
rect 14056 19700 14062 19712
rect 14568 19700 14596 19808
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 17037 19771 17095 19777
rect 17037 19737 17049 19771
rect 17083 19768 17095 19771
rect 17954 19768 17960 19780
rect 17083 19740 17960 19768
rect 17083 19737 17095 19740
rect 17037 19731 17095 19737
rect 17954 19728 17960 19740
rect 18012 19728 18018 19780
rect 19337 19771 19395 19777
rect 19337 19737 19349 19771
rect 19383 19768 19395 19771
rect 20714 19768 20720 19780
rect 19383 19740 20720 19768
rect 19383 19737 19395 19740
rect 19337 19731 19395 19737
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 14056 19672 14596 19700
rect 14056 19660 14062 19672
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 6270 19496 6276 19508
rect 5767 19468 6276 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 6380 19468 7788 19496
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 6380 19428 6408 19468
rect 2547 19400 4844 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 3237 19363 3295 19369
rect 1688 19332 3188 19360
rect 658 19252 664 19304
rect 716 19292 722 19304
rect 1688 19292 1716 19332
rect 716 19264 1716 19292
rect 1765 19295 1823 19301
rect 716 19252 722 19264
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2501 19295 2559 19301
rect 2501 19292 2513 19295
rect 1811 19264 2513 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2501 19261 2513 19264
rect 2547 19261 2559 19295
rect 2501 19255 2559 19261
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 3160 19292 3188 19332
rect 3237 19329 3249 19363
rect 3283 19360 3295 19363
rect 3510 19360 3516 19372
rect 3283 19332 3516 19360
rect 3283 19329 3295 19332
rect 3237 19323 3295 19329
rect 3510 19320 3516 19332
rect 3568 19360 3574 19372
rect 4062 19360 4068 19372
rect 3568 19332 4068 19360
rect 3568 19320 3574 19332
rect 4062 19320 4068 19332
rect 4120 19360 4126 19372
rect 4157 19363 4215 19369
rect 4157 19360 4169 19363
rect 4120 19332 4169 19360
rect 4120 19320 4126 19332
rect 4157 19329 4169 19332
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 4816 19304 4844 19400
rect 6196 19400 6408 19428
rect 5258 19360 5264 19372
rect 5219 19332 5264 19360
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 2648 19264 3004 19292
rect 3160 19264 4752 19292
rect 2648 19252 2654 19264
rect 2866 19224 2872 19236
rect 1964 19196 2872 19224
rect 1964 19165 1992 19196
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 2976 19224 3004 19264
rect 3053 19227 3111 19233
rect 3053 19224 3065 19227
rect 2963 19196 3065 19224
rect 3053 19193 3065 19196
rect 3099 19224 3111 19227
rect 4522 19224 4528 19236
rect 3099 19196 4528 19224
rect 3099 19193 3111 19196
rect 3053 19187 3111 19193
rect 4522 19184 4528 19196
rect 4580 19184 4586 19236
rect 4724 19224 4752 19264
rect 4798 19252 4804 19304
rect 4856 19252 4862 19304
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5166 19292 5172 19304
rect 5123 19264 5172 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 6196 19292 6224 19400
rect 6454 19388 6460 19440
rect 6512 19428 6518 19440
rect 6822 19428 6828 19440
rect 6512 19400 6828 19428
rect 6512 19388 6518 19400
rect 6822 19388 6828 19400
rect 6880 19388 6886 19440
rect 7760 19428 7788 19468
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 8481 19499 8539 19505
rect 8481 19496 8493 19499
rect 8352 19468 8493 19496
rect 8352 19456 8358 19468
rect 8481 19465 8493 19468
rect 8527 19465 8539 19499
rect 8481 19459 8539 19465
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 10965 19499 11023 19505
rect 10008 19468 10824 19496
rect 10008 19456 10014 19468
rect 10796 19428 10824 19468
rect 10965 19465 10977 19499
rect 11011 19496 11023 19499
rect 11054 19496 11060 19508
rect 11011 19468 11060 19496
rect 11011 19465 11023 19468
rect 10965 19459 11023 19465
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11974 19456 11980 19508
rect 12032 19496 12038 19508
rect 12253 19499 12311 19505
rect 12253 19496 12265 19499
rect 12032 19468 12265 19496
rect 12032 19456 12038 19468
rect 12253 19465 12265 19468
rect 12299 19465 12311 19499
rect 13814 19496 13820 19508
rect 13727 19468 13820 19496
rect 12253 19459 12311 19465
rect 13814 19456 13820 19468
rect 13872 19496 13878 19508
rect 20990 19496 20996 19508
rect 13872 19468 14688 19496
rect 20951 19468 20996 19496
rect 13872 19456 13878 19468
rect 11422 19428 11428 19440
rect 7760 19400 8340 19428
rect 10796 19400 11428 19428
rect 6362 19360 6368 19372
rect 6275 19332 6368 19360
rect 6362 19320 6368 19332
rect 6420 19360 6426 19372
rect 6420 19332 6960 19360
rect 6420 19320 6426 19332
rect 6104 19264 6224 19292
rect 4985 19227 5043 19233
rect 4985 19224 4997 19227
rect 4724 19196 4997 19224
rect 4985 19193 4997 19196
rect 5031 19224 5043 19227
rect 6104 19224 6132 19264
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6696 19264 6837 19292
rect 6696 19252 6702 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6932 19292 6960 19332
rect 8312 19292 8340 19400
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 12342 19428 12348 19440
rect 11808 19400 12348 19428
rect 9125 19363 9183 19369
rect 9125 19329 9137 19363
rect 9171 19360 9183 19363
rect 9306 19360 9312 19372
rect 9171 19332 9312 19360
rect 9171 19329 9183 19332
rect 9125 19323 9183 19329
rect 9306 19320 9312 19332
rect 9364 19320 9370 19372
rect 11808 19369 11836 19400
rect 12342 19388 12348 19400
rect 12400 19388 12406 19440
rect 14660 19369 14688 19468
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19329 11851 19363
rect 11793 19323 11851 19329
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 14645 19363 14703 19369
rect 12023 19332 12572 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 12544 19304 12572 19332
rect 14645 19329 14657 19363
rect 14691 19329 14703 19363
rect 14645 19323 14703 19329
rect 16298 19320 16304 19372
rect 16356 19360 16362 19372
rect 16356 19332 16988 19360
rect 16356 19320 16362 19332
rect 8941 19295 8999 19301
rect 8941 19292 8953 19295
rect 6932 19264 8248 19292
rect 8312 19264 8953 19292
rect 6825 19255 6883 19261
rect 5031 19196 6132 19224
rect 6181 19227 6239 19233
rect 5031 19193 5043 19196
rect 4985 19187 5043 19193
rect 6181 19193 6193 19227
rect 6227 19224 6239 19227
rect 6914 19224 6920 19236
rect 6227 19196 6920 19224
rect 6227 19193 6239 19196
rect 6181 19187 6239 19193
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 7092 19227 7150 19233
rect 7092 19193 7104 19227
rect 7138 19224 7150 19227
rect 7558 19224 7564 19236
rect 7138 19196 7564 19224
rect 7138 19193 7150 19196
rect 7092 19187 7150 19193
rect 7558 19184 7564 19196
rect 7616 19224 7622 19236
rect 8110 19224 8116 19236
rect 7616 19196 8116 19224
rect 7616 19184 7622 19196
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 1949 19159 2007 19165
rect 1949 19125 1961 19159
rect 1995 19125 2007 19159
rect 2590 19156 2596 19168
rect 2551 19128 2596 19156
rect 1949 19119 2007 19125
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 3142 19156 3148 19168
rect 3007 19128 3148 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 3142 19116 3148 19128
rect 3200 19116 3206 19168
rect 3602 19156 3608 19168
rect 3563 19128 3608 19156
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3878 19116 3884 19168
rect 3936 19156 3942 19168
rect 3973 19159 4031 19165
rect 3973 19156 3985 19159
rect 3936 19128 3985 19156
rect 3936 19116 3942 19128
rect 3973 19125 3985 19128
rect 4019 19125 4031 19159
rect 3973 19119 4031 19125
rect 4065 19159 4123 19165
rect 4065 19125 4077 19159
rect 4111 19156 4123 19159
rect 4617 19159 4675 19165
rect 4617 19156 4629 19159
rect 4111 19128 4629 19156
rect 4111 19125 4123 19128
rect 4065 19119 4123 19125
rect 4617 19125 4629 19128
rect 4663 19125 4675 19159
rect 4617 19119 4675 19125
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 5810 19156 5816 19168
rect 4856 19128 5816 19156
rect 4856 19116 4862 19128
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 6089 19159 6147 19165
rect 6089 19125 6101 19159
rect 6135 19156 6147 19159
rect 7742 19156 7748 19168
rect 6135 19128 7748 19156
rect 6135 19125 6147 19128
rect 6089 19119 6147 19125
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 8220 19165 8248 19264
rect 8941 19261 8953 19264
rect 8987 19261 8999 19295
rect 8941 19255 8999 19261
rect 8956 19224 8984 19255
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 9490 19292 9496 19304
rect 9272 19264 9496 19292
rect 9272 19252 9278 19264
rect 9490 19252 9496 19264
rect 9548 19292 9554 19304
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 9548 19264 9597 19292
rect 9548 19252 9554 19264
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 10410 19292 10416 19304
rect 9585 19255 9643 19261
rect 9692 19264 10416 19292
rect 9692 19224 9720 19264
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12299 19264 12449 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 12693 19295 12751 19301
rect 12693 19292 12705 19295
rect 12584 19264 12705 19292
rect 12584 19252 12590 19264
rect 12693 19261 12705 19264
rect 12739 19261 12751 19295
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 12693 19255 12751 19261
rect 12820 19264 14473 19292
rect 8956 19196 9720 19224
rect 9852 19227 9910 19233
rect 9852 19193 9864 19227
rect 9898 19224 9910 19227
rect 11146 19224 11152 19236
rect 9898 19196 11152 19224
rect 9898 19193 9910 19196
rect 9852 19187 9910 19193
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 12820 19224 12848 19264
rect 14461 19261 14473 19264
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14792 19264 15117 19292
rect 14792 19252 14798 19264
rect 15105 19261 15117 19264
rect 15151 19261 15163 19295
rect 15378 19292 15384 19304
rect 15339 19264 15384 19292
rect 15105 19255 15163 19261
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 15933 19295 15991 19301
rect 15933 19261 15945 19295
rect 15979 19292 15991 19295
rect 16114 19292 16120 19304
rect 15979 19264 16120 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16209 19295 16267 19301
rect 16209 19261 16221 19295
rect 16255 19292 16267 19295
rect 16574 19292 16580 19304
rect 16255 19264 16580 19292
rect 16255 19261 16267 19264
rect 16209 19255 16267 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 16666 19252 16672 19304
rect 16724 19292 16730 19304
rect 16960 19292 16988 19332
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 16724 19264 16769 19292
rect 16960 19264 17417 19292
rect 16724 19252 16730 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 11348 19196 11928 19224
rect 8205 19159 8263 19165
rect 8205 19125 8217 19159
rect 8251 19125 8263 19159
rect 8205 19119 8263 19125
rect 8662 19116 8668 19168
rect 8720 19156 8726 19168
rect 8849 19159 8907 19165
rect 8849 19156 8861 19159
rect 8720 19128 8861 19156
rect 8720 19116 8726 19128
rect 8849 19125 8861 19128
rect 8895 19156 8907 19159
rect 11238 19156 11244 19168
rect 8895 19128 11244 19156
rect 8895 19125 8907 19128
rect 8849 19119 8907 19125
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 11348 19165 11376 19196
rect 11333 19159 11391 19165
rect 11333 19125 11345 19159
rect 11379 19125 11391 19159
rect 11333 19119 11391 19125
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19156 11759 19159
rect 11790 19156 11796 19168
rect 11747 19128 11796 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 11900 19156 11928 19196
rect 12728 19196 12848 19224
rect 12728 19156 12756 19196
rect 14274 19184 14280 19236
rect 14332 19224 14338 19236
rect 14553 19227 14611 19233
rect 14553 19224 14565 19227
rect 14332 19196 14565 19224
rect 14332 19184 14338 19196
rect 14553 19193 14565 19196
rect 14599 19193 14611 19227
rect 14553 19187 14611 19193
rect 16022 19184 16028 19236
rect 16080 19224 16086 19236
rect 18064 19224 18092 19255
rect 18230 19252 18236 19304
rect 18288 19292 18294 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 18288 19264 19165 19292
rect 18288 19252 18294 19264
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 19705 19295 19763 19301
rect 19705 19261 19717 19295
rect 19751 19292 19763 19295
rect 19794 19292 19800 19304
rect 19751 19264 19800 19292
rect 19751 19261 19763 19264
rect 19705 19255 19763 19261
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 20254 19292 20260 19304
rect 20215 19264 20260 19292
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 20364 19264 20576 19292
rect 16080 19196 18092 19224
rect 16080 19184 16086 19196
rect 11900 19128 12756 19156
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 13446 19156 13452 19168
rect 12860 19128 13452 19156
rect 12860 19116 12866 19128
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 14093 19159 14151 19165
rect 14093 19125 14105 19159
rect 14139 19156 14151 19159
rect 14366 19156 14372 19168
rect 14139 19128 14372 19156
rect 14139 19125 14151 19128
rect 14093 19119 14151 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 16482 19116 16488 19168
rect 16540 19156 16546 19168
rect 16853 19159 16911 19165
rect 16853 19156 16865 19159
rect 16540 19128 16865 19156
rect 16540 19116 16546 19128
rect 16853 19125 16865 19128
rect 16899 19125 16911 19159
rect 16853 19119 16911 19125
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19156 17647 19159
rect 18138 19156 18144 19168
rect 17635 19128 18144 19156
rect 17635 19125 17647 19128
rect 17589 19119 17647 19125
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18874 19156 18880 19168
rect 18279 19128 18880 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 19337 19159 19395 19165
rect 19337 19125 19349 19159
rect 19383 19156 19395 19159
rect 19426 19156 19432 19168
rect 19383 19128 19432 19156
rect 19383 19125 19395 19128
rect 19337 19119 19395 19125
rect 19426 19116 19432 19128
rect 19484 19116 19490 19168
rect 19889 19159 19947 19165
rect 19889 19125 19901 19159
rect 19935 19156 19947 19159
rect 20364 19156 20392 19264
rect 20548 19224 20576 19264
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20772 19264 20821 19292
rect 20772 19252 20778 19264
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 21266 19224 21272 19236
rect 20548 19196 21272 19224
rect 21266 19184 21272 19196
rect 21324 19184 21330 19236
rect 19935 19128 20392 19156
rect 20441 19159 20499 19165
rect 19935 19125 19947 19128
rect 19889 19119 19947 19125
rect 20441 19125 20453 19159
rect 20487 19156 20499 19159
rect 20530 19156 20536 19168
rect 20487 19128 20536 19156
rect 20487 19125 20499 19128
rect 20441 19119 20499 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1854 18952 1860 18964
rect 1815 18924 1860 18952
rect 1854 18912 1860 18924
rect 1912 18912 1918 18964
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18921 3019 18955
rect 2961 18915 3019 18921
rect 1762 18844 1768 18896
rect 1820 18884 1826 18896
rect 2501 18887 2559 18893
rect 2501 18884 2513 18887
rect 1820 18856 2513 18884
rect 1820 18844 1826 18856
rect 2501 18853 2513 18856
rect 2547 18853 2559 18887
rect 2976 18884 3004 18915
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 3292 18924 3341 18952
rect 3292 18912 3298 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 3329 18915 3387 18921
rect 3602 18912 3608 18964
rect 3660 18952 3666 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 3660 18924 4537 18952
rect 3660 18912 3666 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 4525 18915 4583 18921
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 5994 18952 6000 18964
rect 5767 18924 6000 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 5994 18912 6000 18924
rect 6052 18912 6058 18964
rect 6181 18955 6239 18961
rect 6181 18921 6193 18955
rect 6227 18952 6239 18955
rect 6917 18955 6975 18961
rect 6917 18952 6929 18955
rect 6227 18924 6929 18952
rect 6227 18921 6239 18924
rect 6181 18915 6239 18921
rect 6917 18921 6929 18924
rect 6963 18921 6975 18955
rect 6917 18915 6975 18921
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 9677 18955 9735 18961
rect 7064 18924 9628 18952
rect 7064 18912 7070 18924
rect 4433 18887 4491 18893
rect 4433 18884 4445 18887
rect 2976 18856 4445 18884
rect 2501 18847 2559 18853
rect 4433 18853 4445 18856
rect 4479 18853 4491 18887
rect 4433 18847 4491 18853
rect 4614 18844 4620 18896
rect 4672 18884 4678 18896
rect 8846 18884 8852 18896
rect 4672 18856 8852 18884
rect 4672 18844 4678 18856
rect 8846 18844 8852 18856
rect 8904 18844 8910 18896
rect 9600 18884 9628 18924
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 11149 18955 11207 18961
rect 11149 18952 11161 18955
rect 9723 18924 11161 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 11149 18921 11161 18924
rect 11195 18921 11207 18955
rect 13906 18952 13912 18964
rect 11149 18915 11207 18921
rect 12452 18924 13912 18952
rect 12158 18884 12164 18896
rect 9600 18856 12164 18884
rect 12158 18844 12164 18856
rect 12216 18844 12222 18896
rect 1670 18816 1676 18828
rect 1631 18788 1676 18816
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2225 18819 2283 18825
rect 2225 18816 2237 18819
rect 2096 18788 2237 18816
rect 2096 18776 2102 18788
rect 2225 18785 2237 18788
rect 2271 18785 2283 18819
rect 2225 18779 2283 18785
rect 2777 18819 2835 18825
rect 2777 18785 2789 18819
rect 2823 18816 2835 18819
rect 3878 18816 3884 18828
rect 2823 18788 3884 18816
rect 2823 18785 2835 18788
rect 2777 18779 2835 18785
rect 3878 18776 3884 18788
rect 3936 18816 3942 18828
rect 4062 18816 4068 18828
rect 3936 18788 4068 18816
rect 3936 18776 3942 18788
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 5077 18819 5135 18825
rect 5077 18785 5089 18819
rect 5123 18816 5135 18819
rect 5534 18816 5540 18828
rect 5123 18788 5540 18816
rect 5123 18785 5135 18788
rect 5077 18779 5135 18785
rect 5534 18776 5540 18788
rect 5592 18776 5598 18828
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18816 6147 18819
rect 6822 18816 6828 18828
rect 6135 18788 6828 18816
rect 6135 18785 6147 18788
rect 6089 18779 6147 18785
rect 6822 18776 6828 18788
rect 6880 18776 6886 18828
rect 7285 18819 7343 18825
rect 7285 18816 7297 18819
rect 6932 18788 7297 18816
rect 1578 18708 1584 18760
rect 1636 18748 1642 18760
rect 3421 18751 3479 18757
rect 3421 18748 3433 18751
rect 1636 18720 3433 18748
rect 1636 18708 1642 18720
rect 3421 18717 3433 18720
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18717 3663 18751
rect 3605 18711 3663 18717
rect 1118 18640 1124 18692
rect 1176 18680 1182 18692
rect 2777 18683 2835 18689
rect 2777 18680 2789 18683
rect 1176 18652 2789 18680
rect 1176 18640 1182 18652
rect 2777 18649 2789 18652
rect 2823 18649 2835 18683
rect 2777 18643 2835 18649
rect 3436 18612 3464 18711
rect 3510 18640 3516 18692
rect 3568 18680 3574 18692
rect 3620 18680 3648 18711
rect 3694 18708 3700 18760
rect 3752 18748 3758 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 3752 18720 4629 18748
rect 3752 18708 3758 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 5350 18748 5356 18760
rect 5311 18720 5356 18748
rect 4617 18711 4675 18717
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 6362 18748 6368 18760
rect 6323 18720 6368 18748
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18748 6699 18751
rect 6932 18748 6960 18788
rect 7285 18785 7297 18788
rect 7331 18785 7343 18819
rect 7285 18779 7343 18785
rect 8202 18776 8208 18828
rect 8260 18816 8266 18828
rect 8757 18819 8815 18825
rect 8260 18788 8432 18816
rect 8260 18776 8266 18788
rect 7374 18748 7380 18760
rect 6687 18720 6960 18748
rect 7335 18720 7380 18748
rect 6687 18717 6699 18720
rect 6641 18711 6699 18717
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 7558 18748 7564 18760
rect 7519 18720 7564 18748
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7926 18748 7932 18760
rect 7887 18720 7932 18748
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 8404 18748 8432 18788
rect 8757 18785 8769 18819
rect 8803 18816 8815 18819
rect 9582 18816 9588 18828
rect 8803 18788 9588 18816
rect 8803 18785 8815 18788
rect 8757 18779 8815 18785
rect 9582 18776 9588 18788
rect 9640 18776 9646 18828
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10870 18816 10876 18828
rect 10091 18788 10876 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 11054 18816 11060 18828
rect 11015 18788 11060 18816
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11701 18819 11759 18825
rect 11701 18785 11713 18819
rect 11747 18816 11759 18819
rect 12452 18816 12480 18924
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 14366 18952 14372 18964
rect 14327 18924 14372 18952
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 15378 18912 15384 18964
rect 15436 18952 15442 18964
rect 18230 18952 18236 18964
rect 15436 18924 18236 18952
rect 15436 18912 15442 18924
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 18509 18955 18567 18961
rect 18509 18921 18521 18955
rect 18555 18952 18567 18955
rect 19334 18952 19340 18964
rect 18555 18924 19340 18952
rect 18555 18921 18567 18924
rect 18509 18915 18567 18921
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 21082 18952 21088 18964
rect 21043 18924 21088 18952
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 12520 18887 12578 18893
rect 12520 18853 12532 18887
rect 12566 18884 12578 18887
rect 13814 18884 13820 18896
rect 12566 18856 13820 18884
rect 12566 18853 12578 18856
rect 12520 18847 12578 18853
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 13998 18844 14004 18896
rect 14056 18884 14062 18896
rect 15286 18884 15292 18896
rect 14056 18856 15292 18884
rect 14056 18844 14062 18856
rect 15286 18844 15292 18856
rect 15344 18884 15350 18896
rect 18690 18884 18696 18896
rect 15344 18856 18696 18884
rect 15344 18844 15350 18856
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 22646 18884 22652 18896
rect 19484 18856 22652 18884
rect 19484 18844 19490 18856
rect 22646 18844 22652 18856
rect 22704 18844 22710 18896
rect 11747 18788 12480 18816
rect 11747 18785 11759 18788
rect 11701 18779 11759 18785
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 14277 18819 14335 18825
rect 14277 18816 14289 18819
rect 12860 18788 14289 18816
rect 12860 18776 12866 18788
rect 14277 18785 14289 18788
rect 14323 18785 14335 18819
rect 14277 18779 14335 18785
rect 14366 18776 14372 18828
rect 14424 18816 14430 18828
rect 17221 18819 17279 18825
rect 17221 18816 17233 18819
rect 14424 18788 17233 18816
rect 14424 18776 14430 18788
rect 17221 18785 17233 18788
rect 17267 18785 17279 18819
rect 17221 18779 17279 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18816 17555 18819
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 17543 18788 18337 18816
rect 17543 18785 17555 18788
rect 17497 18779 17555 18785
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 19702 18816 19708 18828
rect 19663 18788 19708 18816
rect 18325 18779 18383 18785
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 19886 18776 19892 18828
rect 19944 18816 19950 18828
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 19944 18788 20269 18816
rect 19944 18776 19950 18788
rect 20257 18785 20269 18788
rect 20303 18785 20315 18819
rect 20257 18779 20315 18785
rect 20622 18776 20628 18828
rect 20680 18816 20686 18828
rect 20901 18819 20959 18825
rect 20901 18816 20913 18819
rect 20680 18788 20913 18816
rect 20680 18776 20686 18788
rect 20901 18785 20913 18788
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 8849 18751 8907 18757
rect 8849 18748 8861 18751
rect 8404 18720 8861 18748
rect 8849 18717 8861 18720
rect 8895 18717 8907 18751
rect 8849 18711 8907 18717
rect 9033 18751 9091 18757
rect 9033 18717 9045 18751
rect 9079 18748 9091 18751
rect 9306 18748 9312 18760
rect 9079 18720 9312 18748
rect 9079 18717 9091 18720
rect 9033 18711 9091 18717
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 10134 18748 10140 18760
rect 10095 18720 10140 18748
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10962 18748 10968 18760
rect 10367 18720 10968 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 11146 18708 11152 18760
rect 11204 18748 11210 18760
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 11204 18720 11253 18748
rect 11204 18708 11210 18720
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 11241 18711 11299 18717
rect 11974 18708 11980 18760
rect 12032 18748 12038 18760
rect 12250 18748 12256 18760
rect 12032 18720 12256 18748
rect 12032 18708 12038 18720
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 13538 18708 13544 18760
rect 13596 18748 13602 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 13596 18720 14473 18748
rect 13596 18708 13602 18720
rect 8662 18680 8668 18692
rect 3568 18652 3648 18680
rect 3988 18652 8668 18680
rect 3568 18640 3574 18652
rect 3988 18612 4016 18652
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 8754 18640 8760 18692
rect 8812 18680 8818 18692
rect 9858 18680 9864 18692
rect 8812 18652 9864 18680
rect 8812 18640 8818 18652
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 10686 18680 10692 18692
rect 10647 18652 10692 18680
rect 10686 18640 10692 18652
rect 10744 18640 10750 18692
rect 13648 18689 13676 18720
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 20806 18748 20812 18760
rect 14461 18711 14519 18717
rect 18064 18720 20812 18748
rect 13633 18683 13691 18689
rect 13633 18649 13645 18683
rect 13679 18680 13691 18683
rect 13909 18683 13967 18689
rect 13679 18652 13713 18680
rect 13679 18649 13691 18652
rect 13633 18643 13691 18649
rect 13909 18649 13921 18683
rect 13955 18680 13967 18683
rect 15562 18680 15568 18692
rect 13955 18652 15568 18680
rect 13955 18649 13967 18652
rect 13909 18643 13967 18649
rect 15562 18640 15568 18652
rect 15620 18640 15626 18692
rect 3436 18584 4016 18612
rect 4065 18615 4123 18621
rect 4065 18581 4077 18615
rect 4111 18612 4123 18615
rect 4338 18612 4344 18624
rect 4111 18584 4344 18612
rect 4111 18581 4123 18584
rect 4065 18575 4123 18581
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 6086 18612 6092 18624
rect 5040 18584 6092 18612
rect 5040 18572 5046 18584
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 6641 18615 6699 18621
rect 6641 18581 6653 18615
rect 6687 18612 6699 18615
rect 6730 18612 6736 18624
rect 6687 18584 6736 18612
rect 6687 18581 6699 18584
rect 6641 18575 6699 18581
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 7190 18572 7196 18624
rect 7248 18612 7254 18624
rect 8202 18612 8208 18624
rect 7248 18584 8208 18612
rect 7248 18572 7254 18584
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8389 18615 8447 18621
rect 8389 18612 8401 18615
rect 8352 18584 8401 18612
rect 8352 18572 8358 18584
rect 8389 18581 8401 18584
rect 8435 18581 8447 18615
rect 8389 18575 8447 18581
rect 9122 18572 9128 18624
rect 9180 18612 9186 18624
rect 11698 18612 11704 18624
rect 9180 18584 11704 18612
rect 9180 18572 9186 18584
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 11885 18615 11943 18621
rect 11885 18581 11897 18615
rect 11931 18612 11943 18615
rect 14090 18612 14096 18624
rect 11931 18584 14096 18612
rect 11931 18581 11943 18584
rect 11885 18575 11943 18581
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14274 18572 14280 18624
rect 14332 18612 14338 18624
rect 18064 18612 18092 18720
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 19889 18683 19947 18689
rect 19889 18649 19901 18683
rect 19935 18680 19947 18683
rect 21726 18680 21732 18692
rect 19935 18652 21732 18680
rect 19935 18649 19947 18652
rect 19889 18643 19947 18649
rect 21726 18640 21732 18652
rect 21784 18640 21790 18692
rect 14332 18584 18092 18612
rect 14332 18572 14338 18584
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 19978 18612 19984 18624
rect 18196 18584 19984 18612
rect 18196 18572 18202 18584
rect 19978 18572 19984 18584
rect 20036 18612 20042 18624
rect 20254 18612 20260 18624
rect 20036 18584 20260 18612
rect 20036 18572 20042 18584
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 20346 18572 20352 18624
rect 20404 18612 20410 18624
rect 20441 18615 20499 18621
rect 20441 18612 20453 18615
rect 20404 18584 20453 18612
rect 20404 18572 20410 18584
rect 20441 18581 20453 18584
rect 20487 18581 20499 18615
rect 20441 18575 20499 18581
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2774 18408 2780 18420
rect 2547 18380 2780 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 2869 18411 2927 18417
rect 2869 18377 2881 18411
rect 2915 18408 2927 18411
rect 4798 18408 4804 18420
rect 2915 18380 4804 18408
rect 2915 18377 2927 18380
rect 2869 18371 2927 18377
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 5534 18408 5540 18420
rect 5495 18380 5540 18408
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 6822 18408 6828 18420
rect 6783 18380 6828 18408
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 7742 18368 7748 18420
rect 7800 18408 7806 18420
rect 7929 18411 7987 18417
rect 7929 18408 7941 18411
rect 7800 18380 7941 18408
rect 7800 18368 7806 18380
rect 7929 18377 7941 18380
rect 7975 18377 7987 18411
rect 7929 18371 7987 18377
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 9033 18411 9091 18417
rect 8444 18380 8984 18408
rect 8444 18368 8450 18380
rect 5261 18343 5319 18349
rect 5261 18309 5273 18343
rect 5307 18309 5319 18343
rect 5261 18303 5319 18309
rect 2590 18232 2596 18284
rect 2648 18272 2654 18284
rect 3329 18275 3387 18281
rect 3329 18272 3341 18275
rect 2648 18244 3341 18272
rect 2648 18232 2654 18244
rect 3329 18241 3341 18244
rect 3375 18241 3387 18275
rect 3329 18235 3387 18241
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18272 3571 18275
rect 3694 18272 3700 18284
rect 3559 18244 3700 18272
rect 3559 18241 3571 18244
rect 3513 18235 3571 18241
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 5276 18272 5304 18303
rect 5350 18300 5356 18352
rect 5408 18340 5414 18352
rect 8956 18340 8984 18380
rect 9033 18377 9045 18411
rect 9079 18408 9091 18411
rect 9122 18408 9128 18420
rect 9079 18380 9128 18408
rect 9079 18377 9091 18380
rect 9033 18371 9091 18377
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 10134 18408 10140 18420
rect 9600 18380 10140 18408
rect 9600 18340 9628 18380
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 11054 18408 11060 18420
rect 11015 18380 11060 18408
rect 11054 18368 11060 18380
rect 11112 18368 11118 18420
rect 12529 18411 12587 18417
rect 12529 18377 12541 18411
rect 12575 18408 12587 18411
rect 12802 18408 12808 18420
rect 12575 18380 12808 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 12986 18368 12992 18420
rect 13044 18408 13050 18420
rect 13541 18411 13599 18417
rect 13541 18408 13553 18411
rect 13044 18380 13553 18408
rect 13044 18368 13050 18380
rect 13541 18377 13553 18380
rect 13587 18377 13599 18411
rect 13541 18371 13599 18377
rect 14550 18368 14556 18420
rect 14608 18408 14614 18420
rect 14737 18411 14795 18417
rect 14737 18408 14749 18411
rect 14608 18380 14749 18408
rect 14608 18368 14614 18380
rect 14737 18377 14749 18380
rect 14783 18377 14795 18411
rect 14737 18371 14795 18377
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 19518 18408 19524 18420
rect 14884 18380 19524 18408
rect 14884 18368 14890 18380
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 21266 18408 21272 18420
rect 21227 18380 21272 18408
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 11146 18340 11152 18352
rect 5408 18312 8892 18340
rect 8956 18312 9628 18340
rect 9692 18312 11152 18340
rect 5408 18300 5414 18312
rect 5626 18272 5632 18284
rect 5276 18244 5632 18272
rect 5626 18232 5632 18244
rect 5684 18272 5690 18284
rect 6089 18275 6147 18281
rect 6089 18272 6101 18275
rect 5684 18244 6101 18272
rect 5684 18232 5690 18244
rect 6089 18241 6101 18244
rect 6135 18241 6147 18275
rect 6089 18235 6147 18241
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18272 7527 18275
rect 7558 18272 7564 18284
rect 7515 18244 7564 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 7558 18232 7564 18244
rect 7616 18272 7622 18284
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 7616 18244 8493 18272
rect 7616 18232 7622 18244
rect 8481 18241 8493 18244
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 3878 18164 3884 18216
rect 3936 18204 3942 18216
rect 5166 18204 5172 18216
rect 3936 18176 3981 18204
rect 4080 18176 5172 18204
rect 3936 18164 3942 18176
rect 2866 18096 2872 18148
rect 2924 18136 2930 18148
rect 4080 18136 4108 18176
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 7193 18207 7251 18213
rect 7193 18173 7205 18207
rect 7239 18204 7251 18207
rect 7926 18204 7932 18216
rect 7239 18176 7932 18204
rect 7239 18173 7251 18176
rect 7193 18167 7251 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 8294 18204 8300 18216
rect 8255 18176 8300 18204
rect 8294 18164 8300 18176
rect 8352 18164 8358 18216
rect 8864 18204 8892 18312
rect 9692 18281 9720 18312
rect 11146 18300 11152 18312
rect 11204 18300 11210 18352
rect 12253 18343 12311 18349
rect 12253 18309 12265 18343
rect 12299 18340 12311 18343
rect 18138 18340 18144 18352
rect 12299 18312 18144 18340
rect 12299 18309 12311 18312
rect 12253 18303 12311 18309
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 18248 18312 21128 18340
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 10689 18275 10747 18281
rect 10689 18241 10701 18275
rect 10735 18272 10747 18275
rect 11054 18272 11060 18284
rect 10735 18244 11060 18272
rect 10735 18241 10747 18244
rect 10689 18235 10747 18241
rect 11054 18232 11060 18244
rect 11112 18272 11118 18284
rect 11609 18275 11667 18281
rect 11609 18272 11621 18275
rect 11112 18244 11621 18272
rect 11112 18232 11118 18244
rect 11609 18241 11621 18244
rect 11655 18241 11667 18275
rect 11609 18235 11667 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13814 18272 13820 18284
rect 13219 18244 13820 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14182 18272 14188 18284
rect 14143 18244 14188 18272
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 16666 18232 16672 18284
rect 16724 18272 16730 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16724 18244 16865 18272
rect 16724 18232 16730 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17770 18232 17776 18284
rect 17828 18272 17834 18284
rect 18248 18272 18276 18312
rect 17828 18244 18276 18272
rect 17828 18232 17834 18244
rect 18322 18232 18328 18284
rect 18380 18272 18386 18284
rect 18877 18275 18935 18281
rect 18877 18272 18889 18275
rect 18380 18244 18889 18272
rect 18380 18232 18386 18244
rect 18877 18241 18889 18244
rect 18923 18241 18935 18275
rect 19058 18272 19064 18284
rect 19019 18244 19064 18272
rect 18877 18235 18935 18241
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 19794 18272 19800 18284
rect 19755 18244 19800 18272
rect 19794 18232 19800 18244
rect 19852 18232 19858 18284
rect 20622 18272 20628 18284
rect 20583 18244 20628 18272
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 14553 18207 14611 18213
rect 14553 18204 14565 18207
rect 8864 18176 14565 18204
rect 14553 18173 14565 18176
rect 14599 18173 14611 18207
rect 17954 18204 17960 18216
rect 14553 18167 14611 18173
rect 16132 18176 17960 18204
rect 4154 18145 4160 18148
rect 2924 18108 4108 18136
rect 2924 18096 2930 18108
rect 4148 18099 4160 18145
rect 4212 18136 4218 18148
rect 4212 18108 4248 18136
rect 4154 18096 4160 18099
rect 4212 18096 4218 18108
rect 4430 18096 4436 18148
rect 4488 18136 4494 18148
rect 5997 18139 6055 18145
rect 5997 18136 6009 18139
rect 4488 18108 6009 18136
rect 4488 18096 4494 18108
rect 5997 18105 6009 18108
rect 6043 18105 6055 18139
rect 5997 18099 6055 18105
rect 7466 18096 7472 18148
rect 7524 18136 7530 18148
rect 8478 18136 8484 18148
rect 7524 18108 8484 18136
rect 7524 18096 7530 18108
rect 8478 18096 8484 18108
rect 8536 18096 8542 18148
rect 9401 18139 9459 18145
rect 9401 18105 9413 18139
rect 9447 18136 9459 18139
rect 11330 18136 11336 18148
rect 9447 18108 11336 18136
rect 9447 18105 9459 18108
rect 9401 18099 9459 18105
rect 11330 18096 11336 18108
rect 11388 18096 11394 18148
rect 11425 18139 11483 18145
rect 11425 18105 11437 18139
rect 11471 18136 11483 18139
rect 11698 18136 11704 18148
rect 11471 18108 11704 18136
rect 11471 18105 11483 18108
rect 11425 18099 11483 18105
rect 11698 18096 11704 18108
rect 11756 18096 11762 18148
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 12989 18139 13047 18145
rect 12989 18136 13001 18139
rect 12676 18108 13001 18136
rect 12676 18096 12682 18108
rect 12989 18105 13001 18108
rect 13035 18105 13047 18139
rect 12989 18099 13047 18105
rect 13814 18096 13820 18148
rect 13872 18136 13878 18148
rect 15105 18139 15163 18145
rect 15105 18136 15117 18139
rect 13872 18108 15117 18136
rect 13872 18096 13878 18108
rect 15105 18105 15117 18108
rect 15151 18105 15163 18139
rect 15105 18099 15163 18105
rect 3234 18068 3240 18080
rect 3195 18040 3240 18068
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5905 18071 5963 18077
rect 5905 18068 5917 18071
rect 5592 18040 5917 18068
rect 5592 18028 5598 18040
rect 5905 18037 5917 18040
rect 5951 18037 5963 18071
rect 5905 18031 5963 18037
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 7064 18040 7297 18068
rect 7064 18028 7070 18040
rect 7285 18037 7297 18040
rect 7331 18068 7343 18071
rect 7653 18071 7711 18077
rect 7653 18068 7665 18071
rect 7331 18040 7665 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 7653 18037 7665 18040
rect 7699 18037 7711 18071
rect 8386 18068 8392 18080
rect 8347 18040 8392 18068
rect 7653 18031 7711 18037
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 9493 18071 9551 18077
rect 9493 18037 9505 18071
rect 9539 18068 9551 18071
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9539 18040 10057 18068
rect 9539 18037 9551 18040
rect 9493 18031 9551 18037
rect 10045 18037 10057 18040
rect 10091 18037 10103 18071
rect 10410 18068 10416 18080
rect 10371 18040 10416 18068
rect 10045 18031 10103 18037
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10560 18040 10605 18068
rect 10560 18028 10566 18040
rect 10686 18028 10692 18080
rect 10744 18068 10750 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 10744 18040 11529 18068
rect 10744 18028 10750 18040
rect 11517 18037 11529 18040
rect 11563 18068 11575 18071
rect 12253 18071 12311 18077
rect 12253 18068 12265 18071
rect 11563 18040 12265 18068
rect 11563 18037 11575 18040
rect 11517 18031 11575 18037
rect 12253 18037 12265 18040
rect 12299 18037 12311 18071
rect 12253 18031 12311 18037
rect 12897 18071 12955 18077
rect 12897 18037 12909 18071
rect 12943 18068 12955 18071
rect 13354 18068 13360 18080
rect 12943 18040 13360 18068
rect 12943 18037 12955 18040
rect 12897 18031 12955 18037
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 16132 18068 16160 18176
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18690 18164 18696 18216
rect 18748 18204 18754 18216
rect 18785 18207 18843 18213
rect 18785 18204 18797 18207
rect 18748 18176 18797 18204
rect 18748 18164 18754 18176
rect 18785 18173 18797 18176
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 21100 18213 21128 18312
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 19392 18176 19625 18204
rect 19392 18164 19398 18176
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19613 18167 19671 18173
rect 20349 18207 20407 18213
rect 20349 18173 20361 18207
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 21085 18207 21143 18213
rect 21085 18173 21097 18207
rect 21131 18173 21143 18207
rect 21085 18167 21143 18173
rect 16669 18139 16727 18145
rect 16669 18105 16681 18139
rect 16715 18136 16727 18139
rect 18138 18136 18144 18148
rect 16715 18108 18144 18136
rect 16715 18105 16727 18108
rect 16669 18099 16727 18105
rect 18138 18096 18144 18108
rect 18196 18096 18202 18148
rect 19242 18096 19248 18148
rect 19300 18136 19306 18148
rect 20364 18136 20392 18167
rect 19300 18108 20392 18136
rect 19300 18096 19306 18108
rect 13955 18040 16160 18068
rect 16301 18071 16359 18077
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 16574 18068 16580 18080
rect 16347 18040 16580 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 18417 18071 18475 18077
rect 16816 18040 16861 18068
rect 16816 18028 16822 18040
rect 18417 18037 18429 18071
rect 18463 18068 18475 18071
rect 19058 18068 19064 18080
rect 18463 18040 19064 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 19794 18028 19800 18080
rect 19852 18068 19858 18080
rect 20070 18068 20076 18080
rect 19852 18040 20076 18068
rect 19852 18028 19858 18040
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 3234 17864 3240 17876
rect 3007 17836 3240 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 3234 17824 3240 17836
rect 3292 17824 3298 17876
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 3476 17836 4292 17864
rect 3476 17824 3482 17836
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2225 17799 2283 17805
rect 2225 17796 2237 17799
rect 1820 17768 2237 17796
rect 1820 17756 1826 17768
rect 2225 17765 2237 17768
rect 2271 17765 2283 17799
rect 4264 17796 4292 17836
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4396 17836 4537 17864
rect 4396 17824 4402 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 4525 17827 4583 17833
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7469 17867 7527 17873
rect 7469 17864 7481 17867
rect 7432 17836 7481 17864
rect 7432 17824 7438 17836
rect 7469 17833 7481 17836
rect 7515 17833 7527 17867
rect 7469 17827 7527 17833
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7800 17836 7849 17864
rect 7800 17824 7806 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 11057 17867 11115 17873
rect 11057 17833 11069 17867
rect 11103 17864 11115 17867
rect 11146 17864 11152 17876
rect 11103 17836 11152 17864
rect 11103 17833 11115 17836
rect 11057 17827 11115 17833
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11330 17864 11336 17876
rect 11291 17836 11336 17864
rect 11330 17824 11336 17836
rect 11388 17824 11394 17876
rect 11701 17867 11759 17873
rect 11701 17833 11713 17867
rect 11747 17864 11759 17867
rect 11882 17864 11888 17876
rect 11747 17836 11888 17864
rect 11747 17833 11759 17836
rect 11701 17827 11759 17833
rect 11882 17824 11888 17836
rect 11940 17824 11946 17876
rect 12437 17867 12495 17873
rect 12437 17833 12449 17867
rect 12483 17864 12495 17867
rect 12618 17864 12624 17876
rect 12483 17836 12624 17864
rect 12483 17833 12495 17836
rect 12437 17827 12495 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 13449 17867 13507 17873
rect 13449 17864 13461 17867
rect 13412 17836 13461 17864
rect 13412 17824 13418 17836
rect 13449 17833 13461 17836
rect 13495 17833 13507 17867
rect 13814 17864 13820 17876
rect 13775 17836 13820 17864
rect 13449 17827 13507 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 16301 17867 16359 17873
rect 16301 17833 16313 17867
rect 16347 17864 16359 17867
rect 16758 17864 16764 17876
rect 16347 17836 16764 17864
rect 16347 17833 16359 17836
rect 16301 17827 16359 17833
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 17865 17867 17923 17873
rect 17865 17833 17877 17867
rect 17911 17864 17923 17867
rect 20254 17864 20260 17876
rect 17911 17836 20260 17864
rect 17911 17833 17923 17836
rect 17865 17827 17923 17833
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 21082 17864 21088 17876
rect 21043 17836 21088 17864
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 22002 17864 22008 17876
rect 21963 17836 22008 17864
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 4433 17799 4491 17805
rect 4264 17768 4384 17796
rect 2225 17759 2283 17765
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1938 17731 1996 17737
rect 1938 17728 1950 17731
rect 1397 17691 1455 17697
rect 1872 17700 1950 17728
rect 1412 17524 1440 17691
rect 1872 17660 1900 17700
rect 1938 17697 1950 17700
rect 1984 17697 1996 17731
rect 1938 17691 1996 17697
rect 2130 17688 2136 17740
rect 2188 17728 2194 17740
rect 3329 17731 3387 17737
rect 3329 17728 3341 17731
rect 2188 17700 3341 17728
rect 2188 17688 2194 17700
rect 3329 17697 3341 17700
rect 3375 17697 3387 17731
rect 4356 17728 4384 17768
rect 4433 17765 4445 17799
rect 4479 17796 4491 17799
rect 4798 17796 4804 17808
rect 4479 17768 4804 17796
rect 4479 17765 4491 17768
rect 4433 17759 4491 17765
rect 4798 17756 4804 17768
rect 4856 17756 4862 17808
rect 5626 17805 5632 17808
rect 5620 17796 5632 17805
rect 5587 17768 5632 17796
rect 5620 17759 5632 17768
rect 5626 17756 5632 17759
rect 5684 17756 5690 17808
rect 5718 17756 5724 17808
rect 5776 17796 5782 17808
rect 10502 17796 10508 17808
rect 5776 17768 10508 17796
rect 5776 17756 5782 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 12897 17799 12955 17805
rect 11072 17768 11836 17796
rect 11072 17740 11100 17768
rect 8662 17728 8668 17740
rect 4356 17700 8668 17728
rect 3329 17691 3387 17697
rect 8662 17688 8668 17700
rect 8720 17688 8726 17740
rect 8846 17728 8852 17740
rect 8807 17700 8852 17728
rect 8846 17688 8852 17700
rect 8904 17688 8910 17740
rect 8941 17731 8999 17737
rect 8941 17697 8953 17731
rect 8987 17728 8999 17731
rect 9214 17728 9220 17740
rect 8987 17700 9220 17728
rect 8987 17697 8999 17700
rect 8941 17691 8999 17697
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9933 17731 9991 17737
rect 9933 17728 9945 17731
rect 9456 17700 9945 17728
rect 9456 17688 9462 17700
rect 9933 17697 9945 17700
rect 9979 17728 9991 17731
rect 11054 17728 11060 17740
rect 9979 17700 11060 17728
rect 9979 17697 9991 17700
rect 9933 17691 9991 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 11808 17728 11836 17768
rect 12897 17765 12909 17799
rect 12943 17796 12955 17799
rect 13170 17796 13176 17808
rect 12943 17768 13176 17796
rect 12943 17765 12955 17768
rect 12897 17759 12955 17765
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 16574 17756 16580 17808
rect 16632 17796 16638 17808
rect 17957 17799 18015 17805
rect 17957 17796 17969 17799
rect 16632 17768 17969 17796
rect 16632 17756 16638 17768
rect 17957 17765 17969 17768
rect 18003 17765 18015 17799
rect 17957 17759 18015 17765
rect 18969 17799 19027 17805
rect 18969 17765 18981 17799
rect 19015 17796 19027 17799
rect 19242 17796 19248 17808
rect 19015 17768 19248 17796
rect 19015 17765 19027 17768
rect 18969 17759 19027 17765
rect 19242 17756 19248 17768
rect 19300 17756 19306 17808
rect 20070 17796 20076 17808
rect 19352 17768 20076 17796
rect 12805 17731 12863 17737
rect 11808 17700 11928 17728
rect 2222 17660 2228 17672
rect 1872 17632 2228 17660
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 3510 17660 3516 17672
rect 3471 17632 3516 17660
rect 3510 17620 3516 17632
rect 3568 17620 3574 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 4212 17632 4629 17660
rect 4212 17620 4218 17632
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 5350 17660 5356 17672
rect 5311 17632 5356 17660
rect 4617 17623 4675 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7524 17632 7941 17660
rect 7524 17620 7530 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 9122 17660 9128 17672
rect 8159 17632 8800 17660
rect 9083 17632 9128 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 1762 17552 1768 17604
rect 1820 17592 1826 17604
rect 3694 17592 3700 17604
rect 1820 17564 3700 17592
rect 1820 17552 1826 17564
rect 3694 17552 3700 17564
rect 3752 17552 3758 17604
rect 4065 17595 4123 17601
rect 4065 17561 4077 17595
rect 4111 17592 4123 17595
rect 4430 17592 4436 17604
rect 4111 17564 4436 17592
rect 4111 17561 4123 17564
rect 4065 17555 4123 17561
rect 4430 17552 4436 17564
rect 4488 17552 4494 17604
rect 8772 17592 8800 17632
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 9677 17663 9735 17669
rect 9677 17660 9689 17663
rect 9548 17632 9689 17660
rect 9548 17620 9554 17632
rect 9677 17629 9689 17632
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 10686 17620 10692 17672
rect 10744 17660 10750 17672
rect 11900 17669 11928 17700
rect 12805 17697 12817 17731
rect 12851 17728 12863 17731
rect 13630 17728 13636 17740
rect 12851 17700 13636 17728
rect 12851 17697 12863 17700
rect 12805 17691 12863 17697
rect 13630 17688 13636 17700
rect 13688 17688 13694 17740
rect 14090 17688 14096 17740
rect 14148 17728 14154 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 14148 17700 15669 17728
rect 14148 17688 14154 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17728 15807 17731
rect 16669 17731 16727 17737
rect 15795 17700 16344 17728
rect 15795 17697 15807 17700
rect 15749 17691 15807 17697
rect 16316 17672 16344 17700
rect 16669 17697 16681 17731
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 16761 17731 16819 17737
rect 16761 17697 16773 17731
rect 16807 17728 16819 17731
rect 17310 17728 17316 17740
rect 16807 17700 17316 17728
rect 16807 17697 16819 17700
rect 16761 17691 16819 17697
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 10744 17632 11805 17660
rect 10744 17620 10750 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11885 17663 11943 17669
rect 11885 17629 11897 17663
rect 11931 17629 11943 17663
rect 11885 17623 11943 17629
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 13081 17663 13139 17669
rect 13081 17660 13093 17663
rect 12584 17632 13093 17660
rect 12584 17620 12590 17632
rect 13081 17629 13093 17632
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 9306 17592 9312 17604
rect 6656 17564 8616 17592
rect 8772 17564 9312 17592
rect 6656 17524 6684 17564
rect 1412 17496 6684 17524
rect 6733 17527 6791 17533
rect 6733 17493 6745 17527
rect 6779 17524 6791 17527
rect 6822 17524 6828 17536
rect 6779 17496 6828 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 8294 17484 8300 17536
rect 8352 17524 8358 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8352 17496 8493 17524
rect 8352 17484 8358 17496
rect 8481 17493 8493 17496
rect 8527 17493 8539 17527
rect 8588 17524 8616 17564
rect 9306 17552 9312 17564
rect 9364 17552 9370 17604
rect 13096 17592 13124 17623
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 13909 17663 13967 17669
rect 13909 17660 13921 17663
rect 13872 17632 13921 17660
rect 13872 17620 13878 17632
rect 13909 17629 13921 17632
rect 13955 17629 13967 17663
rect 13909 17623 13967 17629
rect 14001 17663 14059 17669
rect 14001 17629 14013 17663
rect 14047 17629 14059 17663
rect 14001 17623 14059 17629
rect 14016 17592 14044 17623
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 15896 17632 15941 17660
rect 15896 17620 15902 17632
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 16684 17660 16712 17691
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 18877 17731 18935 17737
rect 18877 17728 18889 17731
rect 17420 17700 18889 17728
rect 16632 17632 16712 17660
rect 16945 17663 17003 17669
rect 16632 17620 16638 17632
rect 16945 17629 16957 17663
rect 16991 17660 17003 17663
rect 17126 17660 17132 17672
rect 16991 17632 17132 17660
rect 16991 17629 17003 17632
rect 16945 17623 17003 17629
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 17420 17660 17448 17700
rect 18877 17697 18889 17700
rect 18923 17697 18935 17731
rect 18877 17691 18935 17697
rect 17276 17632 17448 17660
rect 17276 17620 17282 17632
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 18049 17663 18107 17669
rect 18049 17660 18061 17663
rect 17736 17632 18061 17660
rect 17736 17620 17742 17632
rect 18049 17629 18061 17632
rect 18095 17629 18107 17663
rect 18049 17623 18107 17629
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 19061 17663 19119 17669
rect 19061 17660 19073 17663
rect 18748 17632 19073 17660
rect 18748 17620 18754 17632
rect 19061 17629 19073 17632
rect 19107 17629 19119 17663
rect 19061 17623 19119 17629
rect 19150 17620 19156 17672
rect 19208 17660 19214 17672
rect 19352 17660 19380 17768
rect 20070 17756 20076 17768
rect 20128 17756 20134 17808
rect 20165 17799 20223 17805
rect 20165 17765 20177 17799
rect 20211 17796 20223 17799
rect 21634 17796 21640 17808
rect 20211 17768 21640 17796
rect 20211 17765 20223 17768
rect 20165 17759 20223 17765
rect 21634 17756 21640 17768
rect 21692 17756 21698 17808
rect 20898 17728 20904 17740
rect 20859 17700 20904 17728
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 20162 17660 20168 17672
rect 19208 17632 19380 17660
rect 19444 17632 20168 17660
rect 19208 17620 19214 17632
rect 13096 17564 14044 17592
rect 15289 17595 15347 17601
rect 15289 17561 15301 17595
rect 15335 17592 15347 17595
rect 18414 17592 18420 17604
rect 15335 17564 18420 17592
rect 15335 17561 15347 17564
rect 15289 17555 15347 17561
rect 18414 17552 18420 17564
rect 18472 17552 18478 17604
rect 18509 17595 18567 17601
rect 18509 17561 18521 17595
rect 18555 17592 18567 17595
rect 18555 17564 19288 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 11054 17524 11060 17536
rect 8588 17496 11060 17524
rect 8481 17487 8539 17493
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 17402 17524 17408 17536
rect 11204 17496 17408 17524
rect 11204 17484 11210 17496
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 17497 17527 17555 17533
rect 17497 17493 17509 17527
rect 17543 17524 17555 17527
rect 18874 17524 18880 17536
rect 17543 17496 18880 17524
rect 17543 17493 17555 17496
rect 17497 17487 17555 17493
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 19260 17524 19288 17564
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19444 17592 19472 17632
rect 20162 17620 20168 17632
rect 20220 17660 20226 17672
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 20220 17632 20269 17660
rect 20220 17620 20226 17632
rect 20257 17629 20269 17632
rect 20303 17629 20315 17663
rect 20257 17623 20315 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17660 20499 17663
rect 20530 17660 20536 17672
rect 20487 17632 20536 17660
rect 20487 17629 20499 17632
rect 20441 17623 20499 17629
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 21818 17592 21824 17604
rect 19392 17564 19472 17592
rect 19536 17564 21824 17592
rect 19392 17552 19398 17564
rect 19536 17524 19564 17564
rect 21818 17552 21824 17564
rect 21876 17552 21882 17604
rect 19260 17496 19564 17524
rect 19610 17484 19616 17536
rect 19668 17524 19674 17536
rect 19797 17527 19855 17533
rect 19797 17524 19809 17527
rect 19668 17496 19809 17524
rect 19668 17484 19674 17496
rect 19797 17493 19809 17496
rect 19843 17493 19855 17527
rect 19797 17487 19855 17493
rect 20162 17484 20168 17536
rect 20220 17524 20226 17536
rect 20438 17524 20444 17536
rect 20220 17496 20444 17524
rect 20220 17484 20226 17496
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1486 17280 1492 17332
rect 1544 17320 1550 17332
rect 1949 17323 2007 17329
rect 1949 17320 1961 17323
rect 1544 17292 1961 17320
rect 1544 17280 1550 17292
rect 1949 17289 1961 17292
rect 1995 17289 2007 17323
rect 3050 17320 3056 17332
rect 1949 17283 2007 17289
rect 2792 17292 3056 17320
rect 2792 17193 2820 17292
rect 3050 17280 3056 17292
rect 3108 17320 3114 17332
rect 3878 17320 3884 17332
rect 3108 17292 3884 17320
rect 3108 17280 3114 17292
rect 3878 17280 3884 17292
rect 3936 17280 3942 17332
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17320 4218 17332
rect 4341 17323 4399 17329
rect 4341 17320 4353 17323
rect 4212 17292 4353 17320
rect 4212 17280 4218 17292
rect 4341 17289 4353 17292
rect 4387 17289 4399 17323
rect 4341 17283 4399 17289
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 5534 17320 5540 17332
rect 4479 17292 5540 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5718 17320 5724 17332
rect 5679 17292 5724 17320
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 7009 17323 7067 17329
rect 7009 17289 7021 17323
rect 7055 17320 7067 17323
rect 9398 17320 9404 17332
rect 7055 17292 9076 17320
rect 9359 17292 9404 17320
rect 7055 17289 7067 17292
rect 7009 17283 7067 17289
rect 3804 17224 6500 17252
rect 3804 17196 3832 17224
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4985 17187 5043 17193
rect 4985 17184 4997 17187
rect 4387 17156 4997 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 4985 17153 4997 17156
rect 5031 17153 5043 17187
rect 4985 17147 5043 17153
rect 5166 17144 5172 17196
rect 5224 17184 5230 17196
rect 6181 17187 6239 17193
rect 6181 17184 6193 17187
rect 5224 17156 6193 17184
rect 5224 17144 5230 17156
rect 6181 17153 6193 17156
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17153 6423 17187
rect 6472 17184 6500 17224
rect 7374 17184 7380 17196
rect 6472 17156 7380 17184
rect 6365 17147 6423 17153
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 3044 17119 3102 17125
rect 3044 17085 3056 17119
rect 3090 17116 3102 17119
rect 3602 17116 3608 17128
rect 3090 17088 3608 17116
rect 3090 17085 3102 17088
rect 3044 17079 3102 17085
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 6380 17116 6408 17147
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 7558 17184 7564 17196
rect 7519 17156 7564 17184
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7708 17156 8033 17184
rect 7708 17144 7714 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 9048 17184 9076 17292
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 10686 17320 10692 17332
rect 10647 17292 10692 17320
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 11054 17280 11060 17332
rect 11112 17320 11118 17332
rect 12250 17320 12256 17332
rect 11112 17292 12256 17320
rect 11112 17280 11118 17292
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12351 17292 15139 17320
rect 9214 17212 9220 17264
rect 9272 17252 9278 17264
rect 12158 17252 12164 17264
rect 9272 17224 12164 17252
rect 9272 17212 9278 17224
rect 12158 17212 12164 17224
rect 12216 17212 12222 17264
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 9048 17156 10149 17184
rect 8021 17147 8079 17153
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 11422 17184 11428 17196
rect 11379 17156 11428 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 6822 17116 6828 17128
rect 6380 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17116 6886 17128
rect 6880 17088 7972 17116
rect 6880 17076 6886 17088
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 5166 17048 5172 17060
rect 3200 17020 5172 17048
rect 3200 17008 3206 17020
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 5258 17008 5264 17060
rect 5316 17048 5322 17060
rect 6089 17051 6147 17057
rect 6089 17048 6101 17051
rect 5316 17020 6101 17048
rect 5316 17008 5322 17020
rect 6089 17017 6101 17020
rect 6135 17048 6147 17051
rect 6638 17048 6644 17060
rect 6135 17020 6644 17048
rect 6135 17017 6147 17020
rect 6089 17011 6147 17017
rect 6638 17008 6644 17020
rect 6696 17008 6702 17060
rect 6914 17008 6920 17060
rect 6972 17048 6978 17060
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 6972 17020 7481 17048
rect 6972 17008 6978 17020
rect 7469 17017 7481 17020
rect 7515 17017 7527 17051
rect 7944 17048 7972 17088
rect 8570 17076 8576 17128
rect 8628 17116 8634 17128
rect 10244 17116 10272 17147
rect 11054 17116 11060 17128
rect 8628 17088 10272 17116
rect 11015 17088 11060 17116
rect 8628 17076 8634 17088
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 8288 17051 8346 17057
rect 8288 17048 8300 17051
rect 7944 17020 8300 17048
rect 7469 17011 7527 17017
rect 8288 17017 8300 17020
rect 8334 17048 8346 17051
rect 11348 17048 11376 17147
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 12351 17184 12379 17292
rect 15111 17252 15139 17292
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15528 17292 15577 17320
rect 15528 17280 15534 17292
rect 15565 17289 15577 17292
rect 15611 17320 15623 17323
rect 15838 17320 15844 17332
rect 15611 17292 15844 17320
rect 15611 17289 15623 17292
rect 15565 17283 15623 17289
rect 15838 17280 15844 17292
rect 15896 17280 15902 17332
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 16853 17323 16911 17329
rect 16853 17320 16865 17323
rect 16632 17292 16865 17320
rect 16632 17280 16638 17292
rect 16853 17289 16865 17292
rect 16899 17289 16911 17323
rect 16853 17283 16911 17289
rect 18417 17323 18475 17329
rect 18417 17289 18429 17323
rect 18463 17320 18475 17323
rect 18782 17320 18788 17332
rect 18463 17292 18788 17320
rect 18463 17289 18475 17292
rect 18417 17283 18475 17289
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 19702 17320 19708 17332
rect 19076 17292 19708 17320
rect 17586 17252 17592 17264
rect 15111 17224 17356 17252
rect 11848 17156 12379 17184
rect 11848 17144 11854 17156
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 16390 17184 16396 17196
rect 15712 17156 16396 17184
rect 15712 17144 15718 17156
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 17328 17193 17356 17224
rect 17420 17224 17592 17252
rect 17420 17193 17448 17224
rect 17586 17212 17592 17224
rect 17644 17212 17650 17264
rect 19076 17252 19104 17292
rect 19702 17280 19708 17292
rect 19760 17280 19766 17332
rect 18892 17224 19104 17252
rect 18892 17193 18920 17224
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 20622 17252 20628 17264
rect 19208 17224 20628 17252
rect 19208 17212 19214 17224
rect 20622 17212 20628 17224
rect 20680 17212 20686 17264
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17405 17187 17463 17193
rect 17405 17153 17417 17187
rect 17451 17153 17463 17187
rect 18877 17187 18935 17193
rect 18877 17184 18889 17187
rect 17405 17147 17463 17153
rect 17512 17156 18889 17184
rect 12342 17076 12348 17128
rect 12400 17116 12406 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12400 17088 12449 17116
rect 12400 17076 12406 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12704 17119 12762 17125
rect 12704 17085 12716 17119
rect 12750 17116 12762 17119
rect 13538 17116 13544 17128
rect 12750 17088 13544 17116
rect 12750 17085 12762 17088
rect 12704 17079 12762 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 14185 17119 14243 17125
rect 14185 17116 14197 17119
rect 13872 17088 14197 17116
rect 13872 17076 13878 17088
rect 14185 17085 14197 17088
rect 14231 17085 14243 17119
rect 16209 17119 16267 17125
rect 16209 17116 16221 17119
rect 14185 17079 14243 17085
rect 14292 17088 16221 17116
rect 8334 17020 11376 17048
rect 8334 17017 8346 17020
rect 8288 17011 8346 17017
rect 12802 17008 12808 17060
rect 12860 17048 12866 17060
rect 14292 17048 14320 17088
rect 16209 17085 16221 17088
rect 16255 17085 16267 17119
rect 16209 17079 16267 17085
rect 16942 17076 16948 17128
rect 17000 17116 17006 17128
rect 17512 17116 17540 17156
rect 18877 17153 18889 17156
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17184 19395 17187
rect 19889 17187 19947 17193
rect 19889 17184 19901 17187
rect 19383 17156 19901 17184
rect 19383 17153 19395 17156
rect 19337 17147 19395 17153
rect 19889 17153 19901 17156
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20530 17184 20536 17196
rect 20027 17156 20536 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 17000 17088 17540 17116
rect 17000 17076 17006 17088
rect 18598 17076 18604 17128
rect 18656 17116 18662 17128
rect 18984 17116 19012 17147
rect 18656 17088 19012 17116
rect 18656 17076 18662 17088
rect 19150 17076 19156 17128
rect 19208 17116 19214 17128
rect 19996 17116 20024 17147
rect 20530 17144 20536 17156
rect 20588 17184 20594 17196
rect 20993 17187 21051 17193
rect 20993 17184 21005 17187
rect 20588 17156 21005 17184
rect 20588 17144 20594 17156
rect 20993 17153 21005 17156
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 19208 17088 20024 17116
rect 19208 17076 19214 17088
rect 20070 17076 20076 17128
rect 20128 17116 20134 17128
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 20128 17088 20913 17116
rect 20128 17076 20134 17088
rect 20901 17085 20913 17088
rect 20947 17085 20959 17119
rect 20901 17079 20959 17085
rect 12860 17020 14320 17048
rect 14452 17051 14510 17057
rect 12860 17008 12866 17020
rect 14452 17017 14464 17051
rect 14498 17048 14510 17051
rect 14734 17048 14740 17060
rect 14498 17020 14740 17048
rect 14498 17017 14510 17020
rect 14452 17011 14510 17017
rect 14734 17008 14740 17020
rect 14792 17008 14798 17060
rect 16301 17051 16359 17057
rect 16301 17048 16313 17051
rect 14844 17020 16313 17048
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 4801 16983 4859 16989
rect 4801 16980 4813 16983
rect 3016 16952 4813 16980
rect 3016 16940 3022 16952
rect 4801 16949 4813 16952
rect 4847 16949 4859 16983
rect 4801 16943 4859 16949
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 7374 16980 7380 16992
rect 4948 16952 4993 16980
rect 7335 16952 7380 16980
rect 4948 16940 4954 16952
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 9674 16980 9680 16992
rect 9635 16952 9680 16980
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 10042 16980 10048 16992
rect 10003 16952 10048 16980
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 11330 16940 11336 16992
rect 11388 16980 11394 16992
rect 11882 16980 11888 16992
rect 11388 16952 11888 16980
rect 11388 16940 11394 16952
rect 11882 16940 11888 16952
rect 11940 16980 11946 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 11940 16952 13829 16980
rect 11940 16940 11946 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 13906 16940 13912 16992
rect 13964 16980 13970 16992
rect 14844 16980 14872 17020
rect 16301 17017 16313 17020
rect 16347 17017 16359 17051
rect 16301 17011 16359 17017
rect 17221 17051 17279 17057
rect 17221 17017 17233 17051
rect 17267 17048 17279 17051
rect 17494 17048 17500 17060
rect 17267 17020 17500 17048
rect 17267 17017 17279 17020
rect 17221 17011 17279 17017
rect 17494 17008 17500 17020
rect 17552 17008 17558 17060
rect 18046 17008 18052 17060
rect 18104 17048 18110 17060
rect 19337 17051 19395 17057
rect 19337 17048 19349 17051
rect 18104 17020 19349 17048
rect 18104 17008 18110 17020
rect 19337 17017 19349 17020
rect 19383 17017 19395 17051
rect 21910 17048 21916 17060
rect 19337 17011 19395 17017
rect 19444 17020 21916 17048
rect 13964 16952 14872 16980
rect 15841 16983 15899 16989
rect 13964 16940 13970 16952
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 16574 16980 16580 16992
rect 15887 16952 16580 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 17126 16940 17132 16992
rect 17184 16980 17190 16992
rect 17954 16980 17960 16992
rect 17184 16952 17960 16980
rect 17184 16940 17190 16952
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18782 16980 18788 16992
rect 18743 16952 18788 16980
rect 18782 16940 18788 16952
rect 18840 16940 18846 16992
rect 19444 16989 19472 17020
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 19429 16983 19487 16989
rect 19429 16949 19441 16983
rect 19475 16949 19487 16983
rect 19794 16980 19800 16992
rect 19755 16952 19800 16980
rect 19429 16943 19487 16949
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 20441 16983 20499 16989
rect 20441 16949 20453 16983
rect 20487 16980 20499 16983
rect 20530 16980 20536 16992
rect 20487 16952 20536 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 20806 16980 20812 16992
rect 20767 16952 20812 16980
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 2317 16779 2375 16785
rect 2317 16745 2329 16779
rect 2363 16776 2375 16779
rect 2498 16776 2504 16788
rect 2363 16748 2504 16776
rect 2363 16745 2375 16748
rect 2317 16739 2375 16745
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 2958 16776 2964 16788
rect 2919 16748 2964 16776
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 4890 16776 4896 16788
rect 4387 16748 4896 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 6638 16776 6644 16788
rect 6599 16748 6644 16776
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 9950 16776 9956 16788
rect 7432 16748 9956 16776
rect 7432 16736 7438 16748
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10410 16736 10416 16788
rect 10468 16776 10474 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 10468 16748 10885 16776
rect 10468 16736 10474 16748
rect 10873 16745 10885 16748
rect 10919 16745 10931 16779
rect 10873 16739 10931 16745
rect 11885 16779 11943 16785
rect 11885 16745 11897 16779
rect 11931 16745 11943 16779
rect 14274 16776 14280 16788
rect 11885 16739 11943 16745
rect 13280 16748 14280 16776
rect 198 16668 204 16720
rect 256 16708 262 16720
rect 2409 16711 2467 16717
rect 2409 16708 2421 16711
rect 256 16680 2421 16708
rect 256 16668 262 16680
rect 2409 16677 2421 16680
rect 2455 16708 2467 16711
rect 2866 16708 2872 16720
rect 2455 16680 2872 16708
rect 2455 16677 2467 16680
rect 2409 16671 2467 16677
rect 2866 16668 2872 16680
rect 2924 16668 2930 16720
rect 3234 16668 3240 16720
rect 3292 16708 3298 16720
rect 4801 16711 4859 16717
rect 4801 16708 4813 16711
rect 3292 16680 4813 16708
rect 3292 16668 3298 16680
rect 4801 16677 4813 16680
rect 4847 16677 4859 16711
rect 4801 16671 4859 16677
rect 5166 16668 5172 16720
rect 5224 16708 5230 16720
rect 6549 16711 6607 16717
rect 6549 16708 6561 16711
rect 5224 16680 6561 16708
rect 5224 16668 5230 16680
rect 6549 16677 6561 16680
rect 6595 16708 6607 16711
rect 8012 16711 8070 16717
rect 6595 16680 7880 16708
rect 6595 16677 6607 16680
rect 6549 16671 6607 16677
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16640 3387 16643
rect 4062 16640 4068 16652
rect 3375 16612 4068 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 4212 16612 4721 16640
rect 4212 16600 4218 16612
rect 4709 16609 4721 16612
rect 4755 16609 4767 16643
rect 4709 16603 4767 16609
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 5592 16612 6776 16640
rect 5592 16600 5598 16612
rect 2590 16572 2596 16584
rect 2551 16544 2596 16572
rect 2590 16532 2596 16544
rect 2648 16532 2654 16584
rect 3142 16532 3148 16584
rect 3200 16572 3206 16584
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 3200 16544 3433 16572
rect 3200 16532 3206 16544
rect 3421 16541 3433 16544
rect 3467 16541 3479 16575
rect 3602 16572 3608 16584
rect 3563 16544 3608 16572
rect 3421 16535 3479 16541
rect 3602 16532 3608 16544
rect 3660 16572 3666 16584
rect 4798 16572 4804 16584
rect 3660 16544 4804 16572
rect 3660 16532 3666 16544
rect 4798 16532 4804 16544
rect 4856 16572 4862 16584
rect 4893 16575 4951 16581
rect 4893 16572 4905 16575
rect 4856 16544 4905 16572
rect 4856 16532 4862 16544
rect 4893 16541 4905 16544
rect 4939 16541 4951 16575
rect 4893 16535 4951 16541
rect 4982 16532 4988 16584
rect 5040 16572 5046 16584
rect 5350 16572 5356 16584
rect 5040 16544 5356 16572
rect 5040 16532 5046 16544
rect 5350 16532 5356 16544
rect 5408 16572 5414 16584
rect 6748 16581 6776 16612
rect 7650 16600 7656 16652
rect 7708 16640 7714 16652
rect 7745 16643 7803 16649
rect 7745 16640 7757 16643
rect 7708 16612 7757 16640
rect 7708 16600 7714 16612
rect 7745 16609 7757 16612
rect 7791 16609 7803 16643
rect 7852 16640 7880 16680
rect 8012 16677 8024 16711
rect 8058 16708 8070 16711
rect 8570 16708 8576 16720
rect 8058 16680 8576 16708
rect 8058 16677 8070 16680
rect 8012 16671 8070 16677
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 8662 16668 8668 16720
rect 8720 16708 8726 16720
rect 10321 16711 10379 16717
rect 10321 16708 10333 16711
rect 8720 16680 10333 16708
rect 8720 16668 8726 16680
rect 10321 16677 10333 16680
rect 10367 16677 10379 16711
rect 11333 16711 11391 16717
rect 11333 16708 11345 16711
rect 10321 16671 10379 16677
rect 10419 16680 11345 16708
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 7852 16612 10241 16640
rect 7745 16603 7803 16609
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 6733 16575 6791 16581
rect 5408 16544 6408 16572
rect 5408 16532 5414 16544
rect 2314 16464 2320 16516
rect 2372 16504 2378 16516
rect 6380 16504 6408 16544
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 7098 16572 7104 16584
rect 6779 16544 7104 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 10419 16572 10447 16680
rect 11333 16677 11345 16680
rect 11379 16677 11391 16711
rect 11333 16671 11391 16677
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 11900 16640 11928 16739
rect 12253 16711 12311 16717
rect 12253 16677 12265 16711
rect 12299 16708 12311 16711
rect 12434 16708 12440 16720
rect 12299 16680 12440 16708
rect 12299 16677 12311 16680
rect 12253 16671 12311 16677
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 13280 16640 13308 16748
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 14608 16748 15301 16776
rect 14608 16736 14614 16748
rect 15289 16745 15301 16748
rect 15335 16745 15347 16779
rect 15289 16739 15347 16745
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 15657 16779 15715 16785
rect 15657 16776 15669 16779
rect 15620 16748 15669 16776
rect 15620 16736 15626 16748
rect 15657 16745 15669 16748
rect 15703 16745 15715 16779
rect 15657 16739 15715 16745
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 15838 16776 15844 16788
rect 15795 16748 15844 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 15838 16736 15844 16748
rect 15896 16776 15902 16788
rect 16022 16776 16028 16788
rect 15896 16748 16028 16776
rect 15896 16736 15902 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 16298 16776 16304 16788
rect 16259 16748 16304 16776
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 16761 16779 16819 16785
rect 16761 16776 16773 16779
rect 16632 16748 16773 16776
rect 16632 16736 16638 16748
rect 16761 16745 16773 16748
rect 16807 16745 16819 16779
rect 17310 16776 17316 16788
rect 17271 16748 17316 16776
rect 16761 16739 16819 16745
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17402 16736 17408 16788
rect 17460 16776 17466 16788
rect 17681 16779 17739 16785
rect 17681 16776 17693 16779
rect 17460 16748 17693 16776
rect 17460 16736 17466 16748
rect 17681 16745 17693 16748
rect 17727 16745 17739 16779
rect 17681 16739 17739 16745
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 18196 16748 18337 16776
rect 18196 16736 18202 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 18325 16739 18383 16745
rect 19337 16779 19395 16785
rect 19337 16745 19349 16779
rect 19383 16776 19395 16779
rect 20714 16776 20720 16788
rect 19383 16748 20720 16776
rect 19383 16745 19395 16748
rect 19337 16739 19395 16745
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 21085 16779 21143 16785
rect 21085 16745 21097 16779
rect 21131 16776 21143 16779
rect 22005 16779 22063 16785
rect 22005 16776 22017 16779
rect 21131 16748 22017 16776
rect 21131 16745 21143 16748
rect 21085 16739 21143 16745
rect 22005 16745 22017 16748
rect 22051 16745 22063 16779
rect 22005 16739 22063 16745
rect 13998 16668 14004 16720
rect 14056 16708 14062 16720
rect 17773 16711 17831 16717
rect 17773 16708 17785 16711
rect 14056 16680 17785 16708
rect 14056 16668 14062 16680
rect 17773 16677 17785 16680
rect 17819 16677 17831 16711
rect 17773 16671 17831 16677
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 18693 16711 18751 16717
rect 18693 16708 18705 16711
rect 17920 16680 18705 16708
rect 17920 16668 17926 16680
rect 18693 16677 18705 16680
rect 18739 16677 18751 16711
rect 18693 16671 18751 16677
rect 18785 16711 18843 16717
rect 18785 16677 18797 16711
rect 18831 16708 18843 16711
rect 19518 16708 19524 16720
rect 18831 16680 19524 16708
rect 18831 16677 18843 16680
rect 18785 16671 18843 16677
rect 19518 16668 19524 16680
rect 19576 16668 19582 16720
rect 19797 16711 19855 16717
rect 19797 16677 19809 16711
rect 19843 16708 19855 16711
rect 19978 16708 19984 16720
rect 19843 16680 19984 16708
rect 19843 16677 19855 16680
rect 19797 16671 19855 16677
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 11287 16612 11836 16640
rect 11900 16612 13308 16640
rect 13348 16643 13406 16649
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 9272 16544 10447 16572
rect 10505 16575 10563 16581
rect 9272 16532 9278 16544
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 10962 16572 10968 16584
rect 10551 16544 10968 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 10962 16532 10968 16544
rect 11020 16572 11026 16584
rect 11330 16572 11336 16584
rect 11020 16544 11336 16572
rect 11020 16532 11026 16544
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 11422 16532 11428 16584
rect 11480 16572 11486 16584
rect 11480 16544 11525 16572
rect 11480 16532 11486 16544
rect 7374 16504 7380 16516
rect 2372 16476 6316 16504
rect 6380 16476 7380 16504
rect 2372 16464 2378 16476
rect 1946 16436 1952 16448
rect 1907 16408 1952 16436
rect 1946 16396 1952 16408
rect 2004 16396 2010 16448
rect 2866 16396 2872 16448
rect 2924 16436 2930 16448
rect 4982 16436 4988 16448
rect 2924 16408 4988 16436
rect 2924 16396 2930 16408
rect 4982 16396 4988 16408
rect 5040 16396 5046 16448
rect 6178 16436 6184 16448
rect 6139 16408 6184 16436
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 6288 16436 6316 16476
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 11698 16504 11704 16516
rect 8680 16476 11704 16504
rect 8680 16436 8708 16476
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 6288 16408 8708 16436
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9306 16436 9312 16448
rect 9171 16408 9312 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9861 16439 9919 16445
rect 9861 16405 9873 16439
rect 9907 16436 9919 16439
rect 10686 16436 10692 16448
rect 9907 16408 10692 16436
rect 9907 16405 9919 16408
rect 9861 16399 9919 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 11808 16436 11836 16612
rect 13348 16609 13360 16643
rect 13394 16640 13406 16643
rect 13906 16640 13912 16652
rect 13394 16612 13912 16640
rect 13394 16609 13406 16612
rect 13348 16603 13406 16609
rect 13906 16600 13912 16612
rect 13964 16640 13970 16652
rect 14737 16643 14795 16649
rect 13964 16612 14688 16640
rect 13964 16600 13970 16612
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12124 16544 12357 16572
rect 12124 16532 12130 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 14660 16572 14688 16612
rect 14737 16609 14749 16643
rect 14783 16640 14795 16643
rect 16574 16640 16580 16652
rect 14783 16612 16580 16640
rect 14783 16609 14795 16612
rect 14737 16603 14795 16609
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 16669 16643 16727 16649
rect 16669 16609 16681 16643
rect 16715 16640 16727 16643
rect 16758 16640 16764 16652
rect 16715 16612 16764 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 17310 16600 17316 16652
rect 17368 16640 17374 16652
rect 19242 16640 19248 16652
rect 17368 16612 19248 16640
rect 17368 16600 17374 16612
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19705 16643 19763 16649
rect 19705 16640 19717 16643
rect 19484 16612 19717 16640
rect 19484 16600 19490 16612
rect 19705 16609 19717 16612
rect 19751 16609 19763 16643
rect 19705 16603 19763 16609
rect 20901 16643 20959 16649
rect 20901 16609 20913 16643
rect 20947 16640 20959 16643
rect 21174 16640 21180 16652
rect 20947 16612 21180 16640
rect 20947 16609 20959 16612
rect 20901 16603 20959 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 15654 16572 15660 16584
rect 14660 16544 15660 16572
rect 13081 16535 13139 16541
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 12452 16504 12480 16535
rect 12308 16476 12480 16504
rect 12308 16464 12314 16476
rect 12986 16436 12992 16448
rect 11808 16408 12992 16436
rect 12986 16396 12992 16408
rect 13044 16396 13050 16448
rect 13096 16436 13124 16535
rect 15654 16532 15660 16544
rect 15712 16572 15718 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15712 16544 15853 16572
rect 15712 16532 15718 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 15841 16535 15899 16541
rect 15948 16544 16865 16572
rect 14461 16507 14519 16513
rect 14461 16473 14473 16507
rect 14507 16504 14519 16507
rect 14734 16504 14740 16516
rect 14507 16476 14740 16504
rect 14507 16473 14519 16476
rect 14461 16467 14519 16473
rect 14734 16464 14740 16476
rect 14792 16504 14798 16516
rect 15948 16504 15976 16544
rect 16853 16541 16865 16544
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 17865 16575 17923 16581
rect 17865 16572 17877 16575
rect 17644 16544 17877 16572
rect 17644 16532 17650 16544
rect 17865 16541 17877 16544
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 17954 16532 17960 16584
rect 18012 16572 18018 16584
rect 18598 16572 18604 16584
rect 18012 16544 18604 16572
rect 18012 16532 18018 16544
rect 18598 16532 18604 16544
rect 18656 16572 18662 16584
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18656 16544 18889 16572
rect 18656 16532 18662 16544
rect 18877 16541 18889 16544
rect 18923 16572 18935 16575
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 18923 16544 19901 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 14792 16476 15976 16504
rect 14792 16464 14798 16476
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 19334 16504 19340 16516
rect 16080 16476 19340 16504
rect 16080 16464 16086 16476
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 13354 16436 13360 16448
rect 13096 16408 13360 16436
rect 13354 16396 13360 16408
rect 13412 16436 13418 16448
rect 13814 16436 13820 16448
rect 13412 16408 13820 16436
rect 13412 16396 13418 16408
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 14182 16396 14188 16448
rect 14240 16436 14246 16448
rect 15194 16436 15200 16448
rect 14240 16408 15200 16436
rect 14240 16396 14246 16408
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 16117 16439 16175 16445
rect 16117 16436 16129 16439
rect 15712 16408 16129 16436
rect 15712 16396 15718 16408
rect 16117 16405 16129 16408
rect 16163 16405 16175 16439
rect 16117 16399 16175 16405
rect 16482 16396 16488 16448
rect 16540 16436 16546 16448
rect 20806 16436 20812 16448
rect 16540 16408 20812 16436
rect 16540 16396 16546 16408
rect 20806 16396 20812 16408
rect 20864 16396 20870 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 3053 16235 3111 16241
rect 3053 16232 3065 16235
rect 1412 16204 3065 16232
rect 1412 16037 1440 16204
rect 3053 16201 3065 16204
rect 3099 16201 3111 16235
rect 4154 16232 4160 16244
rect 3053 16195 3111 16201
rect 3160 16204 4160 16232
rect 1486 16124 1492 16176
rect 1544 16164 1550 16176
rect 1581 16167 1639 16173
rect 1581 16164 1593 16167
rect 1544 16136 1593 16164
rect 1544 16124 1550 16136
rect 1581 16133 1593 16136
rect 1627 16133 1639 16167
rect 1581 16127 1639 16133
rect 2133 16167 2191 16173
rect 2133 16133 2145 16167
rect 2179 16164 2191 16167
rect 3160 16164 3188 16204
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4525 16235 4583 16241
rect 4525 16201 4537 16235
rect 4571 16232 4583 16235
rect 4798 16232 4804 16244
rect 4571 16204 4804 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 6822 16232 6828 16244
rect 5767 16204 6828 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 7650 16232 7656 16244
rect 6932 16204 7656 16232
rect 2179 16136 3188 16164
rect 2179 16133 2191 16136
rect 2133 16127 2191 16133
rect 6932 16108 6960 16204
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 8386 16192 8392 16244
rect 8444 16232 8450 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8444 16204 8769 16232
rect 8444 16192 8450 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 8938 16192 8944 16244
rect 8996 16232 9002 16244
rect 11146 16232 11152 16244
rect 8996 16204 11152 16232
rect 8996 16192 9002 16204
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 12710 16232 12716 16244
rect 11808 16204 12716 16232
rect 8297 16167 8355 16173
rect 8297 16133 8309 16167
rect 8343 16164 8355 16167
rect 8570 16164 8576 16176
rect 8343 16136 8576 16164
rect 8343 16133 8355 16136
rect 8297 16127 8355 16133
rect 8570 16124 8576 16136
rect 8628 16124 8634 16176
rect 9858 16124 9864 16176
rect 9916 16164 9922 16176
rect 11808 16164 11836 16204
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 13817 16235 13875 16241
rect 13817 16201 13829 16235
rect 13863 16232 13875 16235
rect 13906 16232 13912 16244
rect 13863 16204 13912 16232
rect 13863 16201 13875 16204
rect 13817 16195 13875 16201
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 14090 16232 14096 16244
rect 14051 16204 14096 16232
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 15120 16204 16865 16232
rect 9916 16136 11836 16164
rect 9916 16124 9922 16136
rect 11882 16124 11888 16176
rect 11940 16124 11946 16176
rect 2777 16099 2835 16105
rect 2777 16065 2789 16099
rect 2823 16096 2835 16099
rect 2823 16068 2912 16096
rect 2823 16065 2835 16068
rect 2777 16059 2835 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15960 2099 15963
rect 2593 15963 2651 15969
rect 2593 15960 2605 15963
rect 2087 15932 2605 15960
rect 2087 15929 2099 15932
rect 2041 15923 2099 15929
rect 2593 15929 2605 15932
rect 2639 15960 2651 15963
rect 2774 15960 2780 15972
rect 2639 15932 2780 15960
rect 2639 15929 2651 15932
rect 2593 15923 2651 15929
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 2884 15960 2912 16068
rect 2958 16056 2964 16108
rect 3016 16096 3022 16108
rect 6362 16096 6368 16108
rect 3016 16068 3280 16096
rect 6323 16068 6368 16096
rect 3016 16056 3022 16068
rect 3050 15988 3056 16040
rect 3108 16028 3114 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 3108 16000 3157 16028
rect 3108 15988 3114 16000
rect 3145 15997 3157 16000
rect 3191 15997 3203 16031
rect 3252 16028 3280 16068
rect 6362 16056 6368 16068
rect 6420 16056 6426 16108
rect 6914 16096 6920 16108
rect 6827 16068 6920 16096
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 9306 16096 9312 16108
rect 9267 16068 9312 16096
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 9640 16068 10333 16096
rect 9640 16056 9646 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 11425 16099 11483 16105
rect 10321 16059 10379 16065
rect 10980 16068 11284 16096
rect 5718 16028 5724 16040
rect 3252 16000 5724 16028
rect 3145 15991 3203 15997
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 6089 16031 6147 16037
rect 6089 15997 6101 16031
rect 6135 16028 6147 16031
rect 6178 16028 6184 16040
rect 6135 16000 6184 16028
rect 6135 15997 6147 16000
rect 6089 15991 6147 15997
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 7184 16031 7242 16037
rect 7184 15997 7196 16031
rect 7230 16028 7242 16031
rect 7558 16028 7564 16040
rect 7230 16000 7564 16028
rect 7230 15997 7242 16000
rect 7184 15991 7242 15997
rect 7558 15988 7564 16000
rect 7616 15988 7622 16040
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 7852 16000 9137 16028
rect 3412 15963 3470 15969
rect 3412 15960 3424 15963
rect 2884 15932 3424 15960
rect 3412 15929 3424 15932
rect 3458 15960 3470 15963
rect 3510 15960 3516 15972
rect 3458 15932 3516 15960
rect 3458 15929 3470 15932
rect 3412 15923 3470 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 6822 15960 6828 15972
rect 3620 15932 6828 15960
rect 2498 15892 2504 15904
rect 2459 15864 2504 15892
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 3053 15895 3111 15901
rect 3053 15861 3065 15895
rect 3099 15892 3111 15895
rect 3620 15892 3648 15932
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 4798 15892 4804 15904
rect 3099 15864 3648 15892
rect 4759 15864 4804 15892
rect 3099 15861 3111 15864
rect 3053 15855 3111 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 6181 15895 6239 15901
rect 6181 15892 6193 15895
rect 6052 15864 6193 15892
rect 6052 15852 6058 15864
rect 6181 15861 6193 15864
rect 6227 15861 6239 15895
rect 6181 15855 6239 15861
rect 6270 15852 6276 15904
rect 6328 15892 6334 15904
rect 7852 15892 7880 16000
rect 9125 15997 9137 16000
rect 9171 15997 9183 16031
rect 9125 15991 9183 15997
rect 9490 15988 9496 16040
rect 9548 16028 9554 16040
rect 10980 16028 11008 16068
rect 11146 16028 11152 16040
rect 9548 16000 11008 16028
rect 11107 16000 11152 16028
rect 9548 15988 9554 16000
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 11256 16028 11284 16068
rect 11425 16065 11437 16099
rect 11471 16096 11483 16099
rect 11900 16096 11928 16124
rect 14550 16096 14556 16108
rect 11471 16068 11928 16096
rect 14511 16068 14556 16096
rect 11471 16065 11483 16068
rect 11425 16059 11483 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 14734 16096 14740 16108
rect 14695 16068 14740 16096
rect 14734 16056 14740 16068
rect 14792 16056 14798 16108
rect 11256 16000 11468 16028
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 10137 15963 10195 15969
rect 7984 15932 9904 15960
rect 7984 15920 7990 15932
rect 8662 15892 8668 15904
rect 6328 15864 7880 15892
rect 8623 15864 8668 15892
rect 6328 15852 6334 15864
rect 8662 15852 8668 15864
rect 8720 15892 8726 15904
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 8720 15864 9229 15892
rect 8720 15852 8726 15864
rect 9217 15861 9229 15864
rect 9263 15861 9275 15895
rect 9766 15892 9772 15904
rect 9727 15864 9772 15892
rect 9217 15855 9275 15861
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 9876 15892 9904 15932
rect 10137 15929 10149 15963
rect 10183 15960 10195 15963
rect 10410 15960 10416 15972
rect 10183 15932 10416 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 10410 15920 10416 15932
rect 10468 15920 10474 15972
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 9876 15864 10241 15892
rect 10229 15861 10241 15864
rect 10275 15861 10287 15895
rect 10229 15855 10287 15861
rect 10594 15852 10600 15904
rect 10652 15892 10658 15904
rect 10781 15895 10839 15901
rect 10781 15892 10793 15895
rect 10652 15864 10793 15892
rect 10652 15852 10658 15864
rect 10781 15861 10793 15864
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11241 15895 11299 15901
rect 11241 15892 11253 15895
rect 11204 15864 11253 15892
rect 11204 15852 11210 15864
rect 11241 15861 11253 15864
rect 11287 15861 11299 15895
rect 11440 15892 11468 16000
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 12342 16028 12348 16040
rect 11572 16000 12348 16028
rect 11572 15988 11578 16000
rect 12342 15988 12348 16000
rect 12400 16028 12406 16040
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 12400 16000 12449 16028
rect 12400 15988 12406 16000
rect 12437 15997 12449 16000
rect 12483 16028 12495 16031
rect 14461 16031 14519 16037
rect 12483 16000 13400 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 13372 15972 13400 16000
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 15120 16028 15148 16204
rect 16853 16201 16865 16204
rect 16899 16201 16911 16235
rect 16853 16195 16911 16201
rect 19260 16204 20208 16232
rect 16666 16124 16672 16176
rect 16724 16164 16730 16176
rect 16942 16164 16948 16176
rect 16724 16136 16948 16164
rect 16724 16124 16730 16136
rect 16942 16124 16948 16136
rect 17000 16164 17006 16176
rect 19260 16164 19288 16204
rect 17000 16136 19288 16164
rect 19337 16167 19395 16173
rect 17000 16124 17006 16136
rect 19337 16133 19349 16167
rect 19383 16164 19395 16167
rect 19886 16164 19892 16176
rect 19383 16136 19892 16164
rect 19383 16133 19395 16136
rect 19337 16127 19395 16133
rect 19886 16124 19892 16136
rect 19944 16124 19950 16176
rect 20180 16164 20208 16204
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 20349 16235 20407 16241
rect 20349 16232 20361 16235
rect 20312 16204 20361 16232
rect 20312 16192 20318 16204
rect 20349 16201 20361 16204
rect 20395 16201 20407 16235
rect 20349 16195 20407 16201
rect 20180 16136 20944 16164
rect 16390 16056 16396 16108
rect 16448 16096 16454 16108
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 16448 16068 17417 16096
rect 16448 16056 16454 16068
rect 17405 16065 17417 16068
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 18506 16056 18512 16108
rect 18564 16096 18570 16108
rect 18601 16099 18659 16105
rect 18601 16096 18613 16099
rect 18564 16068 18613 16096
rect 18564 16056 18570 16068
rect 18601 16065 18613 16068
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 19702 16096 19708 16108
rect 19300 16068 19708 16096
rect 19300 16056 19306 16068
rect 19702 16056 19708 16068
rect 19760 16056 19766 16108
rect 19978 16096 19984 16108
rect 19939 16068 19984 16096
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 20622 16056 20628 16108
rect 20680 16096 20686 16108
rect 20916 16105 20944 16136
rect 20809 16099 20867 16105
rect 20809 16096 20821 16099
rect 20680 16068 20821 16096
rect 20680 16056 20686 16068
rect 20809 16065 20821 16068
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 14507 16000 15148 16028
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 15470 16037 15476 16040
rect 15464 16028 15476 16037
rect 15252 16000 15297 16028
rect 15431 16000 15476 16028
rect 15252 15988 15258 16000
rect 15464 15991 15476 16000
rect 15470 15988 15476 15991
rect 15528 15988 15534 16040
rect 16574 15988 16580 16040
rect 16632 16028 16638 16040
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 16632 16000 17233 16028
rect 16632 15988 16638 16000
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 18417 16031 18475 16037
rect 18417 15997 18429 16031
rect 18463 16028 18475 16031
rect 19334 16028 19340 16040
rect 18463 16000 19340 16028
rect 18463 15997 18475 16000
rect 18417 15991 18475 15997
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 20714 16028 20720 16040
rect 20675 16000 20720 16028
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 12710 15969 12716 15972
rect 12704 15960 12716 15969
rect 12671 15932 12716 15960
rect 12704 15923 12716 15932
rect 12710 15920 12716 15923
rect 12768 15920 12774 15972
rect 13354 15920 13360 15972
rect 13412 15920 13418 15972
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 18509 15963 18567 15969
rect 18509 15960 18521 15963
rect 18196 15932 18521 15960
rect 18196 15920 18202 15932
rect 18509 15929 18521 15932
rect 18555 15929 18567 15963
rect 18509 15923 18567 15929
rect 16482 15892 16488 15904
rect 11440 15864 16488 15892
rect 11241 15855 11299 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 16577 15895 16635 15901
rect 16577 15861 16589 15895
rect 16623 15892 16635 15895
rect 16666 15892 16672 15904
rect 16623 15864 16672 15892
rect 16623 15861 16635 15864
rect 16577 15855 16635 15861
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 17184 15864 17325 15892
rect 17184 15852 17190 15864
rect 17313 15861 17325 15864
rect 17359 15892 17371 15895
rect 17770 15892 17776 15904
rect 17359 15864 17776 15892
rect 17359 15861 17371 15864
rect 17313 15855 17371 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 18046 15892 18052 15904
rect 18007 15864 18052 15892
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 19702 15892 19708 15904
rect 19663 15864 19708 15892
rect 19702 15852 19708 15864
rect 19760 15852 19766 15904
rect 19794 15852 19800 15904
rect 19852 15892 19858 15904
rect 19852 15864 19897 15892
rect 19852 15852 19858 15864
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2866 15688 2872 15700
rect 2827 15660 2872 15688
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 2961 15691 3019 15697
rect 2961 15657 2973 15691
rect 3007 15688 3019 15691
rect 3142 15688 3148 15700
rect 3007 15660 3148 15688
rect 3007 15657 3019 15660
rect 2961 15651 3019 15657
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 3418 15688 3424 15700
rect 3379 15660 3424 15688
rect 3418 15648 3424 15660
rect 3476 15648 3482 15700
rect 4062 15688 4068 15700
rect 4023 15660 4068 15688
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4433 15691 4491 15697
rect 4433 15657 4445 15691
rect 4479 15688 4491 15691
rect 4798 15688 4804 15700
rect 4479 15660 4804 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 5552 15660 7512 15688
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 2317 15623 2375 15629
rect 2317 15620 2329 15623
rect 1452 15592 2329 15620
rect 1452 15580 1458 15592
rect 2317 15589 2329 15592
rect 2363 15589 2375 15623
rect 2317 15583 2375 15589
rect 2774 15580 2780 15632
rect 2832 15620 2838 15632
rect 5552 15620 5580 15660
rect 2832 15592 5580 15620
rect 7484 15620 7512 15660
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 8478 15688 8484 15700
rect 7616 15660 8484 15688
rect 7616 15648 7622 15660
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 10229 15691 10287 15697
rect 10229 15657 10241 15691
rect 10275 15657 10287 15691
rect 10594 15688 10600 15700
rect 10555 15660 10600 15688
rect 10229 15651 10287 15657
rect 8573 15623 8631 15629
rect 8573 15620 8585 15623
rect 7484 15592 8585 15620
rect 2832 15580 2838 15592
rect 8573 15589 8585 15592
rect 8619 15589 8631 15623
rect 9030 15620 9036 15632
rect 8991 15592 9036 15620
rect 8573 15583 8631 15589
rect 9030 15580 9036 15592
rect 9088 15580 9094 15632
rect 10244 15620 10272 15651
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 11149 15691 11207 15697
rect 10744 15660 10789 15688
rect 10744 15648 10750 15660
rect 11149 15657 11161 15691
rect 11195 15688 11207 15691
rect 12618 15688 12624 15700
rect 11195 15660 12624 15688
rect 11195 15657 11207 15660
rect 11149 15651 11207 15657
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 12897 15691 12955 15697
rect 12897 15657 12909 15691
rect 12943 15688 12955 15691
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 12943 15660 14381 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 14369 15657 14381 15660
rect 14415 15657 14427 15691
rect 14369 15651 14427 15657
rect 15289 15691 15347 15697
rect 15289 15657 15301 15691
rect 15335 15688 15347 15691
rect 16758 15688 16764 15700
rect 15335 15660 16764 15688
rect 15335 15657 15347 15660
rect 15289 15651 15347 15657
rect 16758 15648 16764 15660
rect 16816 15648 16822 15700
rect 18046 15648 18052 15700
rect 18104 15688 18110 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 18104 15660 18705 15688
rect 18104 15648 18110 15660
rect 18693 15657 18705 15660
rect 18739 15657 18751 15691
rect 18693 15651 18751 15657
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 20438 15688 20444 15700
rect 18840 15660 20300 15688
rect 20399 15660 20444 15688
rect 18840 15648 18846 15660
rect 13357 15623 13415 15629
rect 13357 15620 13369 15623
rect 10244 15592 13369 15620
rect 13357 15589 13369 15592
rect 13403 15589 13415 15623
rect 14274 15620 14280 15632
rect 14235 15592 14280 15620
rect 13357 15583 13415 15589
rect 14274 15580 14280 15592
rect 14332 15580 14338 15632
rect 15657 15623 15715 15629
rect 15657 15589 15669 15623
rect 15703 15620 15715 15623
rect 16206 15620 16212 15632
rect 15703 15592 16212 15620
rect 15703 15589 15715 15592
rect 15657 15583 15715 15589
rect 1486 15552 1492 15564
rect 1447 15524 1492 15552
rect 1486 15512 1492 15524
rect 1544 15512 1550 15564
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15552 2099 15555
rect 2685 15555 2743 15561
rect 2685 15552 2697 15555
rect 2087 15524 2697 15552
rect 2087 15521 2099 15524
rect 2041 15515 2099 15521
rect 2685 15521 2697 15524
rect 2731 15521 2743 15555
rect 2685 15515 2743 15521
rect 2866 15512 2872 15564
rect 2924 15552 2930 15564
rect 3329 15555 3387 15561
rect 3329 15552 3341 15555
rect 2924 15524 3341 15552
rect 2924 15512 2930 15524
rect 3329 15521 3341 15524
rect 3375 15521 3387 15555
rect 3329 15515 3387 15521
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 4890 15552 4896 15564
rect 4571 15524 4896 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5701 15555 5759 15561
rect 5701 15552 5713 15555
rect 5592 15524 5713 15552
rect 5592 15512 5598 15524
rect 5701 15521 5713 15524
rect 5747 15521 5759 15555
rect 5701 15515 5759 15521
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 6972 15524 7113 15552
rect 6972 15512 6978 15524
rect 7101 15521 7113 15524
rect 7147 15521 7159 15555
rect 7368 15555 7426 15561
rect 7368 15552 7380 15555
rect 7101 15515 7159 15521
rect 7208 15524 7380 15552
rect 1504 15484 1532 15512
rect 2130 15484 2136 15496
rect 1504 15456 2136 15484
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 3510 15444 3516 15496
rect 3568 15484 3574 15496
rect 3786 15484 3792 15496
rect 3568 15456 3792 15484
rect 3568 15444 3574 15456
rect 3786 15444 3792 15456
rect 3844 15484 3850 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 3844 15456 4629 15484
rect 3844 15444 3850 15456
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 5442 15484 5448 15496
rect 5403 15456 5448 15484
rect 4617 15447 4675 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 7208 15484 7236 15524
rect 7368 15521 7380 15524
rect 7414 15552 7426 15555
rect 8757 15555 8815 15561
rect 7414 15524 8708 15552
rect 7414 15521 7426 15524
rect 7368 15515 7426 15521
rect 6840 15456 7236 15484
rect 8680 15484 8708 15524
rect 8757 15521 8769 15555
rect 8803 15552 8815 15555
rect 9674 15552 9680 15564
rect 8803 15524 9680 15552
rect 8803 15521 8815 15524
rect 8757 15515 8815 15521
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 10410 15512 10416 15564
rect 10468 15552 10474 15564
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 10468 15524 11253 15552
rect 10468 15512 10474 15524
rect 11241 15521 11253 15524
rect 11287 15552 11299 15555
rect 11330 15552 11336 15564
rect 11287 15524 11336 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 11508 15555 11566 15561
rect 11508 15521 11520 15555
rect 11554 15552 11566 15555
rect 12250 15552 12256 15564
rect 11554 15524 12256 15552
rect 11554 15521 11566 15524
rect 11508 15515 11566 15521
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 13262 15552 13268 15564
rect 13223 15524 13268 15552
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 15672 15552 15700 15583
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 16844 15623 16902 15629
rect 16844 15589 16856 15623
rect 16890 15620 16902 15623
rect 18506 15620 18512 15632
rect 16890 15592 18512 15620
rect 16890 15589 16902 15592
rect 16844 15583 16902 15589
rect 18506 15580 18512 15592
rect 18564 15620 18570 15632
rect 19150 15620 19156 15632
rect 18564 15592 19156 15620
rect 18564 15580 18570 15592
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 19242 15580 19248 15632
rect 19300 15620 19306 15632
rect 19705 15623 19763 15629
rect 19705 15620 19717 15623
rect 19300 15592 19717 15620
rect 19300 15580 19306 15592
rect 19705 15589 19717 15592
rect 19751 15589 19763 15623
rect 19705 15583 19763 15589
rect 16298 15552 16304 15564
rect 13372 15524 15700 15552
rect 15948 15524 16304 15552
rect 8938 15484 8944 15496
rect 8680 15456 8944 15484
rect 2685 15419 2743 15425
rect 2685 15385 2697 15419
rect 2731 15416 2743 15419
rect 2731 15388 5488 15416
rect 2731 15385 2743 15388
rect 2685 15379 2743 15385
rect 2498 15308 2504 15360
rect 2556 15348 2562 15360
rect 2958 15348 2964 15360
rect 2556 15320 2964 15348
rect 2556 15308 2562 15320
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 5460 15348 5488 15388
rect 6454 15376 6460 15428
rect 6512 15416 6518 15428
rect 6840 15425 6868 15456
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 10778 15484 10784 15496
rect 10739 15456 10784 15484
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 13372 15484 13400 15524
rect 12676 15456 13400 15484
rect 13449 15487 13507 15493
rect 12676 15444 12682 15456
rect 13449 15453 13461 15487
rect 13495 15453 13507 15487
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 13449 15447 13507 15453
rect 13556 15456 14473 15484
rect 6825 15419 6883 15425
rect 6825 15416 6837 15419
rect 6512 15388 6837 15416
rect 6512 15376 6518 15388
rect 6825 15385 6837 15388
rect 6871 15385 6883 15419
rect 6825 15379 6883 15385
rect 8573 15419 8631 15425
rect 8573 15385 8585 15419
rect 8619 15416 8631 15419
rect 11149 15419 11207 15425
rect 11149 15416 11161 15419
rect 8619 15388 11161 15416
rect 8619 15385 8631 15388
rect 8573 15379 8631 15385
rect 9048 15360 9076 15388
rect 11149 15385 11161 15388
rect 11195 15385 11207 15419
rect 11149 15379 11207 15385
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 13464 15416 13492 15447
rect 12308 15388 13492 15416
rect 12308 15376 12314 15388
rect 8202 15348 8208 15360
rect 5460 15320 8208 15348
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 12621 15351 12679 15357
rect 12621 15317 12633 15351
rect 12667 15348 12679 15351
rect 12710 15348 12716 15360
rect 12667 15320 12716 15348
rect 12667 15317 12679 15320
rect 12621 15311 12679 15317
rect 12710 15308 12716 15320
rect 12768 15348 12774 15360
rect 13556 15348 13584 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 15838 15484 15844 15496
rect 15795 15456 15844 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 15948 15493 15976 15524
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15552 16543 15555
rect 16577 15555 16635 15561
rect 16577 15552 16589 15555
rect 16531 15524 16589 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 16577 15521 16589 15524
rect 16623 15521 16635 15555
rect 18598 15552 18604 15564
rect 18559 15524 18604 15552
rect 16577 15515 16635 15521
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 20272 15561 20300 15660
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 18748 15524 19625 15552
rect 18748 15512 18754 15524
rect 19613 15521 19625 15524
rect 19659 15552 19671 15555
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 19659 15524 20085 15552
rect 19659 15521 19671 15524
rect 19613 15515 19671 15521
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20073 15515 20131 15521
rect 20257 15555 20315 15561
rect 20257 15521 20269 15555
rect 20303 15521 20315 15555
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20257 15515 20315 15521
rect 20364 15524 20913 15552
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15484 18199 15487
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 18187 15456 18797 15484
rect 18187 15453 18199 15456
rect 18141 15447 18199 15453
rect 18785 15453 18797 15456
rect 18831 15453 18843 15487
rect 18785 15447 18843 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 20162 15484 20168 15496
rect 19935 15456 20168 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 13909 15419 13967 15425
rect 13909 15385 13921 15419
rect 13955 15416 13967 15419
rect 14366 15416 14372 15428
rect 13955 15388 14372 15416
rect 13955 15385 13967 15388
rect 13909 15379 13967 15385
rect 14366 15376 14372 15388
rect 14424 15376 14430 15428
rect 18233 15419 18291 15425
rect 18233 15385 18245 15419
rect 18279 15416 18291 15419
rect 20364 15416 20392 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 20806 15444 20812 15496
rect 20864 15484 20870 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 20864 15456 21097 15484
rect 20864 15444 20870 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 18279 15388 20392 15416
rect 18279 15385 18291 15388
rect 18233 15379 18291 15385
rect 12768 15320 13584 15348
rect 12768 15308 12774 15320
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15470 15348 15476 15360
rect 15252 15320 15476 15348
rect 15252 15308 15258 15320
rect 15470 15308 15476 15320
rect 15528 15348 15534 15360
rect 16482 15348 16488 15360
rect 15528 15320 16488 15348
rect 15528 15308 15534 15320
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 17770 15308 17776 15360
rect 17828 15348 17834 15360
rect 17957 15351 18015 15357
rect 17957 15348 17969 15351
rect 17828 15320 17969 15348
rect 17828 15308 17834 15320
rect 17957 15317 17969 15320
rect 18003 15348 18015 15351
rect 18049 15351 18107 15357
rect 18049 15348 18061 15351
rect 18003 15320 18061 15348
rect 18003 15317 18015 15320
rect 17957 15311 18015 15317
rect 18049 15317 18061 15320
rect 18095 15317 18107 15351
rect 19242 15348 19248 15360
rect 19203 15320 19248 15348
rect 18049 15311 18107 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 20073 15351 20131 15357
rect 20073 15317 20085 15351
rect 20119 15348 20131 15351
rect 21174 15348 21180 15360
rect 20119 15320 21180 15348
rect 20119 15317 20131 15320
rect 20073 15311 20131 15317
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1854 15144 1860 15156
rect 1815 15116 1860 15144
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 3234 15144 3240 15156
rect 3195 15116 3240 15144
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 3418 15104 3424 15156
rect 3476 15144 3482 15156
rect 3970 15144 3976 15156
rect 3476 15116 3976 15144
rect 3476 15104 3482 15116
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 6270 15144 6276 15156
rect 4080 15116 6276 15144
rect 4080 15076 4108 15116
rect 6270 15104 6276 15116
rect 6328 15144 6334 15156
rect 6638 15144 6644 15156
rect 6328 15116 6644 15144
rect 6328 15104 6334 15116
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7098 15144 7104 15156
rect 6972 15116 7104 15144
rect 6972 15104 6978 15116
rect 7098 15104 7104 15116
rect 7156 15144 7162 15156
rect 7834 15144 7840 15156
rect 7156 15116 7840 15144
rect 7156 15104 7162 15116
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 7929 15147 7987 15153
rect 7929 15113 7941 15147
rect 7975 15144 7987 15147
rect 10042 15144 10048 15156
rect 7975 15116 10048 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 11885 15147 11943 15153
rect 11885 15113 11897 15147
rect 11931 15144 11943 15147
rect 12250 15144 12256 15156
rect 11931 15116 12256 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12492 15116 12537 15144
rect 12492 15104 12498 15116
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13412 15116 13461 15144
rect 13412 15104 13418 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 14090 15144 14096 15156
rect 14051 15116 14096 15144
rect 13449 15107 13507 15113
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 14274 15104 14280 15156
rect 14332 15144 14338 15156
rect 15378 15144 15384 15156
rect 14332 15116 15384 15144
rect 14332 15104 14338 15116
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 17954 15144 17960 15156
rect 15519 15116 17960 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 19429 15147 19487 15153
rect 19429 15144 19441 15147
rect 19208 15116 19441 15144
rect 19208 15104 19214 15116
rect 19429 15113 19441 15116
rect 19475 15113 19487 15147
rect 20990 15144 20996 15156
rect 20951 15116 20996 15144
rect 19429 15107 19487 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 1688 15048 4108 15076
rect 4249 15079 4307 15085
rect 1688 14949 1716 15048
rect 4249 15045 4261 15079
rect 4295 15045 4307 15079
rect 4249 15039 4307 15045
rect 3786 15008 3792 15020
rect 3747 14980 3792 15008
rect 3786 14968 3792 14980
rect 3844 14968 3850 15020
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14909 1731 14943
rect 1673 14903 1731 14909
rect 2225 14943 2283 14949
rect 2225 14909 2237 14943
rect 2271 14940 2283 14943
rect 4264 14940 4292 15039
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 7558 15076 7564 15088
rect 6880 15048 7564 15076
rect 6880 15036 6886 15048
rect 7558 15036 7564 15048
rect 7616 15036 7622 15088
rect 7650 15036 7656 15088
rect 7708 15076 7714 15088
rect 10134 15076 10140 15088
rect 7708 15048 10140 15076
rect 7708 15036 7714 15048
rect 10134 15036 10140 15048
rect 10192 15036 10198 15088
rect 11514 15036 11520 15088
rect 11572 15076 11578 15088
rect 11572 15048 15424 15076
rect 11572 15036 11578 15048
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5626 15008 5632 15020
rect 4939 14980 5632 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 5905 15011 5963 15017
rect 5776 14980 5821 15008
rect 5776 14968 5782 14980
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6270 15008 6276 15020
rect 5951 14980 6276 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 8478 15008 8484 15020
rect 8439 14980 8484 15008
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8754 14968 8760 15020
rect 8812 15008 8818 15020
rect 9582 15008 9588 15020
rect 8812 14980 9588 15008
rect 8812 14968 8818 14980
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 9732 14980 9777 15008
rect 9732 14968 9738 14980
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12492 14980 13001 15008
rect 12492 14968 12498 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 14642 15008 14648 15020
rect 14603 14980 14648 15008
rect 12989 14971 13047 14977
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 2271 14912 4292 14940
rect 2271 14909 2283 14912
rect 2225 14903 2283 14909
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 6454 14940 6460 14952
rect 5316 14912 5672 14940
rect 6367 14912 6460 14940
rect 5316 14900 5322 14912
rect 1762 14832 1768 14884
rect 1820 14872 1826 14884
rect 5644 14881 5672 14912
rect 6454 14900 6460 14912
rect 6512 14940 6518 14952
rect 7193 14943 7251 14949
rect 6512 14912 6776 14940
rect 6512 14900 6518 14912
rect 2501 14875 2559 14881
rect 2501 14872 2513 14875
rect 1820 14844 2513 14872
rect 1820 14832 1826 14844
rect 2501 14841 2513 14844
rect 2547 14841 2559 14875
rect 2501 14835 2559 14841
rect 3145 14875 3203 14881
rect 3145 14841 3157 14875
rect 3191 14872 3203 14875
rect 5629 14875 5687 14881
rect 3191 14844 3740 14872
rect 3191 14841 3203 14844
rect 3145 14835 3203 14841
rect 3326 14764 3332 14816
rect 3384 14804 3390 14816
rect 3602 14804 3608 14816
rect 3384 14776 3608 14804
rect 3384 14764 3390 14776
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 3712 14813 3740 14844
rect 5629 14841 5641 14875
rect 5675 14841 5687 14875
rect 5629 14835 5687 14841
rect 5810 14832 5816 14884
rect 5868 14872 5874 14884
rect 5994 14872 6000 14884
rect 5868 14844 6000 14872
rect 5868 14832 5874 14844
rect 5994 14832 6000 14844
rect 6052 14832 6058 14884
rect 6748 14872 6776 14912
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 8018 14940 8024 14952
rect 7239 14912 8024 14940
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 8294 14940 8300 14952
rect 8255 14912 8300 14940
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 8386 14900 8392 14952
rect 8444 14940 8450 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 8444 14912 8489 14940
rect 8588 14912 10333 14940
rect 8444 14900 8450 14912
rect 8588 14872 8616 14912
rect 10321 14909 10333 14912
rect 10367 14909 10379 14943
rect 10321 14903 10379 14909
rect 10410 14900 10416 14952
rect 10468 14940 10474 14952
rect 10778 14949 10784 14952
rect 10505 14943 10563 14949
rect 10505 14940 10517 14943
rect 10468 14912 10517 14940
rect 10468 14900 10474 14912
rect 10505 14909 10517 14912
rect 10551 14909 10563 14943
rect 10772 14940 10784 14949
rect 10691 14912 10784 14940
rect 10505 14903 10563 14909
rect 10772 14903 10784 14912
rect 10836 14940 10842 14952
rect 12452 14940 12480 14968
rect 10836 14912 12480 14940
rect 10778 14900 10784 14903
rect 10836 14900 10842 14912
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 12676 14912 12817 14940
rect 12676 14900 12682 14912
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13722 14940 13728 14952
rect 13679 14912 13728 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 15286 14940 15292 14952
rect 15247 14912 15292 14940
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 6748 14844 8616 14872
rect 9033 14875 9091 14881
rect 9033 14841 9045 14875
rect 9079 14872 9091 14875
rect 9585 14875 9643 14881
rect 9585 14872 9597 14875
rect 9079 14844 9597 14872
rect 9079 14841 9091 14844
rect 9033 14835 9091 14841
rect 9585 14841 9597 14844
rect 9631 14872 9643 14875
rect 15102 14872 15108 14884
rect 9631 14844 10364 14872
rect 9631 14841 9643 14844
rect 9585 14835 9643 14841
rect 3697 14807 3755 14813
rect 3697 14773 3709 14807
rect 3743 14804 3755 14807
rect 4062 14804 4068 14816
rect 3743 14776 4068 14804
rect 3743 14773 3755 14776
rect 3697 14767 3755 14773
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4338 14764 4344 14816
rect 4396 14804 4402 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4396 14776 4629 14804
rect 4396 14764 4402 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 4617 14767 4675 14773
rect 4709 14807 4767 14813
rect 4709 14773 4721 14807
rect 4755 14804 4767 14807
rect 5074 14804 5080 14816
rect 4755 14776 5080 14804
rect 4755 14773 4767 14776
rect 4709 14767 4767 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 5261 14807 5319 14813
rect 5261 14804 5273 14807
rect 5224 14776 5273 14804
rect 5224 14764 5230 14776
rect 5261 14773 5273 14776
rect 5307 14773 5319 14807
rect 5261 14767 5319 14773
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 6273 14807 6331 14813
rect 6273 14804 6285 14807
rect 5500 14776 6285 14804
rect 5500 14764 5506 14776
rect 6273 14773 6285 14776
rect 6319 14804 6331 14807
rect 6362 14804 6368 14816
rect 6319 14776 6368 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 8478 14804 8484 14816
rect 7331 14776 8484 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9122 14804 9128 14816
rect 9083 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9490 14804 9496 14816
rect 9451 14776 9496 14804
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 10336 14804 10364 14844
rect 10888 14844 15108 14872
rect 10888 14804 10916 14844
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 15396 14872 15424 15048
rect 20162 15036 20168 15088
rect 20220 15076 20226 15088
rect 20220 15048 20392 15076
rect 20220 15036 20226 15048
rect 20364 15020 20392 15048
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 20346 15008 20352 15020
rect 17460 14980 18184 15008
rect 20307 14980 20352 15008
rect 17460 14968 17466 14980
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 15841 14943 15899 14949
rect 15841 14940 15853 14943
rect 15528 14912 15853 14940
rect 15528 14900 15534 14912
rect 15841 14909 15853 14912
rect 15887 14909 15899 14943
rect 15841 14903 15899 14909
rect 16108 14943 16166 14949
rect 16108 14909 16120 14943
rect 16154 14940 16166 14943
rect 17770 14940 17776 14952
rect 16154 14912 17776 14940
rect 16154 14909 16166 14912
rect 16108 14903 16166 14909
rect 17770 14900 17776 14912
rect 17828 14900 17834 14952
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14909 18107 14943
rect 18156 14940 18184 14980
rect 20346 14968 20352 14980
rect 20404 14968 20410 15020
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 18156 14912 20177 14940
rect 18049 14903 18107 14909
rect 20165 14909 20177 14912
rect 20211 14940 20223 14943
rect 20254 14940 20260 14952
rect 20211 14912 20260 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 16942 14872 16948 14884
rect 15396 14844 16948 14872
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 18064 14872 18092 14903
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 20806 14940 20812 14952
rect 20767 14912 20812 14940
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 17144 14844 18092 14872
rect 18316 14875 18374 14881
rect 10336 14776 10916 14804
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12584 14776 12909 14804
rect 12584 14764 12590 14776
rect 12897 14773 12909 14776
rect 12943 14804 12955 14807
rect 13906 14804 13912 14816
rect 12943 14776 13912 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14458 14804 14464 14816
rect 14419 14776 14464 14804
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 14608 14776 14653 14804
rect 14608 14764 14614 14776
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 16298 14804 16304 14816
rect 14792 14776 16304 14804
rect 14792 14764 14798 14776
rect 16298 14764 16304 14776
rect 16356 14764 16362 14816
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 17144 14804 17172 14844
rect 18316 14841 18328 14875
rect 18362 14872 18374 14875
rect 18690 14872 18696 14884
rect 18362 14844 18696 14872
rect 18362 14841 18374 14844
rect 18316 14835 18374 14841
rect 18690 14832 18696 14844
rect 18748 14832 18754 14884
rect 20073 14875 20131 14881
rect 20073 14872 20085 14875
rect 18800 14844 20085 14872
rect 16540 14776 17172 14804
rect 17221 14807 17279 14813
rect 16540 14764 16546 14776
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 17402 14804 17408 14816
rect 17267 14776 17408 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 17497 14807 17555 14813
rect 17497 14773 17509 14807
rect 17543 14804 17555 14807
rect 18800 14804 18828 14844
rect 20073 14841 20085 14844
rect 20119 14841 20131 14875
rect 20073 14835 20131 14841
rect 17543 14776 18828 14804
rect 19705 14807 19763 14813
rect 17543 14773 17555 14776
rect 17497 14767 17555 14773
rect 19705 14773 19717 14807
rect 19751 14804 19763 14807
rect 20162 14804 20168 14816
rect 19751 14776 20168 14804
rect 19751 14773 19763 14776
rect 19705 14767 19763 14773
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 3510 14600 3516 14612
rect 3471 14572 3516 14600
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 4304 14572 4375 14600
rect 4304 14560 4310 14572
rect 2777 14535 2835 14541
rect 2777 14501 2789 14535
rect 2823 14532 2835 14535
rect 3970 14532 3976 14544
rect 2823 14504 3976 14532
rect 2823 14501 2835 14504
rect 2777 14495 2835 14501
rect 3970 14492 3976 14504
rect 4028 14492 4034 14544
rect 4347 14541 4375 14572
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 5776 14572 6776 14600
rect 5776 14560 5782 14572
rect 4332 14535 4390 14541
rect 4332 14501 4344 14535
rect 4378 14532 4390 14535
rect 5534 14532 5540 14544
rect 4378 14504 5540 14532
rect 4378 14501 4390 14504
rect 4332 14495 4390 14501
rect 5534 14492 5540 14504
rect 5592 14532 5598 14544
rect 6641 14535 6699 14541
rect 6641 14532 6653 14535
rect 5592 14504 6653 14532
rect 5592 14492 5598 14504
rect 6641 14501 6653 14504
rect 6687 14501 6699 14535
rect 6748 14532 6776 14572
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 6880 14572 7205 14600
rect 6880 14560 6886 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 8754 14600 8760 14612
rect 7193 14563 7251 14569
rect 8220 14572 8760 14600
rect 8220 14532 8248 14572
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8904 14572 8953 14600
rect 8904 14560 8910 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 11514 14600 11520 14612
rect 9640 14572 11520 14600
rect 9640 14560 9646 14572
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 12710 14600 12716 14612
rect 11839 14572 12716 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 15289 14603 15347 14609
rect 12912 14572 14587 14600
rect 6748 14504 8248 14532
rect 8297 14535 8355 14541
rect 6641 14495 6699 14501
rect 8297 14501 8309 14535
rect 8343 14532 8355 14535
rect 10042 14532 10048 14544
rect 8343 14504 10048 14532
rect 8343 14501 8355 14504
rect 8297 14495 8355 14501
rect 10042 14492 10048 14504
rect 10100 14492 10106 14544
rect 10404 14535 10462 14541
rect 10404 14501 10416 14535
rect 10450 14532 10462 14535
rect 10962 14532 10968 14544
rect 10450 14504 10968 14532
rect 10450 14501 10462 14504
rect 10404 14495 10462 14501
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2406 14424 2412 14476
rect 2464 14464 2470 14476
rect 2685 14467 2743 14473
rect 2685 14464 2697 14467
rect 2464 14436 2697 14464
rect 2464 14424 2470 14436
rect 2685 14433 2697 14436
rect 2731 14433 2743 14467
rect 2685 14427 2743 14433
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14464 3387 14467
rect 6089 14467 6147 14473
rect 3375 14436 6040 14464
rect 3375 14433 3387 14436
rect 3329 14427 3387 14433
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 4065 14399 4123 14405
rect 3007 14368 3372 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3344 14340 3372 14368
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 3326 14288 3332 14340
rect 3384 14288 3390 14340
rect 2038 14220 2044 14272
rect 2096 14260 2102 14272
rect 2317 14263 2375 14269
rect 2317 14260 2329 14263
rect 2096 14232 2329 14260
rect 2096 14220 2102 14232
rect 2317 14229 2329 14232
rect 2363 14229 2375 14263
rect 2317 14223 2375 14229
rect 3050 14220 3056 14272
rect 3108 14260 3114 14272
rect 4080 14260 4108 14359
rect 6012 14328 6040 14436
rect 6089 14433 6101 14467
rect 6135 14464 6147 14467
rect 6914 14464 6920 14476
rect 6135 14436 6920 14464
rect 6135 14433 6147 14436
rect 6089 14427 6147 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7098 14464 7104 14476
rect 7059 14436 7104 14464
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 9674 14464 9680 14476
rect 8435 14436 9680 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 10134 14464 10140 14476
rect 10095 14436 10140 14464
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 10778 14464 10784 14476
rect 10244 14436 10784 14464
rect 6178 14396 6184 14408
rect 6139 14368 6184 14396
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 6411 14368 6653 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 6641 14365 6653 14368
rect 6687 14396 6699 14399
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 6687 14368 7297 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 8478 14396 8484 14408
rect 8439 14368 8484 14396
rect 7285 14359 7343 14365
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 10244 14396 10272 14436
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 12158 14464 12164 14476
rect 12119 14436 12164 14464
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12250 14396 12256 14408
rect 8996 14368 10272 14396
rect 12211 14368 12256 14396
rect 8996 14356 9002 14368
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 12434 14396 12440 14408
rect 12395 14368 12440 14396
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 6546 14328 6552 14340
rect 6012 14300 6552 14328
rect 6546 14288 6552 14300
rect 6604 14328 6610 14340
rect 9490 14328 9496 14340
rect 6604 14300 9496 14328
rect 6604 14288 6610 14300
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 11517 14331 11575 14337
rect 11517 14297 11529 14331
rect 11563 14328 11575 14331
rect 11698 14328 11704 14340
rect 11563 14300 11704 14328
rect 11563 14297 11575 14300
rect 11517 14291 11575 14297
rect 11698 14288 11704 14300
rect 11756 14328 11762 14340
rect 12452 14328 12480 14356
rect 11756 14300 12480 14328
rect 11756 14288 11762 14300
rect 4798 14260 4804 14272
rect 3108 14232 4804 14260
rect 3108 14220 3114 14232
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 5442 14260 5448 14272
rect 5403 14232 5448 14260
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5718 14260 5724 14272
rect 5679 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6733 14263 6791 14269
rect 6733 14260 6745 14263
rect 5868 14232 6745 14260
rect 5868 14220 5874 14232
rect 6733 14229 6745 14232
rect 6779 14229 6791 14263
rect 6733 14223 6791 14229
rect 7929 14263 7987 14269
rect 7929 14229 7941 14263
rect 7975 14260 7987 14263
rect 8846 14260 8852 14272
rect 7975 14232 8852 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 8938 14220 8944 14272
rect 8996 14260 9002 14272
rect 12912 14260 12940 14572
rect 13630 14492 13636 14544
rect 13688 14492 13694 14544
rect 14274 14492 14280 14544
rect 14332 14532 14338 14544
rect 14461 14535 14519 14541
rect 14461 14532 14473 14535
rect 14332 14504 14473 14532
rect 14332 14492 14338 14504
rect 14461 14501 14473 14504
rect 14507 14501 14519 14535
rect 14461 14495 14519 14501
rect 13354 14464 13360 14476
rect 13315 14436 13360 14464
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13648 14396 13676 14492
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 14559 14464 14587 14572
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 16761 14603 16819 14609
rect 16761 14600 16773 14603
rect 15335 14572 16773 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 16761 14569 16773 14572
rect 16807 14569 16819 14603
rect 16761 14563 16819 14569
rect 18598 14560 18604 14612
rect 18656 14600 18662 14612
rect 18785 14603 18843 14609
rect 18785 14600 18797 14603
rect 18656 14572 18797 14600
rect 18656 14560 18662 14572
rect 18785 14569 18797 14572
rect 18831 14569 18843 14603
rect 19242 14600 19248 14612
rect 19203 14572 19248 14600
rect 18785 14563 18843 14569
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19797 14603 19855 14609
rect 19797 14600 19809 14603
rect 19392 14572 19809 14600
rect 19392 14560 19398 14572
rect 19797 14569 19809 14572
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 20162 14560 20168 14612
rect 20220 14560 20226 14612
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 14826 14492 14832 14544
rect 14884 14532 14890 14544
rect 15470 14532 15476 14544
rect 14884 14504 15476 14532
rect 14884 14492 14890 14504
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 15654 14532 15660 14544
rect 15615 14504 15660 14532
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 15749 14535 15807 14541
rect 15749 14501 15761 14535
rect 15795 14532 15807 14535
rect 15838 14532 15844 14544
rect 15795 14504 15844 14532
rect 15795 14501 15807 14504
rect 15749 14495 15807 14501
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 18233 14535 18291 14541
rect 18233 14532 18245 14535
rect 15948 14504 18245 14532
rect 15948 14464 15976 14504
rect 18233 14501 18245 14504
rect 18279 14501 18291 14535
rect 18233 14495 18291 14501
rect 19153 14535 19211 14541
rect 19153 14501 19165 14535
rect 19199 14532 19211 14535
rect 20180 14532 20208 14560
rect 19199 14504 20208 14532
rect 19199 14501 19211 14504
rect 19153 14495 19211 14501
rect 14424 14436 14469 14464
rect 14559 14436 15976 14464
rect 14424 14424 14430 14436
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16669 14467 16727 14473
rect 16669 14464 16681 14467
rect 16632 14436 16681 14464
rect 16632 14424 16638 14436
rect 16669 14433 16681 14436
rect 16715 14433 16727 14467
rect 16669 14427 16727 14433
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 18104 14436 18153 14464
rect 18104 14424 18110 14436
rect 18141 14433 18153 14436
rect 18187 14433 18199 14467
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 18141 14427 18199 14433
rect 18248 14436 20177 14464
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 13587 14368 14565 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 14553 14365 14565 14368
rect 14599 14396 14611 14399
rect 15838 14396 15844 14408
rect 14599 14368 15844 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 13464 14328 13492 14359
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 16356 14368 16865 14396
rect 16356 14356 16362 14368
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 18248 14396 18276 14436
rect 20165 14433 20177 14436
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20772 14436 20913 14464
rect 20772 14424 20778 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 17092 14368 18276 14396
rect 18417 14399 18475 14405
rect 17092 14356 17098 14368
rect 18417 14365 18429 14399
rect 18463 14396 18475 14399
rect 18598 14396 18604 14408
rect 18463 14368 18604 14396
rect 18463 14365 18475 14368
rect 18417 14359 18475 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14365 19395 14399
rect 19337 14359 19395 14365
rect 13906 14328 13912 14340
rect 13464 14300 13912 14328
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 15930 14288 15936 14340
rect 15988 14328 15994 14340
rect 15988 14300 16804 14328
rect 15988 14288 15994 14300
rect 16776 14272 16804 14300
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19352 14328 19380 14359
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 20128 14368 20269 14396
rect 20128 14356 20134 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20404 14368 20449 14396
rect 20404 14356 20410 14368
rect 19208 14300 19380 14328
rect 19208 14288 19214 14300
rect 8996 14232 12940 14260
rect 12989 14263 13047 14269
rect 8996 14220 9002 14232
rect 12989 14229 13001 14263
rect 13035 14260 13047 14263
rect 13814 14260 13820 14272
rect 13035 14232 13820 14260
rect 13035 14229 13047 14232
rect 12989 14223 13047 14229
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 13998 14260 14004 14272
rect 13959 14232 14004 14260
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14550 14220 14556 14272
rect 14608 14260 14614 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 14608 14232 16313 14260
rect 14608 14220 14614 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 16758 14220 16764 14272
rect 16816 14220 16822 14272
rect 17770 14260 17776 14272
rect 17731 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 4433 14059 4491 14065
rect 4433 14056 4445 14059
rect 4304 14028 4445 14056
rect 4304 14016 4310 14028
rect 4433 14025 4445 14028
rect 4479 14025 4491 14059
rect 4433 14019 4491 14025
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 6089 14059 6147 14065
rect 6089 14056 6101 14059
rect 5684 14028 6101 14056
rect 5684 14016 5690 14028
rect 6089 14025 6101 14028
rect 6135 14025 6147 14059
rect 6454 14056 6460 14068
rect 6415 14028 6460 14056
rect 6089 14019 6147 14025
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3050 13920 3056 13932
rect 3011 13892 3056 13920
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 6104 13920 6132 14019
rect 6454 14016 6460 14028
rect 6512 14016 6518 14068
rect 8386 14016 8392 14068
rect 8444 14056 8450 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 8444 14028 11161 14056
rect 8444 14016 8450 14028
rect 11149 14025 11161 14028
rect 11195 14025 11207 14059
rect 11149 14019 11207 14025
rect 13081 14059 13139 14065
rect 13081 14025 13093 14059
rect 13127 14056 13139 14059
rect 13722 14056 13728 14068
rect 13127 14028 13728 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 13722 14016 13728 14028
rect 13780 14056 13786 14068
rect 15194 14056 15200 14068
rect 13780 14028 15200 14056
rect 13780 14016 13786 14028
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 16577 14059 16635 14065
rect 16577 14056 16589 14059
rect 15896 14028 16589 14056
rect 15896 14016 15902 14028
rect 16577 14025 16589 14028
rect 16623 14025 16635 14059
rect 16577 14019 16635 14025
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16816 14028 16865 14056
rect 16816 14016 16822 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 18690 14016 18696 14068
rect 18748 14056 18754 14068
rect 18748 14028 19472 14056
rect 18748 14016 18754 14028
rect 8481 13991 8539 13997
rect 8481 13957 8493 13991
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 9125 13991 9183 13997
rect 9125 13957 9137 13991
rect 9171 13988 9183 13991
rect 9398 13988 9404 14000
rect 9171 13960 9404 13988
rect 9171 13957 9183 13960
rect 9125 13951 9183 13957
rect 8496 13920 8524 13951
rect 9398 13948 9404 13960
rect 9456 13948 9462 14000
rect 10137 13991 10195 13997
rect 10137 13957 10149 13991
rect 10183 13957 10195 13991
rect 10137 13951 10195 13957
rect 9582 13920 9588 13932
rect 6104 13892 7236 13920
rect 8496 13892 9588 13920
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 2409 13855 2467 13861
rect 1443 13824 2360 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 2332 13784 2360 13824
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2958 13852 2964 13864
rect 2455 13824 2964 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 3602 13812 3608 13864
rect 3660 13852 3666 13864
rect 4246 13852 4252 13864
rect 3660 13824 4252 13852
rect 3660 13812 3666 13824
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4982 13861 4988 13864
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13821 4767 13855
rect 4976 13852 4988 13861
rect 4895 13824 4988 13852
rect 4709 13815 4767 13821
rect 4976 13815 4988 13824
rect 5040 13852 5046 13864
rect 5442 13852 5448 13864
rect 5040 13824 5448 13852
rect 3142 13784 3148 13796
rect 2332 13756 3148 13784
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 3320 13787 3378 13793
rect 3320 13753 3332 13787
rect 3366 13784 3378 13787
rect 3694 13784 3700 13796
rect 3366 13756 3700 13784
rect 3366 13753 3378 13756
rect 3320 13747 3378 13753
rect 3694 13744 3700 13756
rect 3752 13744 3758 13796
rect 4724 13784 4752 13815
rect 4982 13812 4988 13815
rect 5040 13812 5046 13824
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13852 6699 13855
rect 7006 13852 7012 13864
rect 6687 13824 7012 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13821 7159 13855
rect 7208 13852 7236 13892
rect 9582 13880 9588 13892
rect 9640 13920 9646 13932
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 9640 13892 9689 13920
rect 9640 13880 9646 13892
rect 9677 13889 9689 13892
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 10152 13920 10180 13951
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 12526 13988 12532 14000
rect 10376 13960 12532 13988
rect 10376 13948 10382 13960
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 12710 13948 12716 14000
rect 12768 13988 12774 14000
rect 13262 13988 13268 14000
rect 12768 13960 13268 13988
rect 12768 13948 12774 13960
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 14550 13948 14556 14000
rect 14608 13988 14614 14000
rect 14737 13991 14795 13997
rect 14737 13988 14749 13991
rect 14608 13960 14749 13988
rect 14608 13948 14614 13960
rect 14737 13957 14749 13960
rect 14783 13957 14795 13991
rect 14737 13951 14795 13957
rect 16298 13948 16304 14000
rect 16356 13988 16362 14000
rect 19444 13988 19472 14028
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 19760 14028 20085 14056
rect 19760 14016 19766 14028
rect 20073 14025 20085 14028
rect 20119 14025 20131 14059
rect 20073 14019 20131 14025
rect 19797 13991 19855 13997
rect 19797 13988 19809 13991
rect 16356 13960 18460 13988
rect 19444 13960 19809 13988
rect 16356 13948 16362 13960
rect 10778 13920 10784 13932
rect 10008 13892 10180 13920
rect 10691 13892 10784 13920
rect 10008 13880 10014 13892
rect 10778 13880 10784 13892
rect 10836 13920 10842 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 10836 13892 11713 13920
rect 10836 13880 10842 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12618 13920 12624 13932
rect 12483 13892 12624 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 17402 13920 17408 13932
rect 17363 13892 17408 13920
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 18432 13929 18460 13960
rect 19797 13957 19809 13960
rect 19843 13988 19855 13991
rect 20346 13988 20352 14000
rect 19843 13960 20352 13988
rect 19843 13957 19855 13960
rect 19797 13951 19855 13957
rect 20346 13948 20352 13960
rect 20404 13948 20410 14000
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20496 13892 20637 13920
rect 20496 13880 20502 13892
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 7357 13855 7415 13861
rect 7357 13852 7369 13855
rect 7208 13824 7369 13852
rect 7101 13815 7159 13821
rect 7357 13821 7369 13824
rect 7403 13821 7415 13855
rect 7357 13815 7415 13821
rect 4798 13784 4804 13796
rect 4711 13756 4804 13784
rect 4798 13744 4804 13756
rect 4856 13784 4862 13796
rect 6362 13784 6368 13796
rect 4856 13756 6368 13784
rect 4856 13744 4862 13756
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 7116 13784 7144 13815
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 10597 13855 10655 13861
rect 10597 13852 10609 13855
rect 9180 13824 10609 13852
rect 9180 13812 9186 13824
rect 10597 13821 10609 13824
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 11609 13855 11667 13861
rect 11609 13821 11621 13855
rect 11655 13852 11667 13855
rect 12342 13852 12348 13864
rect 11655 13824 12348 13852
rect 11655 13821 11667 13824
rect 11609 13815 11667 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13624 13855 13682 13861
rect 13412 13824 13457 13852
rect 13412 13812 13418 13824
rect 13624 13821 13636 13855
rect 13670 13852 13682 13855
rect 14734 13852 14740 13864
rect 13670 13824 14740 13852
rect 13670 13821 13682 13824
rect 13624 13815 13682 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 14826 13812 14832 13864
rect 14884 13852 14890 13864
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 14884 13824 15209 13852
rect 14884 13812 14890 13824
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 15464 13855 15522 13861
rect 15464 13821 15476 13855
rect 15510 13852 15522 13855
rect 15930 13852 15936 13864
rect 15510 13824 15936 13852
rect 15510 13821 15522 13824
rect 15464 13815 15522 13821
rect 15930 13812 15936 13824
rect 15988 13852 15994 13864
rect 17420 13852 17448 13880
rect 15988 13824 17448 13852
rect 15988 13812 15994 13824
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20312 13824 20545 13852
rect 20312 13812 20318 13824
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 21085 13855 21143 13861
rect 21085 13821 21097 13855
rect 21131 13852 21143 13855
rect 21174 13852 21180 13864
rect 21131 13824 21180 13852
rect 21131 13821 21143 13824
rect 21085 13815 21143 13821
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 7650 13784 7656 13796
rect 7116 13756 7656 13784
rect 7650 13744 7656 13756
rect 7708 13784 7714 13796
rect 8386 13784 8392 13796
rect 7708 13756 8392 13784
rect 7708 13744 7714 13756
rect 8386 13744 8392 13756
rect 8444 13744 8450 13796
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 9493 13787 9551 13793
rect 9493 13784 9505 13787
rect 9364 13756 9505 13784
rect 9364 13744 9370 13756
rect 9493 13753 9505 13756
rect 9539 13784 9551 13787
rect 9539 13756 9720 13784
rect 9539 13753 9551 13756
rect 9493 13747 9551 13753
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2130 13716 2136 13728
rect 1995 13688 2136 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2130 13676 2136 13688
rect 2188 13676 2194 13728
rect 2314 13716 2320 13728
rect 2275 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 8938 13676 8944 13728
rect 8996 13716 9002 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 8996 13688 9597 13716
rect 8996 13676 9002 13688
rect 9585 13685 9597 13688
rect 9631 13685 9643 13719
rect 9692 13716 9720 13756
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10505 13787 10563 13793
rect 10505 13784 10517 13787
rect 9824 13756 10517 13784
rect 9824 13744 9830 13756
rect 10505 13753 10517 13756
rect 10551 13753 10563 13787
rect 10505 13747 10563 13753
rect 11422 13744 11428 13796
rect 11480 13784 11486 13796
rect 11517 13787 11575 13793
rect 11517 13784 11529 13787
rect 11480 13756 11529 13784
rect 11480 13744 11486 13756
rect 11517 13753 11529 13756
rect 11563 13753 11575 13787
rect 11517 13747 11575 13753
rect 12986 13744 12992 13796
rect 13044 13784 13050 13796
rect 14182 13784 14188 13796
rect 13044 13756 14188 13784
rect 13044 13744 13050 13756
rect 14182 13744 14188 13756
rect 14240 13744 14246 13796
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 17313 13787 17371 13793
rect 17313 13784 17325 13787
rect 14700 13756 17325 13784
rect 14700 13744 14706 13756
rect 17313 13753 17325 13756
rect 17359 13753 17371 13787
rect 17313 13747 17371 13753
rect 18598 13744 18604 13796
rect 18656 13793 18662 13796
rect 18656 13787 18720 13793
rect 18656 13753 18674 13787
rect 18708 13784 18720 13787
rect 19334 13784 19340 13796
rect 18708 13756 19340 13784
rect 18708 13753 18720 13756
rect 18656 13747 18720 13753
rect 18656 13744 18662 13747
rect 19334 13744 19340 13756
rect 19392 13744 19398 13796
rect 19886 13744 19892 13796
rect 19944 13784 19950 13796
rect 20806 13784 20812 13796
rect 19944 13756 20812 13784
rect 19944 13744 19950 13756
rect 20806 13744 20812 13756
rect 20864 13744 20870 13796
rect 16482 13716 16488 13728
rect 9692 13688 16488 13716
rect 9585 13679 9643 13685
rect 16482 13676 16488 13688
rect 16540 13676 16546 13728
rect 16942 13676 16948 13728
rect 17000 13716 17006 13728
rect 17221 13719 17279 13725
rect 17221 13716 17233 13719
rect 17000 13688 17233 13716
rect 17000 13676 17006 13688
rect 17221 13685 17233 13688
rect 17267 13685 17279 13719
rect 17221 13679 17279 13685
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20441 13719 20499 13725
rect 20441 13716 20453 13719
rect 20220 13688 20453 13716
rect 20220 13676 20226 13688
rect 20441 13685 20453 13688
rect 20487 13685 20499 13719
rect 21266 13716 21272 13728
rect 21227 13688 21272 13716
rect 20441 13679 20499 13685
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 4338 13512 4344 13524
rect 4299 13484 4344 13512
rect 4338 13472 4344 13484
rect 4396 13472 4402 13524
rect 5074 13472 5080 13524
rect 5132 13512 5138 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 5132 13484 5181 13512
rect 5132 13472 5138 13484
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5718 13512 5724 13524
rect 5583 13484 5724 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 6236 13484 6377 13512
rect 6236 13472 6242 13484
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 6365 13475 6423 13481
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7377 13515 7435 13521
rect 7377 13512 7389 13515
rect 7156 13484 7389 13512
rect 7156 13472 7162 13484
rect 7377 13481 7389 13484
rect 7423 13481 7435 13515
rect 7377 13475 7435 13481
rect 7558 13472 7564 13524
rect 7616 13512 7622 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 7616 13484 7757 13512
rect 7616 13472 7622 13484
rect 7745 13481 7757 13484
rect 7791 13481 7803 13515
rect 7745 13475 7803 13481
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8389 13515 8447 13521
rect 8389 13512 8401 13515
rect 8352 13484 8401 13512
rect 8352 13472 8358 13484
rect 8389 13481 8401 13484
rect 8435 13481 8447 13515
rect 8846 13512 8852 13524
rect 8807 13484 8852 13512
rect 8389 13475 8447 13481
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 9214 13512 9220 13524
rect 8956 13484 9220 13512
rect 2498 13444 2504 13456
rect 2332 13416 2504 13444
rect 1581 13379 1639 13385
rect 1581 13345 1593 13379
rect 1627 13376 1639 13379
rect 2038 13376 2044 13388
rect 1627 13348 2044 13376
rect 1627 13345 1639 13348
rect 1581 13339 1639 13345
rect 2038 13336 2044 13348
rect 2096 13336 2102 13388
rect 2332 13385 2360 13416
rect 2498 13404 2504 13416
rect 2556 13444 2562 13456
rect 3050 13444 3056 13456
rect 2556 13416 3056 13444
rect 2556 13404 2562 13416
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13444 5687 13447
rect 5810 13444 5816 13456
rect 5675 13416 5816 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 5810 13404 5816 13416
rect 5868 13404 5874 13456
rect 6273 13447 6331 13453
rect 6273 13413 6285 13447
rect 6319 13444 6331 13447
rect 6454 13444 6460 13456
rect 6319 13416 6460 13444
rect 6319 13413 6331 13416
rect 6273 13407 6331 13413
rect 6454 13404 6460 13416
rect 6512 13444 6518 13456
rect 6733 13447 6791 13453
rect 6733 13444 6745 13447
rect 6512 13416 6745 13444
rect 6512 13404 6518 13416
rect 6733 13413 6745 13416
rect 6779 13444 6791 13447
rect 6822 13444 6828 13456
rect 6779 13416 6828 13444
rect 6779 13413 6791 13416
rect 6733 13407 6791 13413
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 2590 13385 2596 13388
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13345 2375 13379
rect 2584 13376 2596 13385
rect 2551 13348 2596 13376
rect 2317 13339 2375 13345
rect 2584 13339 2596 13348
rect 2590 13336 2596 13339
rect 2648 13336 2654 13388
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4709 13379 4767 13385
rect 4709 13376 4721 13379
rect 4212 13348 4721 13376
rect 4212 13336 4218 13348
rect 4709 13345 4721 13348
rect 4755 13345 4767 13379
rect 7576 13376 7604 13472
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 8757 13447 8815 13453
rect 8757 13444 8769 13447
rect 7708 13416 8769 13444
rect 7708 13404 7714 13416
rect 8757 13413 8769 13416
rect 8803 13413 8815 13447
rect 8757 13407 8815 13413
rect 8846 13376 8852 13388
rect 4709 13339 4767 13345
rect 5000 13348 5764 13376
rect 7576 13348 8852 13376
rect 5000 13320 5028 13348
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 1452 13280 1777 13308
rect 1452 13268 1458 13280
rect 1765 13277 1777 13280
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 4338 13308 4344 13320
rect 3936 13280 4344 13308
rect 3936 13268 3942 13280
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4798 13308 4804 13320
rect 4759 13280 4804 13308
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 4982 13308 4988 13320
rect 4943 13280 4988 13308
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 5736 13317 5764 13348
rect 8846 13336 8852 13348
rect 8904 13376 8910 13388
rect 8956 13376 8984 13484
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 10008 13484 10149 13512
rect 10008 13472 10014 13484
rect 10137 13481 10149 13484
rect 10183 13481 10195 13515
rect 10137 13475 10195 13481
rect 10594 13472 10600 13524
rect 10652 13512 10658 13524
rect 10778 13512 10784 13524
rect 10652 13484 10784 13512
rect 10652 13472 10658 13484
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11057 13515 11115 13521
rect 11057 13481 11069 13515
rect 11103 13512 11115 13515
rect 12066 13512 12072 13524
rect 11103 13484 12072 13512
rect 11103 13481 11115 13484
rect 11057 13475 11115 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 12161 13515 12219 13521
rect 12161 13481 12173 13515
rect 12207 13512 12219 13515
rect 12250 13512 12256 13524
rect 12207 13484 12256 13512
rect 12207 13481 12219 13484
rect 12161 13475 12219 13481
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 15289 13515 15347 13521
rect 12575 13484 14688 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 10318 13444 10324 13456
rect 8904 13348 8984 13376
rect 9048 13416 10324 13444
rect 8904 13336 8910 13348
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13277 5779 13311
rect 5721 13271 5779 13277
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6052 13280 6837 13308
rect 6052 13268 6058 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7374 13308 7380 13320
rect 7055 13280 7380 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 3694 13240 3700 13252
rect 3607 13212 3700 13240
rect 3694 13200 3700 13212
rect 3752 13240 3758 13252
rect 7024 13240 7052 13271
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 7834 13308 7840 13320
rect 7795 13280 7840 13308
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 3752 13212 7052 13240
rect 7392 13240 7420 13268
rect 7944 13240 7972 13271
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8260 13280 8953 13308
rect 8260 13268 8266 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9048 13240 9076 13416
rect 10318 13404 10324 13416
rect 10376 13404 10382 13456
rect 11422 13444 11428 13456
rect 11383 13416 11428 13444
rect 11422 13404 11428 13416
rect 11480 13404 11486 13456
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 11572 13416 11617 13444
rect 11572 13404 11578 13416
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9950 13376 9956 13388
rect 9456 13348 9956 13376
rect 9456 13336 9462 13348
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13376 10103 13379
rect 11146 13376 11152 13388
rect 10091 13348 11152 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 12544 13376 12572 13475
rect 13630 13453 13636 13456
rect 13624 13407 13636 13453
rect 13688 13444 13694 13456
rect 13688 13416 13724 13444
rect 13630 13404 13636 13407
rect 13688 13404 13694 13416
rect 11532 13348 12572 13376
rect 10318 13308 10324 13320
rect 10279 13280 10324 13308
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 11422 13308 11428 13320
rect 11112 13280 11428 13308
rect 11112 13268 11118 13280
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 7392 13212 7972 13240
rect 8036 13212 9076 13240
rect 3752 13200 3758 13212
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 8036 13172 8064 13212
rect 9398 13200 9404 13252
rect 9456 13240 9462 13252
rect 11532 13240 11560 13348
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 14660 13376 14688 13484
rect 15289 13481 15301 13515
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 15304 13444 15332 13475
rect 15654 13472 15660 13524
rect 15712 13512 15718 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15712 13484 16313 13512
rect 15712 13472 15718 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 17770 13472 17776 13524
rect 17828 13512 17834 13524
rect 18233 13515 18291 13521
rect 18233 13512 18245 13515
rect 17828 13484 18245 13512
rect 17828 13472 17834 13484
rect 18233 13481 18245 13484
rect 18279 13481 18291 13515
rect 18233 13475 18291 13481
rect 18785 13515 18843 13521
rect 18785 13481 18797 13515
rect 18831 13481 18843 13515
rect 19794 13512 19800 13524
rect 19755 13484 19800 13512
rect 18785 13475 18843 13481
rect 16574 13444 16580 13456
rect 15304 13416 16580 13444
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 18141 13447 18199 13453
rect 18141 13413 18153 13447
rect 18187 13444 18199 13447
rect 18800 13444 18828 13475
rect 19794 13472 19800 13484
rect 19852 13472 19858 13524
rect 18187 13416 18828 13444
rect 19153 13447 19211 13453
rect 18187 13413 18199 13416
rect 18141 13407 18199 13413
rect 19153 13413 19165 13447
rect 19199 13444 19211 13447
rect 19702 13444 19708 13456
rect 19199 13416 19708 13444
rect 19199 13413 19211 13416
rect 19153 13407 19211 13413
rect 19702 13404 19708 13416
rect 19760 13404 19766 13456
rect 20257 13447 20315 13453
rect 20257 13413 20269 13447
rect 20303 13444 20315 13447
rect 20346 13444 20352 13456
rect 20303 13416 20352 13444
rect 20303 13413 20315 13416
rect 20257 13407 20315 13413
rect 20346 13404 20352 13416
rect 20404 13404 20410 13456
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 12676 13348 14596 13376
rect 14660 13348 15669 13376
rect 12676 13336 12682 13348
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13277 12771 13311
rect 13354 13308 13360 13320
rect 13315 13280 13360 13308
rect 12713 13271 12771 13277
rect 12728 13240 12756 13271
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 9456 13212 11560 13240
rect 12084 13212 12756 13240
rect 9456 13200 9462 13212
rect 3568 13144 8064 13172
rect 3568 13132 3574 13144
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10502 13172 10508 13184
rect 10192 13144 10508 13172
rect 10192 13132 10198 13144
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 12084 13172 12112 13212
rect 11020 13144 12112 13172
rect 14568 13172 14596 13348
rect 15657 13345 15669 13348
rect 15703 13376 15715 13379
rect 16390 13376 16396 13388
rect 15703 13348 16396 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13376 16727 13379
rect 18046 13376 18052 13388
rect 16715 13348 18052 13376
rect 16715 13345 16727 13348
rect 16669 13339 16727 13345
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 19794 13336 19800 13388
rect 19852 13376 19858 13388
rect 20165 13379 20223 13385
rect 20165 13376 20177 13379
rect 19852 13348 20177 13376
rect 19852 13336 19858 13348
rect 20165 13345 20177 13348
rect 20211 13345 20223 13379
rect 20165 13339 20223 13345
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20864 13348 20913 13376
rect 20864 13336 20870 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 14826 13308 14832 13320
rect 14700 13280 14832 13308
rect 14700 13268 14706 13280
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 15344 13280 15761 13308
rect 15344 13268 15350 13280
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15749 13271 15807 13277
rect 15856 13280 15945 13308
rect 15856 13252 15884 13280
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13308 17003 13311
rect 17402 13308 17408 13320
rect 16991 13280 17408 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 14734 13240 14740 13252
rect 14695 13212 14740 13240
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 15378 13200 15384 13252
rect 15436 13240 15442 13252
rect 15654 13240 15660 13252
rect 15436 13212 15660 13240
rect 15436 13200 15442 13212
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 15838 13200 15844 13252
rect 15896 13200 15902 13252
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 16776 13240 16804 13271
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13308 18475 13311
rect 18690 13308 18696 13320
rect 18463 13280 18696 13308
rect 18463 13277 18475 13280
rect 18417 13271 18475 13277
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 18840 13280 19257 13308
rect 18840 13268 18846 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 20438 13308 20444 13320
rect 19392 13280 19437 13308
rect 20399 13280 20444 13308
rect 19392 13268 19398 13280
rect 20438 13268 20444 13280
rect 20496 13308 20502 13320
rect 20496 13280 20576 13308
rect 20496 13268 20502 13280
rect 16448 13212 16804 13240
rect 16448 13200 16454 13212
rect 17126 13200 17132 13252
rect 17184 13240 17190 13252
rect 17310 13240 17316 13252
rect 17184 13212 17316 13240
rect 17184 13200 17190 13212
rect 17310 13200 17316 13212
rect 17368 13200 17374 13252
rect 17773 13243 17831 13249
rect 17773 13209 17785 13243
rect 17819 13240 17831 13243
rect 18138 13240 18144 13252
rect 17819 13212 18144 13240
rect 17819 13209 17831 13212
rect 17773 13203 17831 13209
rect 18138 13200 18144 13212
rect 18196 13200 18202 13252
rect 19702 13200 19708 13252
rect 19760 13240 19766 13252
rect 20548 13240 20576 13280
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 20772 13280 21097 13308
rect 20772 13268 20778 13280
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 21266 13240 21272 13252
rect 19760 13212 20024 13240
rect 20548 13212 21272 13240
rect 19760 13200 19766 13212
rect 18690 13172 18696 13184
rect 14568 13144 18696 13172
rect 11020 13132 11026 13144
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 19886 13172 19892 13184
rect 19576 13144 19892 13172
rect 19576 13132 19582 13144
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 19996 13172 20024 13212
rect 21266 13200 21272 13212
rect 21324 13200 21330 13252
rect 20898 13172 20904 13184
rect 19996 13144 20904 13172
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1544 12940 2544 12968
rect 1544 12928 1550 12940
rect 2516 12900 2544 12940
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 2961 12971 3019 12977
rect 2961 12968 2973 12971
rect 2648 12940 2973 12968
rect 2648 12928 2654 12940
rect 2961 12937 2973 12940
rect 3007 12937 3019 12971
rect 4154 12968 4160 12980
rect 4115 12940 4160 12968
rect 2961 12931 3019 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4798 12928 4804 12980
rect 4856 12968 4862 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4856 12940 5181 12968
rect 4856 12928 4862 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 8205 12971 8263 12977
rect 5169 12931 5227 12937
rect 6748 12940 8156 12968
rect 4706 12900 4712 12912
rect 2516 12872 4712 12900
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 4985 12903 5043 12909
rect 4985 12869 4997 12903
rect 5031 12900 5043 12903
rect 5031 12872 6224 12900
rect 5031 12869 5043 12872
rect 4985 12863 5043 12869
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 3200 12804 3433 12832
rect 3200 12792 3206 12804
rect 3421 12801 3433 12804
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3694 12792 3700 12844
rect 3752 12832 3758 12844
rect 4062 12832 4068 12844
rect 3752 12804 4068 12832
rect 3752 12792 3758 12804
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12832 4859 12835
rect 5534 12832 5540 12844
rect 4847 12804 5540 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 5534 12792 5540 12804
rect 5592 12832 5598 12844
rect 6196 12841 6224 12872
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5592 12804 5733 12832
rect 5592 12792 5598 12804
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12801 6239 12835
rect 6181 12795 6239 12801
rect 1578 12764 1584 12776
rect 1539 12736 1584 12764
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 2130 12724 2136 12776
rect 2188 12764 2194 12776
rect 3237 12767 3295 12773
rect 3237 12764 3249 12767
rect 2188 12736 3249 12764
rect 2188 12724 2194 12736
rect 3237 12733 3249 12736
rect 3283 12733 3295 12767
rect 3237 12727 3295 12733
rect 3786 12724 3792 12776
rect 3844 12764 3850 12776
rect 5258 12764 5264 12776
rect 3844 12736 5264 12764
rect 3844 12724 3850 12736
rect 5258 12724 5264 12736
rect 5316 12764 5322 12776
rect 5629 12767 5687 12773
rect 5316 12736 5580 12764
rect 5316 12724 5322 12736
rect 1848 12699 1906 12705
rect 1848 12665 1860 12699
rect 1894 12696 1906 12699
rect 2038 12696 2044 12708
rect 1894 12668 2044 12696
rect 1894 12665 1906 12668
rect 1848 12659 1906 12665
rect 2038 12656 2044 12668
rect 2096 12656 2102 12708
rect 5552 12705 5580 12736
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 6748 12764 6776 12940
rect 8128 12832 8156 12940
rect 8205 12937 8217 12971
rect 8251 12968 8263 12971
rect 8478 12968 8484 12980
rect 8251 12940 8484 12968
rect 8251 12937 8263 12940
rect 8205 12931 8263 12937
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10137 12971 10195 12977
rect 10137 12968 10149 12971
rect 10100 12940 10149 12968
rect 10100 12928 10106 12940
rect 10137 12937 10149 12940
rect 10183 12937 10195 12971
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 10137 12931 10195 12937
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11756 12940 12020 12968
rect 11756 12928 11762 12940
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 11992 12900 12020 12940
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12618 12968 12624 12980
rect 12124 12940 12624 12968
rect 12124 12928 12130 12940
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 14458 12968 14464 12980
rect 13771 12940 14464 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 15286 12968 15292 12980
rect 15247 12940 15292 12968
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 17034 12968 17040 12980
rect 15856 12940 17040 12968
rect 12158 12900 12164 12912
rect 9640 12872 11744 12900
rect 11992 12872 12164 12900
rect 9640 12860 9646 12872
rect 10318 12832 10324 12844
rect 8128 12804 8616 12832
rect 5675 12736 6776 12764
rect 6825 12767 6883 12773
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7374 12764 7380 12776
rect 6871 12736 7380 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7374 12724 7380 12736
rect 7432 12764 7438 12776
rect 8386 12764 8392 12776
rect 7432 12736 8392 12764
rect 7432 12724 7438 12736
rect 8386 12724 8392 12736
rect 8444 12764 8450 12776
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 8444 12736 8493 12764
rect 8444 12724 8450 12736
rect 8481 12733 8493 12736
rect 8527 12733 8539 12767
rect 8588 12764 8616 12804
rect 9876 12804 10324 12832
rect 9674 12764 9680 12776
rect 8588 12736 9680 12764
rect 8481 12727 8539 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12696 4583 12699
rect 4985 12699 5043 12705
rect 4985 12696 4997 12699
rect 4571 12668 4997 12696
rect 4571 12665 4583 12668
rect 4525 12659 4583 12665
rect 4985 12665 4997 12668
rect 5031 12665 5043 12699
rect 4985 12659 5043 12665
rect 5537 12699 5595 12705
rect 5537 12665 5549 12699
rect 5583 12665 5595 12699
rect 5537 12659 5595 12665
rect 7092 12699 7150 12705
rect 7092 12665 7104 12699
rect 7138 12665 7150 12699
rect 7092 12659 7150 12665
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 3108 12600 4629 12628
rect 3108 12588 3114 12600
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 7107 12628 7135 12659
rect 7834 12656 7840 12708
rect 7892 12696 7898 12708
rect 8294 12696 8300 12708
rect 7892 12668 8300 12696
rect 7892 12656 7898 12668
rect 8294 12656 8300 12668
rect 8352 12696 8358 12708
rect 8570 12696 8576 12708
rect 8352 12668 8576 12696
rect 8352 12656 8358 12668
rect 8570 12656 8576 12668
rect 8628 12656 8634 12708
rect 8748 12699 8806 12705
rect 8748 12665 8760 12699
rect 8794 12696 8806 12699
rect 9214 12696 9220 12708
rect 8794 12668 9220 12696
rect 8794 12665 8806 12668
rect 8748 12659 8806 12665
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 7558 12628 7564 12640
rect 7107 12600 7564 12628
rect 4617 12591 4675 12597
rect 7558 12588 7564 12600
rect 7616 12628 7622 12640
rect 9876 12637 9904 12804
rect 10318 12792 10324 12804
rect 10376 12832 10382 12844
rect 11716 12841 11744 12872
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 12894 12900 12900 12912
rect 12452 12872 12900 12900
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10376 12804 10701 12832
rect 10376 12792 10382 12804
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 11882 12764 11888 12776
rect 10520 12736 11888 12764
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 7616 12600 9873 12628
rect 7616 12588 7622 12600
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10520 12637 10548 12736
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12696 11575 12699
rect 12452 12696 12480 12872
rect 12894 12860 12900 12872
rect 12952 12860 12958 12912
rect 13262 12860 13268 12912
rect 13320 12900 13326 12912
rect 13449 12903 13507 12909
rect 13449 12900 13461 12903
rect 13320 12872 13461 12900
rect 13320 12860 13326 12872
rect 13449 12869 13461 12872
rect 13495 12900 13507 12903
rect 14642 12900 14648 12912
rect 13495 12872 14648 12900
rect 13495 12869 13507 12872
rect 13449 12863 13507 12869
rect 14642 12860 14648 12872
rect 14700 12860 14706 12912
rect 15856 12900 15884 12940
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 17678 12968 17684 12980
rect 17639 12940 17684 12968
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 19518 12968 19524 12980
rect 17788 12940 19524 12968
rect 15764 12872 15884 12900
rect 12986 12832 12992 12844
rect 12947 12804 12992 12832
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 14056 12804 14197 12832
rect 14056 12792 14062 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 14734 12832 14740 12844
rect 14415 12804 14740 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 15764 12841 15792 12872
rect 17586 12860 17592 12912
rect 17644 12900 17650 12912
rect 17788 12900 17816 12940
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 19886 12968 19892 12980
rect 19751 12940 19892 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19886 12928 19892 12940
rect 19944 12928 19950 12980
rect 17644 12872 17816 12900
rect 18417 12903 18475 12909
rect 17644 12860 17650 12872
rect 18417 12869 18429 12903
rect 18463 12900 18475 12903
rect 20070 12900 20076 12912
rect 18463 12872 20076 12900
rect 18463 12869 18475 12872
rect 18417 12863 18475 12869
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 20438 12900 20444 12912
rect 20364 12872 20444 12900
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12801 15807 12835
rect 15930 12832 15936 12844
rect 15891 12804 15936 12832
rect 15749 12795 15807 12801
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 16298 12832 16304 12844
rect 16259 12804 16304 12832
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 18506 12832 18512 12844
rect 17368 12804 18512 12832
rect 17368 12792 17374 12804
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 19061 12835 19119 12841
rect 18616 12804 19012 12832
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 12584 12736 13645 12764
rect 12584 12724 12590 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 13872 12736 14105 12764
rect 13872 12724 13878 12736
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 18616 12764 18644 12804
rect 14516 12736 18644 12764
rect 14516 12724 14522 12736
rect 18874 12724 18880 12776
rect 18932 12724 18938 12776
rect 18984 12764 19012 12804
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 19150 12832 19156 12844
rect 19107 12804 19156 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 19150 12792 19156 12804
rect 19208 12832 19214 12844
rect 19334 12832 19340 12844
rect 19208 12804 19340 12832
rect 19208 12792 19214 12804
rect 19334 12792 19340 12804
rect 19392 12792 19398 12844
rect 20364 12841 20392 12872
rect 20438 12860 20444 12872
rect 20496 12860 20502 12912
rect 20349 12835 20407 12841
rect 19444 12804 20300 12832
rect 19444 12764 19472 12804
rect 18984 12736 19472 12764
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 20165 12767 20223 12773
rect 20165 12764 20177 12767
rect 19576 12736 20177 12764
rect 19576 12724 19582 12736
rect 20165 12733 20177 12736
rect 20211 12733 20223 12767
rect 20272 12764 20300 12804
rect 20349 12801 20361 12835
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 20438 12764 20444 12776
rect 20272 12736 20444 12764
rect 20165 12727 20223 12733
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 20717 12767 20775 12773
rect 20717 12733 20729 12767
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 11563 12668 12480 12696
rect 12805 12699 12863 12705
rect 11563 12665 11575 12668
rect 11517 12659 11575 12665
rect 12805 12665 12817 12699
rect 12851 12696 12863 12699
rect 12851 12668 13676 12696
rect 12851 12665 12863 12668
rect 12805 12659 12863 12665
rect 13648 12640 13676 12668
rect 14274 12656 14280 12708
rect 14332 12696 14338 12708
rect 14737 12699 14795 12705
rect 14737 12696 14749 12699
rect 14332 12668 14749 12696
rect 14332 12656 14338 12668
rect 14737 12665 14749 12668
rect 14783 12665 14795 12699
rect 14737 12659 14795 12665
rect 16568 12699 16626 12705
rect 16568 12665 16580 12699
rect 16614 12696 16626 12699
rect 17310 12696 17316 12708
rect 16614 12668 17316 12696
rect 16614 12665 16626 12668
rect 16568 12659 16626 12665
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 18785 12699 18843 12705
rect 18785 12696 18797 12699
rect 17828 12668 18797 12696
rect 17828 12656 17834 12668
rect 18785 12665 18797 12668
rect 18831 12665 18843 12699
rect 18892 12696 18920 12724
rect 18892 12668 19196 12696
rect 18785 12659 18843 12665
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 10008 12600 10517 12628
rect 10008 12588 10014 12600
rect 10505 12597 10517 12600
rect 10551 12597 10563 12631
rect 10505 12591 10563 12597
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 10652 12600 10697 12628
rect 10652 12588 10658 12600
rect 10962 12588 10968 12640
rect 11020 12628 11026 12640
rect 11238 12628 11244 12640
rect 11020 12600 11244 12628
rect 11020 12588 11026 12600
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 11609 12631 11667 12637
rect 11609 12597 11621 12631
rect 11655 12628 11667 12631
rect 11974 12628 11980 12640
rect 11655 12600 11980 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12894 12628 12900 12640
rect 12492 12600 12537 12628
rect 12855 12600 12900 12628
rect 12492 12588 12498 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13630 12588 13636 12640
rect 13688 12588 13694 12640
rect 15378 12588 15384 12640
rect 15436 12628 15442 12640
rect 15657 12631 15715 12637
rect 15657 12628 15669 12631
rect 15436 12600 15669 12628
rect 15436 12588 15442 12600
rect 15657 12597 15669 12600
rect 15703 12597 15715 12631
rect 15657 12591 15715 12597
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 18138 12628 18144 12640
rect 16816 12600 18144 12628
rect 16816 12588 16822 12600
rect 18138 12588 18144 12600
rect 18196 12628 18202 12640
rect 18690 12628 18696 12640
rect 18196 12600 18696 12628
rect 18196 12588 18202 12600
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 19168 12628 19196 12668
rect 19242 12656 19248 12708
rect 19300 12696 19306 12708
rect 19613 12699 19671 12705
rect 19613 12696 19625 12699
rect 19300 12668 19625 12696
rect 19300 12656 19306 12668
rect 19613 12665 19625 12668
rect 19659 12696 19671 12699
rect 20073 12699 20131 12705
rect 20073 12696 20085 12699
rect 19659 12668 20085 12696
rect 19659 12665 19671 12668
rect 19613 12659 19671 12665
rect 20073 12665 20085 12668
rect 20119 12665 20131 12699
rect 20073 12659 20131 12665
rect 20732 12628 20760 12727
rect 20993 12699 21051 12705
rect 20993 12665 21005 12699
rect 21039 12696 21051 12699
rect 21082 12696 21088 12708
rect 21039 12668 21088 12696
rect 21039 12665 21051 12668
rect 20993 12659 21051 12665
rect 21082 12656 21088 12668
rect 21140 12656 21146 12708
rect 18932 12600 18977 12628
rect 19168 12600 20760 12628
rect 18932 12588 18938 12600
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 3602 12424 3608 12436
rect 3563 12396 3608 12424
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 4065 12427 4123 12433
rect 4065 12393 4077 12427
rect 4111 12393 4123 12427
rect 4065 12387 4123 12393
rect 2032 12359 2090 12365
rect 2032 12325 2044 12359
rect 2078 12356 2090 12359
rect 2222 12356 2228 12368
rect 2078 12328 2228 12356
rect 2078 12325 2090 12328
rect 2032 12319 2090 12325
rect 2222 12316 2228 12328
rect 2280 12316 2286 12368
rect 2958 12316 2964 12368
rect 3016 12356 3022 12368
rect 4080 12356 4108 12387
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 8202 12424 8208 12436
rect 5132 12396 5177 12424
rect 8163 12396 8208 12424
rect 5132 12384 5138 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8588 12396 13584 12424
rect 3016 12328 4108 12356
rect 7092 12359 7150 12365
rect 3016 12316 3022 12328
rect 7092 12325 7104 12359
rect 7138 12356 7150 12359
rect 8478 12356 8484 12368
rect 7138 12328 8484 12356
rect 7138 12325 7150 12328
rect 7092 12319 7150 12325
rect 8478 12316 8484 12328
rect 8536 12316 8542 12368
rect 1578 12248 1584 12300
rect 1636 12288 1642 12300
rect 1765 12291 1823 12297
rect 1765 12288 1777 12291
rect 1636 12260 1777 12288
rect 1636 12248 1642 12260
rect 1765 12257 1777 12260
rect 1811 12288 1823 12291
rect 2498 12288 2504 12300
rect 1811 12260 2504 12288
rect 1811 12257 1823 12260
rect 1765 12251 1823 12257
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3200 12260 3433 12288
rect 3200 12248 3206 12260
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 4120 12260 4445 12288
rect 4120 12248 4126 12260
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 5258 12288 5264 12300
rect 4571 12260 5264 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5442 12288 5448 12300
rect 5403 12260 5448 12288
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 6825 12291 6883 12297
rect 6825 12288 6837 12291
rect 6420 12260 6837 12288
rect 6420 12248 6426 12260
rect 6825 12257 6837 12260
rect 6871 12257 6883 12291
rect 8588 12288 8616 12396
rect 11977 12359 12035 12365
rect 10520 12328 11928 12356
rect 8938 12288 8944 12300
rect 6825 12251 6883 12257
rect 6932 12260 8616 12288
rect 8851 12260 8944 12288
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 3160 12192 4629 12220
rect 3160 12161 3188 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 4982 12180 4988 12232
rect 5040 12220 5046 12232
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 5040 12192 5549 12220
rect 5040 12180 5046 12192
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 6932 12220 6960 12260
rect 8938 12248 8944 12260
rect 8996 12288 9002 12300
rect 9122 12288 9128 12300
rect 8996 12260 9128 12288
rect 8996 12248 9002 12260
rect 9122 12248 9128 12260
rect 9180 12248 9186 12300
rect 5684 12192 5729 12220
rect 5828 12192 6960 12220
rect 5684 12180 5690 12192
rect 3145 12155 3203 12161
rect 3145 12121 3157 12155
rect 3191 12121 3203 12155
rect 3145 12115 3203 12121
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 3160 12084 3188 12115
rect 3878 12112 3884 12164
rect 3936 12152 3942 12164
rect 5828 12152 5856 12192
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 9033 12223 9091 12229
rect 9033 12220 9045 12223
rect 8628 12192 9045 12220
rect 8628 12180 8634 12192
rect 9033 12189 9045 12192
rect 9079 12189 9091 12223
rect 9214 12220 9220 12232
rect 9175 12192 9220 12220
rect 9033 12183 9091 12189
rect 9214 12180 9220 12192
rect 9272 12220 9278 12232
rect 9582 12220 9588 12232
rect 9272 12192 9588 12220
rect 9272 12180 9278 12192
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 10410 12220 10416 12232
rect 10323 12192 10416 12220
rect 10410 12180 10416 12192
rect 10468 12220 10474 12232
rect 10520 12220 10548 12328
rect 10680 12291 10738 12297
rect 10680 12257 10692 12291
rect 10726 12288 10738 12291
rect 11146 12288 11152 12300
rect 10726 12260 11152 12288
rect 10726 12257 10738 12260
rect 10680 12251 10738 12257
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 11900 12288 11928 12328
rect 11977 12325 11989 12359
rect 12023 12356 12035 12359
rect 12314 12359 12372 12365
rect 12314 12356 12326 12359
rect 12023 12328 12326 12356
rect 12023 12325 12035 12328
rect 11977 12319 12035 12325
rect 12314 12325 12326 12328
rect 12360 12356 12372 12359
rect 12986 12356 12992 12368
rect 12360 12328 12992 12356
rect 12360 12325 12372 12328
rect 12314 12319 12372 12325
rect 12986 12316 12992 12328
rect 13044 12316 13050 12368
rect 13556 12356 13584 12396
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13688 12396 13737 12424
rect 13688 12384 13694 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 13725 12387 13783 12393
rect 17310 12384 17316 12436
rect 17368 12424 17374 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17368 12396 17509 12424
rect 17368 12384 17374 12396
rect 17497 12393 17509 12396
rect 17543 12424 17555 12427
rect 17862 12424 17868 12436
rect 17543 12396 17868 12424
rect 17543 12393 17555 12396
rect 17497 12387 17555 12393
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 19208 12396 19441 12424
rect 19208 12384 19214 12396
rect 19429 12393 19441 12396
rect 19475 12393 19487 12427
rect 19429 12387 19487 12393
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 20806 12424 20812 12436
rect 19567 12396 20812 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 14185 12359 14243 12365
rect 14185 12356 14197 12359
rect 13556 12328 14197 12356
rect 14185 12325 14197 12328
rect 14231 12356 14243 12359
rect 14366 12356 14372 12368
rect 14231 12328 14372 12356
rect 14231 12325 14243 12328
rect 14185 12319 14243 12325
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 15286 12316 15292 12368
rect 15344 12356 15350 12368
rect 15562 12356 15568 12368
rect 15344 12328 15568 12356
rect 15344 12316 15350 12328
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 16298 12356 16304 12368
rect 16132 12328 16304 12356
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11900 12260 12081 12288
rect 12069 12257 12081 12260
rect 12115 12288 12127 12291
rect 12158 12288 12164 12300
rect 12115 12260 12164 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 14093 12291 14151 12297
rect 14093 12288 14105 12291
rect 12676 12260 14105 12288
rect 12676 12248 12682 12260
rect 14093 12257 14105 12260
rect 14139 12257 14151 12291
rect 14093 12251 14151 12257
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15252 12260 15669 12288
rect 15252 12248 15258 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 14366 12220 14372 12232
rect 10468 12192 10548 12220
rect 14327 12192 14372 12220
rect 10468 12180 10474 12192
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 16132 12229 16160 12328
rect 16298 12316 16304 12328
rect 16356 12356 16362 12368
rect 16356 12328 16528 12356
rect 16356 12316 16362 12328
rect 16390 12297 16396 12300
rect 16384 12288 16396 12297
rect 16351 12260 16396 12288
rect 16384 12251 16396 12260
rect 16390 12248 16396 12251
rect 16448 12248 16454 12300
rect 16500 12288 16528 12328
rect 16574 12316 16580 12368
rect 16632 12356 16638 12368
rect 17126 12356 17132 12368
rect 16632 12328 17132 12356
rect 16632 12316 16638 12328
rect 17126 12316 17132 12328
rect 17184 12316 17190 12368
rect 17678 12316 17684 12368
rect 17736 12356 17742 12368
rect 18294 12359 18352 12365
rect 18294 12356 18306 12359
rect 17736 12328 18306 12356
rect 17736 12316 17742 12328
rect 18294 12325 18306 12328
rect 18340 12325 18352 12359
rect 19981 12359 20039 12365
rect 19981 12356 19993 12359
rect 18294 12319 18352 12325
rect 19720 12328 19993 12356
rect 17773 12291 17831 12297
rect 16500 12260 17172 12288
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12220 15439 12223
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 15427 12192 16129 12220
rect 15427 12189 15439 12192
rect 15381 12183 15439 12189
rect 16117 12189 16129 12192
rect 16163 12189 16175 12223
rect 17144 12220 17172 12260
rect 17773 12257 17785 12291
rect 17819 12288 17831 12291
rect 19242 12288 19248 12300
rect 17819 12260 19248 12288
rect 17819 12257 17831 12260
rect 17773 12251 17831 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19720 12288 19748 12328
rect 19981 12325 19993 12328
rect 20027 12325 20039 12359
rect 19981 12319 20039 12325
rect 19886 12288 19892 12300
rect 19392 12260 19748 12288
rect 19847 12260 19892 12288
rect 19392 12248 19398 12260
rect 19886 12248 19892 12260
rect 19944 12248 19950 12300
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 17144 12192 18061 12220
rect 16117 12183 16175 12189
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 18049 12183 18107 12189
rect 19352 12192 20085 12220
rect 9306 12152 9312 12164
rect 3936 12124 5856 12152
rect 8496 12124 9312 12152
rect 3936 12112 3942 12124
rect 2096 12056 3188 12084
rect 2096 12044 2102 12056
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 8496 12084 8524 12124
rect 9306 12112 9312 12124
rect 9364 12152 9370 12164
rect 10042 12152 10048 12164
rect 9364 12124 10048 12152
rect 9364 12112 9370 12124
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 11977 12155 12035 12161
rect 11977 12152 11989 12155
rect 11839 12124 11989 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 11977 12121 11989 12124
rect 12023 12121 12035 12155
rect 11977 12115 12035 12121
rect 13078 12112 13084 12164
rect 13136 12152 13142 12164
rect 13354 12152 13360 12164
rect 13136 12124 13360 12152
rect 13136 12112 13142 12124
rect 13354 12112 13360 12124
rect 13412 12112 13418 12164
rect 19242 12112 19248 12164
rect 19300 12152 19306 12164
rect 19352 12152 19380 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20990 12180 20996 12232
rect 21048 12220 21054 12232
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 21048 12192 21097 12220
rect 21048 12180 21054 12192
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 19300 12124 19380 12152
rect 19300 12112 19306 12124
rect 3476 12056 8524 12084
rect 8573 12087 8631 12093
rect 3476 12044 3482 12056
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 10594 12084 10600 12096
rect 8619 12056 10600 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 13446 12084 13452 12096
rect 13407 12056 13452 12084
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 15381 12087 15439 12093
rect 15381 12053 15393 12087
rect 15427 12084 15439 12087
rect 15470 12084 15476 12096
rect 15427 12056 15476 12084
rect 15427 12053 15439 12056
rect 15381 12047 15439 12053
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 17954 12084 17960 12096
rect 16448 12056 17960 12084
rect 16448 12044 16454 12056
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1397 11883 1455 11889
rect 1397 11849 1409 11883
rect 1443 11880 1455 11883
rect 2314 11880 2320 11892
rect 1443 11852 2320 11880
rect 1443 11849 1455 11852
rect 1397 11843 1455 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 6825 11883 6883 11889
rect 3568 11852 5948 11880
rect 3568 11840 3574 11852
rect 3789 11815 3847 11821
rect 3789 11781 3801 11815
rect 3835 11812 3847 11815
rect 4614 11812 4620 11824
rect 3835 11784 4620 11812
rect 3835 11781 3847 11784
rect 3789 11775 3847 11781
rect 2038 11744 2044 11756
rect 1999 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2409 11679 2467 11685
rect 2409 11645 2421 11679
rect 2455 11676 2467 11679
rect 2498 11676 2504 11688
rect 2455 11648 2504 11676
rect 2455 11645 2467 11648
rect 2409 11639 2467 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 2676 11611 2734 11617
rect 2676 11577 2688 11611
rect 2722 11608 2734 11611
rect 3602 11608 3608 11620
rect 2722 11580 3608 11608
rect 2722 11577 2734 11580
rect 2676 11571 2734 11577
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 1946 11540 1952 11552
rect 1903 11512 1952 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 3804 11540 3832 11775
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 5258 11812 5264 11824
rect 5219 11784 5264 11812
rect 5258 11772 5264 11784
rect 5316 11772 5322 11824
rect 5920 11812 5948 11852
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 7650 11880 7656 11892
rect 6871 11852 7656 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8478 11880 8484 11892
rect 7760 11852 8484 11880
rect 7374 11812 7380 11824
rect 5920 11784 7380 11812
rect 7374 11772 7380 11784
rect 7432 11772 7438 11824
rect 7760 11812 7788 11852
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 10502 11880 10508 11892
rect 8628 11852 10508 11880
rect 8628 11840 8634 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11698 11880 11704 11892
rect 10652 11852 11704 11880
rect 10652 11840 10658 11852
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 15470 11880 15476 11892
rect 14292 11852 15476 11880
rect 7484 11784 7788 11812
rect 9217 11815 9275 11821
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11744 4951 11747
rect 5626 11744 5632 11756
rect 4939 11716 5632 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 7484 11753 7512 11784
rect 9217 11781 9229 11815
rect 9263 11781 9275 11815
rect 9217 11775 9275 11781
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11713 7527 11747
rect 7834 11744 7840 11756
rect 7795 11716 7840 11744
rect 7469 11707 7527 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 9232 11744 9260 11775
rect 9490 11772 9496 11824
rect 9548 11812 9554 11824
rect 9548 11784 10272 11812
rect 9548 11772 9554 11784
rect 10134 11744 10140 11756
rect 9232 11716 10140 11744
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10244 11744 10272 11784
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 10689 11815 10747 11821
rect 10689 11812 10701 11815
rect 10376 11784 10701 11812
rect 10376 11772 10382 11784
rect 10689 11781 10701 11784
rect 10735 11781 10747 11815
rect 10689 11775 10747 11781
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 11974 11812 11980 11824
rect 11020 11784 11980 11812
rect 11020 11772 11026 11784
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 13817 11815 13875 11821
rect 13817 11781 13829 11815
rect 13863 11812 13875 11815
rect 14182 11812 14188 11824
rect 13863 11784 14188 11812
rect 13863 11781 13875 11784
rect 13817 11775 13875 11781
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 10244 11716 11253 11744
rect 11241 11713 11253 11716
rect 11287 11744 11299 11747
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11287 11716 12081 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 12158 11704 12164 11756
rect 12216 11744 12222 11756
rect 14292 11753 14320 11852
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 16758 11880 16764 11892
rect 16356 11852 16764 11880
rect 16356 11840 16362 11852
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 19794 11880 19800 11892
rect 16991 11852 19800 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 21269 11883 21327 11889
rect 21269 11849 21281 11883
rect 21315 11880 21327 11883
rect 21450 11880 21456 11892
rect 21315 11852 21456 11880
rect 21315 11849 21327 11852
rect 21269 11843 21327 11849
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 19061 11815 19119 11821
rect 19061 11812 19073 11815
rect 17420 11784 19073 11812
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 12216 11716 12449 11744
rect 12216 11704 12222 11716
rect 12437 11713 12449 11716
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16206 11744 16212 11756
rect 16080 11716 16212 11744
rect 16080 11704 16086 11716
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 16482 11744 16488 11756
rect 16443 11716 16488 11744
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 17420 11753 17448 11784
rect 19061 11781 19073 11784
rect 19107 11781 19119 11815
rect 19061 11775 19119 11781
rect 20438 11772 20444 11824
rect 20496 11812 20502 11824
rect 21542 11812 21548 11824
rect 20496 11784 21548 11812
rect 20496 11772 20502 11784
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11713 17463 11747
rect 17586 11744 17592 11756
rect 17547 11716 17592 11744
rect 17405 11707 17463 11713
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 18506 11704 18512 11756
rect 18564 11744 18570 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18564 11716 18613 11744
rect 18564 11704 18570 11716
rect 18601 11713 18613 11716
rect 18647 11744 18659 11747
rect 19242 11744 19248 11756
rect 18647 11716 19248 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 19242 11704 19248 11716
rect 19300 11744 19306 11756
rect 20548 11753 20576 11784
rect 21542 11772 21548 11784
rect 21600 11772 21606 11824
rect 19613 11747 19671 11753
rect 19613 11744 19625 11747
rect 19300 11716 19625 11744
rect 19300 11704 19306 11716
rect 19613 11713 19625 11716
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11713 20683 11747
rect 20625 11707 20683 11713
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4522 11676 4528 11688
rect 4304 11648 4528 11676
rect 4304 11636 4310 11648
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 4798 11676 4804 11688
rect 4755 11648 4804 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 10318 11676 10324 11688
rect 5767 11648 10324 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 10870 11676 10876 11688
rect 10744 11648 10876 11676
rect 10744 11636 10750 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 11020 11648 11069 11676
rect 11020 11636 11026 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11388 11648 11897 11676
rect 11388 11636 11394 11648
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 11977 11679 12035 11685
rect 11977 11645 11989 11679
rect 12023 11676 12035 11679
rect 12342 11676 12348 11688
rect 12023 11648 12348 11676
rect 12023 11645 12035 11648
rect 11977 11639 12035 11645
rect 5629 11611 5687 11617
rect 5629 11608 5641 11611
rect 4264 11580 5641 11608
rect 4264 11549 4292 11580
rect 5629 11577 5641 11580
rect 5675 11577 5687 11611
rect 5629 11571 5687 11577
rect 8104 11611 8162 11617
rect 8104 11577 8116 11611
rect 8150 11608 8162 11611
rect 8202 11608 8208 11620
rect 8150 11580 8208 11608
rect 8150 11577 8162 11580
rect 8104 11571 8162 11577
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 8662 11568 8668 11620
rect 8720 11608 8726 11620
rect 9030 11608 9036 11620
rect 8720 11580 9036 11608
rect 8720 11568 8726 11580
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 9953 11611 10011 11617
rect 9953 11577 9965 11611
rect 9999 11608 10011 11611
rect 11790 11608 11796 11620
rect 9999 11580 11796 11608
rect 9999 11577 10011 11580
rect 9953 11571 10011 11577
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 2280 11512 3832 11540
rect 4249 11543 4307 11549
rect 2280 11500 2286 11512
rect 4249 11509 4261 11543
rect 4295 11509 4307 11543
rect 4249 11503 4307 11509
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4580 11512 4629 11540
rect 4580 11500 4586 11512
rect 4617 11509 4629 11512
rect 4663 11540 4675 11543
rect 5258 11540 5264 11552
rect 4663 11512 5264 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 6273 11543 6331 11549
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6822 11540 6828 11552
rect 6319 11512 6828 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7190 11540 7196 11552
rect 7151 11512 7196 11540
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 9493 11543 9551 11549
rect 7340 11512 7385 11540
rect 7340 11500 7346 11512
rect 9493 11509 9505 11543
rect 9539 11540 9551 11543
rect 9766 11540 9772 11552
rect 9539 11512 9772 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10778 11540 10784 11552
rect 9907 11512 10784 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 10928 11512 11161 11540
rect 10928 11500 10934 11512
rect 11149 11509 11161 11512
rect 11195 11509 11207 11543
rect 11514 11540 11520 11552
rect 11475 11512 11520 11540
rect 11149 11503 11207 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11992 11540 12020 11639
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 12710 11685 12716 11688
rect 12704 11676 12716 11685
rect 12623 11648 12716 11676
rect 12704 11639 12716 11648
rect 12768 11676 12774 11688
rect 13446 11676 13452 11688
rect 12768 11648 13452 11676
rect 12710 11636 12716 11639
rect 12768 11636 12774 11648
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 14550 11685 14556 11688
rect 14544 11639 14556 11685
rect 14608 11676 14614 11688
rect 16298 11676 16304 11688
rect 14608 11648 14644 11676
rect 16259 11648 16304 11676
rect 14550 11636 14556 11639
rect 14608 11636 14614 11648
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 18046 11676 18052 11688
rect 16448 11648 18052 11676
rect 16448 11636 16454 11648
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18690 11636 18696 11688
rect 18748 11676 18754 11688
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 18748 11648 19441 11676
rect 18748 11636 18754 11648
rect 19429 11645 19441 11648
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 19521 11679 19579 11685
rect 19521 11645 19533 11679
rect 19567 11676 19579 11679
rect 19702 11676 19708 11688
rect 19567 11648 19708 11676
rect 19567 11645 19579 11648
rect 19521 11639 19579 11645
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 16666 11608 16672 11620
rect 12216 11580 16672 11608
rect 12216 11568 12222 11580
rect 16666 11568 16672 11580
rect 16724 11568 16730 11620
rect 17313 11611 17371 11617
rect 17313 11577 17325 11611
rect 17359 11608 17371 11611
rect 18509 11611 18567 11617
rect 17359 11580 18092 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 11664 11512 12020 11540
rect 15657 11543 15715 11549
rect 11664 11500 11670 11512
rect 15657 11509 15669 11543
rect 15703 11540 15715 11543
rect 15746 11540 15752 11552
rect 15703 11512 15752 11540
rect 15703 11509 15715 11512
rect 15657 11503 15715 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 18064 11549 18092 11580
rect 18509 11577 18521 11611
rect 18555 11608 18567 11611
rect 18598 11608 18604 11620
rect 18555 11580 18604 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 18598 11568 18604 11580
rect 18656 11608 18662 11620
rect 18877 11611 18935 11617
rect 18877 11608 18889 11611
rect 18656 11580 18889 11608
rect 18656 11568 18662 11580
rect 18877 11577 18889 11580
rect 18923 11577 18935 11611
rect 20640 11608 20668 11707
rect 21082 11676 21088 11688
rect 21043 11648 21088 11676
rect 21082 11636 21088 11648
rect 21140 11636 21146 11688
rect 18877 11571 18935 11577
rect 18984 11580 20668 11608
rect 18049 11543 18107 11549
rect 18049 11509 18061 11543
rect 18095 11509 18107 11543
rect 18414 11540 18420 11552
rect 18375 11512 18420 11540
rect 18049 11503 18107 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 18984 11540 19012 11580
rect 18748 11512 19012 11540
rect 18748 11500 18754 11512
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 20073 11543 20131 11549
rect 20073 11540 20085 11543
rect 19760 11512 20085 11540
rect 19760 11500 19766 11512
rect 20073 11509 20085 11512
rect 20119 11509 20131 11543
rect 20438 11540 20444 11552
rect 20399 11512 20444 11540
rect 20073 11503 20131 11509
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2363 11308 2973 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 2961 11299 3019 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 5166 11336 5172 11348
rect 4479 11308 5172 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5776 11308 5825 11336
rect 5776 11296 5782 11308
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 5813 11299 5871 11305
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 7190 11336 7196 11348
rect 6871 11308 7196 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 7285 11339 7343 11345
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 7374 11336 7380 11348
rect 7331 11308 7380 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 11514 11336 11520 11348
rect 7699 11308 11520 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 12158 11336 12164 11348
rect 11900 11308 12164 11336
rect 2409 11271 2467 11277
rect 2409 11237 2421 11271
rect 2455 11268 2467 11271
rect 5074 11268 5080 11280
rect 2455 11240 5080 11268
rect 2455 11237 2467 11240
rect 2409 11231 2467 11237
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 6273 11271 6331 11277
rect 6273 11237 6285 11271
rect 6319 11268 6331 11271
rect 8202 11268 8208 11280
rect 6319 11240 8208 11268
rect 6319 11237 6331 11240
rect 6273 11231 6331 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 8941 11271 8999 11277
rect 8941 11237 8953 11271
rect 8987 11268 8999 11271
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 8987 11240 9413 11268
rect 8987 11237 8999 11240
rect 8941 11231 8999 11237
rect 9401 11237 9413 11240
rect 9447 11237 9459 11271
rect 9401 11231 9459 11237
rect 9582 11228 9588 11280
rect 9640 11268 9646 11280
rect 10042 11268 10048 11280
rect 9640 11240 10048 11268
rect 9640 11228 9646 11240
rect 10042 11228 10048 11240
rect 10100 11268 10106 11280
rect 11900 11268 11928 11308
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 12492 11308 12541 11336
rect 12492 11296 12498 11308
rect 12529 11305 12541 11308
rect 12575 11305 12587 11339
rect 12529 11299 12587 11305
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 12860 11308 14565 11336
rect 12860 11296 12866 11308
rect 14553 11305 14565 11308
rect 14599 11305 14611 11339
rect 14553 11299 14611 11305
rect 14645 11339 14703 11345
rect 14645 11305 14657 11339
rect 14691 11336 14703 11339
rect 18414 11336 18420 11348
rect 14691 11308 18420 11336
rect 14691 11305 14703 11308
rect 14645 11299 14703 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 18969 11339 19027 11345
rect 18969 11305 18981 11339
rect 19015 11305 19027 11339
rect 19702 11336 19708 11348
rect 19663 11308 19708 11336
rect 18969 11299 19027 11305
rect 10100 11240 11928 11268
rect 10100 11228 10106 11240
rect 11974 11228 11980 11280
rect 12032 11268 12038 11280
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 12032 11240 15669 11268
rect 12032 11228 12038 11240
rect 15657 11237 15669 11240
rect 15703 11237 15715 11271
rect 15657 11231 15715 11237
rect 17770 11228 17776 11280
rect 17828 11277 17834 11280
rect 17828 11271 17892 11277
rect 17828 11237 17846 11271
rect 17880 11237 17892 11271
rect 17828 11231 17892 11237
rect 17828 11228 17834 11231
rect 17954 11228 17960 11280
rect 18012 11268 18018 11280
rect 18984 11268 19012 11299
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 20441 11339 20499 11345
rect 20441 11305 20453 11339
rect 20487 11336 20499 11339
rect 20622 11336 20628 11348
rect 20487 11308 20628 11336
rect 20487 11305 20499 11308
rect 20441 11299 20499 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 21174 11268 21180 11280
rect 18012 11240 19012 11268
rect 21135 11240 21180 11268
rect 18012 11228 18018 11240
rect 21174 11228 21180 11240
rect 21232 11228 21238 11280
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 2682 11160 2688 11212
rect 2740 11200 2746 11212
rect 3050 11200 3056 11212
rect 2740 11172 3056 11200
rect 2740 11160 2746 11172
rect 3050 11160 3056 11172
rect 3108 11200 3114 11212
rect 3329 11203 3387 11209
rect 3329 11200 3341 11203
rect 3108 11172 3341 11200
rect 3108 11160 3114 11172
rect 3329 11169 3341 11172
rect 3375 11169 3387 11203
rect 5626 11200 5632 11212
rect 3329 11163 3387 11169
rect 3620 11172 5632 11200
rect 3620 11144 3648 11172
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 6880 11172 7205 11200
rect 6880 11160 6886 11172
rect 7193 11169 7205 11172
rect 7239 11169 7251 11203
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 7193 11163 7251 11169
rect 7300 11172 7665 11200
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2280 11104 2513 11132
rect 2280 11092 2286 11104
rect 2501 11101 2513 11104
rect 2547 11101 2559 11135
rect 3418 11132 3424 11144
rect 3379 11104 3424 11132
rect 2501 11095 2559 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3602 11132 3608 11144
rect 3515 11104 3608 11132
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 2774 11064 2780 11076
rect 1627 11036 2780 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4540 11064 4568 11095
rect 4614 11092 4620 11144
rect 4672 11132 4678 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 4672 11104 4721 11132
rect 4672 11092 4678 11104
rect 4709 11101 4721 11104
rect 4755 11132 4767 11135
rect 5810 11132 5816 11144
rect 4755 11104 5816 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 7300 11132 7328 11172
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 7653 11163 7711 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 9033 11203 9091 11209
rect 9033 11169 9045 11203
rect 9079 11200 9091 11203
rect 9674 11200 9680 11212
rect 9079 11172 9680 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 6420 11104 6465 11132
rect 6564 11104 7328 11132
rect 7469 11135 7527 11141
rect 6420 11092 6426 11104
rect 6564 11064 6592 11104
rect 7469 11101 7481 11135
rect 7515 11132 7527 11135
rect 7558 11132 7564 11144
rect 7515 11104 7564 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 4120 11036 4200 11064
rect 4540 11036 6592 11064
rect 4120 11024 4126 11036
rect 4172 10996 4200 11036
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7834 11064 7840 11076
rect 7064 11036 7840 11064
rect 7064 11024 7070 11036
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8036 11064 8064 11163
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10318 11200 10324 11212
rect 10279 11172 10324 11200
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 12526 11200 12532 11212
rect 11624 11172 12532 11200
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9582 11132 9588 11144
rect 9263 11104 9588 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10502 11132 10508 11144
rect 10284 11104 10508 11132
rect 10284 11092 10290 11104
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 11624 11073 11652 11172
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 12860 11172 13001 11200
rect 12860 11160 12866 11172
rect 12989 11169 13001 11172
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 13256 11203 13314 11209
rect 13256 11169 13268 11203
rect 13302 11200 13314 11203
rect 13998 11200 14004 11212
rect 13302 11172 14004 11200
rect 13302 11169 13314 11172
rect 13256 11163 13314 11169
rect 13998 11160 14004 11172
rect 14056 11200 14062 11212
rect 14182 11200 14188 11212
rect 14056 11172 14188 11200
rect 14056 11160 14062 11172
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 14550 11200 14556 11212
rect 14463 11172 14556 11200
rect 14550 11160 14556 11172
rect 14608 11200 14614 11212
rect 15749 11203 15807 11209
rect 15749 11200 15761 11203
rect 14608 11172 15761 11200
rect 14608 11160 14614 11172
rect 15749 11169 15761 11172
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 17126 11200 17132 11212
rect 16715 11172 17132 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 19150 11160 19156 11212
rect 19208 11200 19214 11212
rect 19334 11200 19340 11212
rect 19208 11172 19340 11200
rect 19208 11160 19214 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19613 11203 19671 11209
rect 19613 11169 19625 11203
rect 19659 11200 19671 11203
rect 19702 11200 19708 11212
rect 19659 11172 19708 11200
rect 19659 11169 19671 11172
rect 19613 11163 19671 11169
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 20257 11203 20315 11209
rect 20257 11169 20269 11203
rect 20303 11200 20315 11203
rect 20714 11200 20720 11212
rect 20303 11172 20720 11200
rect 20303 11169 20315 11172
rect 20257 11163 20315 11169
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 20901 11203 20959 11209
rect 20901 11169 20913 11203
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 12492 11104 12633 11132
rect 12492 11092 12498 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 15838 11132 15844 11144
rect 12768 11104 12813 11132
rect 15799 11104 15844 11132
rect 12768 11092 12774 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 16758 11132 16764 11144
rect 16719 11104 16764 11132
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16853 11135 16911 11141
rect 16853 11101 16865 11135
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11101 17647 11135
rect 17589 11095 17647 11101
rect 11609 11067 11667 11073
rect 11609 11064 11621 11067
rect 8036 11036 11621 11064
rect 11609 11033 11621 11036
rect 11655 11033 11667 11067
rect 11609 11027 11667 11033
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 14369 11067 14427 11073
rect 11848 11036 13032 11064
rect 11848 11024 11854 11036
rect 4890 10996 4896 11008
rect 4172 10968 4896 10996
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 6270 10956 6276 11008
rect 6328 10996 6334 11008
rect 7466 10996 7472 11008
rect 6328 10968 7472 10996
rect 6328 10956 6334 10968
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 8570 10996 8576 11008
rect 8531 10968 8576 10996
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 9401 10999 9459 11005
rect 9401 10965 9413 10999
rect 9447 10996 9459 10999
rect 10042 10996 10048 11008
rect 9447 10968 10048 10996
rect 9447 10965 9459 10968
rect 9401 10959 9459 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 12158 10996 12164 11008
rect 12119 10968 12164 10996
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 13004 10996 13032 11036
rect 14369 11033 14381 11067
rect 14415 11064 14427 11067
rect 14458 11064 14464 11076
rect 14415 11036 14464 11064
rect 14415 11033 14427 11036
rect 14369 11027 14427 11033
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 15289 11067 15347 11073
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 16666 11064 16672 11076
rect 15335 11036 16672 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 13906 10996 13912 11008
rect 13004 10968 13912 10996
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 14240 10968 16313 10996
rect 14240 10956 14246 10968
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 16301 10959 16359 10965
rect 16482 10956 16488 11008
rect 16540 10996 16546 11008
rect 16868 10996 16896 11095
rect 16540 10968 16896 10996
rect 17604 10996 17632 11095
rect 19242 11092 19248 11144
rect 19300 11132 19306 11144
rect 19797 11135 19855 11141
rect 19797 11132 19809 11135
rect 19300 11104 19809 11132
rect 19300 11092 19306 11104
rect 19797 11101 19809 11104
rect 19843 11101 19855 11135
rect 19797 11095 19855 11101
rect 20622 11092 20628 11144
rect 20680 11132 20686 11144
rect 20916 11132 20944 11163
rect 20680 11104 20944 11132
rect 20680 11092 20686 11104
rect 18782 10996 18788 11008
rect 17604 10968 18788 10996
rect 16540 10956 16546 10968
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 19242 10996 19248 11008
rect 19203 10968 19248 10996
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1820 10764 1961 10792
rect 1820 10752 1826 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 5537 10795 5595 10801
rect 4120 10764 5120 10792
rect 4120 10752 4126 10764
rect 5092 10724 5120 10764
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5626 10792 5632 10804
rect 5583 10764 5632 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6236 10764 6837 10792
rect 6236 10752 6242 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 9214 10792 9220 10804
rect 6825 10755 6883 10761
rect 6932 10764 9220 10792
rect 6932 10724 6960 10764
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9674 10792 9680 10804
rect 9635 10764 9680 10792
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 16482 10792 16488 10804
rect 11848 10764 16488 10792
rect 11848 10752 11854 10764
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 16761 10795 16819 10801
rect 16761 10761 16773 10795
rect 16807 10792 16819 10795
rect 16942 10792 16948 10804
rect 16807 10764 16948 10792
rect 16807 10761 16819 10764
rect 16761 10755 16819 10761
rect 16942 10752 16948 10764
rect 17000 10792 17006 10804
rect 17678 10792 17684 10804
rect 17000 10764 17684 10792
rect 17000 10752 17006 10764
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 21177 10795 21235 10801
rect 17972 10764 18184 10792
rect 11606 10724 11612 10736
rect 5092 10696 6960 10724
rect 9324 10696 11612 10724
rect 2222 10616 2228 10668
rect 2280 10656 2286 10668
rect 2501 10659 2559 10665
rect 2501 10656 2513 10659
rect 2280 10628 2513 10656
rect 2280 10616 2286 10628
rect 2501 10625 2513 10628
rect 2547 10625 2559 10659
rect 3602 10656 3608 10668
rect 3563 10628 3608 10656
rect 2501 10619 2559 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 7374 10656 7380 10668
rect 7335 10628 7380 10656
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 7466 10616 7472 10668
rect 7524 10656 7530 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 7524 10628 8217 10656
rect 7524 10616 7530 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 9324 10656 9352 10696
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 12158 10684 12164 10736
rect 12216 10724 12222 10736
rect 12216 10696 12848 10724
rect 12216 10684 12222 10696
rect 12820 10668 12848 10696
rect 9272 10628 9352 10656
rect 9272 10616 9278 10628
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10192 10628 10333 10656
rect 10192 10616 10198 10628
rect 10321 10625 10333 10628
rect 10367 10656 10379 10659
rect 11425 10659 11483 10665
rect 11425 10656 11437 10659
rect 10367 10628 11437 10656
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 11425 10625 11437 10628
rect 11471 10625 11483 10659
rect 11425 10619 11483 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 12618 10656 12624 10668
rect 11747 10628 12624 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14424 10628 15025 10656
rect 14424 10616 14430 10628
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15838 10656 15844 10668
rect 15436 10628 15844 10656
rect 15436 10616 15442 10628
rect 15838 10616 15844 10628
rect 15896 10656 15902 10668
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 15896 10628 16221 10656
rect 15896 10616 15902 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16500 10656 16528 10752
rect 17586 10684 17592 10736
rect 17644 10724 17650 10736
rect 17972 10724 18000 10764
rect 17644 10696 18000 10724
rect 18049 10727 18107 10733
rect 17644 10684 17650 10696
rect 18049 10693 18061 10727
rect 18095 10693 18107 10727
rect 18049 10687 18107 10693
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 16500 10628 17417 10656
rect 16209 10619 16267 10625
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 2958 10548 2964 10600
rect 3016 10588 3022 10600
rect 3329 10591 3387 10597
rect 3329 10588 3341 10591
rect 3016 10560 3341 10588
rect 3016 10548 3022 10560
rect 3329 10557 3341 10560
rect 3375 10557 3387 10591
rect 3329 10551 3387 10557
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10588 3479 10591
rect 3510 10588 3516 10600
rect 3467 10560 3516 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 4154 10588 4160 10600
rect 4115 10560 4160 10588
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 4948 10560 7420 10588
rect 4948 10548 4954 10560
rect 4424 10523 4482 10529
rect 4424 10489 4436 10523
rect 4470 10520 4482 10523
rect 4706 10520 4712 10532
rect 4470 10492 4712 10520
rect 4470 10489 4482 10492
rect 4424 10483 4482 10489
rect 4706 10480 4712 10492
rect 4764 10480 4770 10532
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 6730 10520 6736 10532
rect 5592 10492 6736 10520
rect 5592 10480 5598 10492
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 6972 10492 7297 10520
rect 6972 10480 6978 10492
rect 7285 10489 7297 10492
rect 7331 10489 7343 10523
rect 7392 10520 7420 10560
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7892 10560 8033 10588
rect 7892 10548 7898 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 8472 10591 8530 10597
rect 8472 10557 8484 10591
rect 8518 10588 8530 10591
rect 10152 10588 10180 10616
rect 8518 10560 10180 10588
rect 8518 10557 8530 10560
rect 8472 10551 8530 10557
rect 11238 10548 11244 10600
rect 11296 10548 11302 10600
rect 11330 10548 11336 10600
rect 11388 10588 11394 10600
rect 13072 10591 13130 10597
rect 11388 10560 11433 10588
rect 11388 10548 11394 10560
rect 13072 10557 13084 10591
rect 13118 10588 13130 10591
rect 14458 10588 14464 10600
rect 13118 10560 14464 10588
rect 13118 10557 13130 10560
rect 13072 10551 13130 10557
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10588 14979 10591
rect 15930 10588 15936 10600
rect 14967 10560 15936 10588
rect 14967 10557 14979 10560
rect 14921 10551 14979 10557
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10588 16083 10591
rect 17494 10588 17500 10600
rect 16071 10560 17500 10588
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 17494 10548 17500 10560
rect 17552 10548 17558 10600
rect 9122 10520 9128 10532
rect 7392 10492 9128 10520
rect 7285 10483 7343 10489
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 9214 10480 9220 10532
rect 9272 10520 9278 10532
rect 9398 10520 9404 10532
rect 9272 10492 9404 10520
rect 9272 10480 9278 10492
rect 9398 10480 9404 10492
rect 9456 10520 9462 10532
rect 10045 10523 10103 10529
rect 10045 10520 10057 10523
rect 9456 10492 10057 10520
rect 9456 10480 9462 10492
rect 10045 10489 10057 10492
rect 10091 10489 10103 10523
rect 10045 10483 10103 10489
rect 10137 10523 10195 10529
rect 10137 10489 10149 10523
rect 10183 10520 10195 10523
rect 11256 10520 11284 10548
rect 10183 10492 11284 10520
rect 10183 10489 10195 10492
rect 10137 10483 10195 10489
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 14829 10523 14887 10529
rect 13228 10492 14504 10520
rect 13228 10480 13234 10492
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 2317 10455 2375 10461
rect 2317 10452 2329 10455
rect 2280 10424 2329 10452
rect 2280 10412 2286 10424
rect 2317 10421 2329 10424
rect 2363 10421 2375 10455
rect 2317 10415 2375 10421
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2455 10424 2973 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 5350 10452 5356 10464
rect 3936 10424 5356 10452
rect 3936 10412 3942 10424
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 7006 10452 7012 10464
rect 6319 10424 7012 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7190 10452 7196 10464
rect 7151 10424 7196 10452
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7837 10455 7895 10461
rect 7837 10421 7849 10455
rect 7883 10452 7895 10455
rect 8386 10452 8392 10464
rect 7883 10424 8392 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 9582 10452 9588 10464
rect 9543 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 10284 10424 10885 10452
rect 10284 10412 10290 10424
rect 10873 10421 10885 10424
rect 10919 10421 10931 10455
rect 10873 10415 10931 10421
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11698 10452 11704 10464
rect 11287 10424 11704 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11698 10412 11704 10424
rect 11756 10452 11762 10464
rect 12710 10452 12716 10464
rect 11756 10424 12716 10452
rect 11756 10412 11762 10424
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14476 10461 14504 10492
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 17218 10520 17224 10532
rect 14875 10492 16896 10520
rect 17179 10492 17224 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 14185 10455 14243 10461
rect 14185 10452 14197 10455
rect 13872 10424 14197 10452
rect 13872 10412 13878 10424
rect 14185 10421 14197 10424
rect 14231 10421 14243 10455
rect 14185 10415 14243 10421
rect 14461 10455 14519 10461
rect 14461 10421 14473 10455
rect 14507 10421 14519 10455
rect 15654 10452 15660 10464
rect 15615 10424 15660 10452
rect 14461 10415 14519 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 15930 10412 15936 10464
rect 15988 10452 15994 10464
rect 16868 10461 16896 10492
rect 17218 10480 17224 10492
rect 17276 10520 17282 10532
rect 17862 10520 17868 10532
rect 17276 10492 17868 10520
rect 17276 10480 17282 10492
rect 17862 10480 17868 10492
rect 17920 10480 17926 10532
rect 18064 10520 18092 10687
rect 18156 10656 18184 10764
rect 21177 10761 21189 10795
rect 21223 10792 21235 10795
rect 21358 10792 21364 10804
rect 21223 10764 21364 10792
rect 21223 10761 21235 10764
rect 21177 10755 21235 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18156 10628 18613 10656
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18782 10616 18788 10668
rect 18840 10656 18846 10668
rect 19337 10659 19395 10665
rect 19337 10656 19349 10659
rect 18840 10628 19349 10656
rect 18840 10616 18846 10628
rect 19337 10625 19349 10628
rect 19383 10625 19395 10659
rect 19337 10619 19395 10625
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 19604 10591 19662 10597
rect 18555 10560 19564 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 19426 10520 19432 10532
rect 18064 10492 19432 10520
rect 19426 10480 19432 10492
rect 19484 10480 19490 10532
rect 19536 10520 19564 10560
rect 19604 10557 19616 10591
rect 19650 10588 19662 10591
rect 20070 10588 20076 10600
rect 19650 10560 20076 10588
rect 19650 10557 19662 10560
rect 19604 10551 19662 10557
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 20990 10588 20996 10600
rect 20951 10560 20996 10588
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 20806 10520 20812 10532
rect 19536 10492 20812 10520
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 16117 10455 16175 10461
rect 16117 10452 16129 10455
rect 15988 10424 16129 10452
rect 15988 10412 15994 10424
rect 16117 10421 16129 10424
rect 16163 10421 16175 10455
rect 16117 10415 16175 10421
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10421 16911 10455
rect 16853 10415 16911 10421
rect 17313 10455 17371 10461
rect 17313 10421 17325 10455
rect 17359 10452 17371 10455
rect 17678 10452 17684 10464
rect 17359 10424 17684 10452
rect 17359 10421 17371 10424
rect 17313 10415 17371 10421
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 17828 10424 20729 10452
rect 17828 10412 17834 10424
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 20717 10415 20775 10421
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 5534 10248 5540 10260
rect 3936 10220 5540 10248
rect 3936 10208 3942 10220
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6362 10248 6368 10260
rect 6319 10220 6368 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6362 10208 6368 10220
rect 6420 10248 6426 10260
rect 7098 10248 7104 10260
rect 6420 10220 7104 10248
rect 6420 10208 6426 10220
rect 7098 10208 7104 10220
rect 7156 10208 7162 10260
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10217 7987 10251
rect 8202 10248 8208 10260
rect 8163 10220 8208 10248
rect 7929 10211 7987 10217
rect 5160 10183 5218 10189
rect 5160 10149 5172 10183
rect 5206 10180 5218 10183
rect 7374 10180 7380 10192
rect 5206 10152 7380 10180
rect 5206 10149 5218 10152
rect 5160 10143 5218 10149
rect 7374 10140 7380 10152
rect 7432 10180 7438 10192
rect 7944 10180 7972 10211
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8570 10248 8576 10260
rect 8531 10220 8576 10248
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8665 10251 8723 10257
rect 8665 10217 8677 10251
rect 8711 10248 8723 10251
rect 9769 10251 9827 10257
rect 9769 10248 9781 10251
rect 8711 10220 9781 10248
rect 8711 10217 8723 10220
rect 8665 10211 8723 10217
rect 9769 10217 9781 10220
rect 9815 10217 9827 10251
rect 10226 10248 10232 10260
rect 10187 10220 10232 10248
rect 9769 10211 9827 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11204 10220 11989 10248
rect 11204 10208 11210 10220
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 7432 10152 7972 10180
rect 7432 10140 7438 10152
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10112 2651 10115
rect 3237 10115 3295 10121
rect 3237 10112 3249 10115
rect 2639 10084 3249 10112
rect 2639 10081 2651 10084
rect 2593 10075 2651 10081
rect 3237 10081 3249 10084
rect 3283 10081 3295 10115
rect 3237 10075 3295 10081
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4212 10084 4905 10112
rect 4212 10072 4218 10084
rect 4893 10081 4905 10084
rect 4939 10112 4951 10115
rect 4939 10084 5948 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10013 2743 10047
rect 2685 10007 2743 10013
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 3602 10044 3608 10056
rect 2915 10016 3608 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 2700 9976 2728 10007
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 5920 10044 5948 10084
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 6805 10115 6863 10121
rect 6805 10112 6817 10115
rect 6420 10084 6817 10112
rect 6420 10072 6426 10084
rect 6805 10081 6817 10084
rect 6851 10112 6863 10115
rect 6851 10084 7880 10112
rect 6851 10081 6863 10084
rect 6805 10075 6863 10081
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 5920 10016 6561 10044
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 2648 9948 2728 9976
rect 7852 9976 7880 10084
rect 7944 10044 7972 10152
rect 8938 10140 8944 10192
rect 8996 10180 9002 10192
rect 9122 10180 9128 10192
rect 8996 10152 9128 10180
rect 8996 10140 9002 10152
rect 9122 10140 9128 10152
rect 9180 10140 9186 10192
rect 10864 10183 10922 10189
rect 10864 10149 10876 10183
rect 10910 10180 10922 10183
rect 11238 10180 11244 10192
rect 10910 10152 11244 10180
rect 10910 10149 10922 10152
rect 10864 10143 10922 10149
rect 11238 10140 11244 10152
rect 11296 10180 11302 10192
rect 11790 10180 11796 10192
rect 11296 10152 11796 10180
rect 11296 10140 11302 10152
rect 11790 10140 11796 10152
rect 11848 10140 11854 10192
rect 11992 10180 12020 10211
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 13265 10251 13323 10257
rect 13265 10248 13277 10251
rect 12952 10220 13277 10248
rect 12952 10208 12958 10220
rect 13265 10217 13277 10220
rect 13311 10217 13323 10251
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13265 10211 13323 10217
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 17405 10251 17463 10257
rect 17405 10217 17417 10251
rect 17451 10248 17463 10251
rect 17451 10220 18368 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 12713 10183 12771 10189
rect 11992 10152 12572 10180
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 9824 10084 10149 10112
rect 9824 10072 9830 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10112 10655 10115
rect 12158 10112 12164 10124
rect 10643 10084 12164 10112
rect 10643 10081 10655 10084
rect 10597 10075 10655 10081
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 7944 10016 8769 10044
rect 8757 10013 8769 10016
rect 8803 10013 8815 10047
rect 8757 10007 8815 10013
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 12544 10044 12572 10152
rect 12713 10149 12725 10183
rect 12759 10180 12771 10183
rect 14182 10180 14188 10192
rect 12759 10152 14188 10180
rect 12759 10149 12771 10152
rect 12713 10143 12771 10149
rect 14182 10140 14188 10152
rect 14240 10140 14246 10192
rect 15746 10180 15752 10192
rect 15304 10152 15752 10180
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10112 12679 10115
rect 12667 10084 13032 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 13004 10056 13032 10084
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 15304 10121 15332 10152
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 15856 10152 17632 10180
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13596 10084 13737 10112
rect 13596 10072 13602 10084
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15556 10115 15614 10121
rect 15556 10112 15568 10115
rect 15436 10084 15568 10112
rect 15436 10072 15442 10084
rect 15556 10081 15568 10084
rect 15602 10112 15614 10115
rect 15856 10112 15884 10152
rect 15602 10084 15884 10112
rect 17313 10115 17371 10121
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 17313 10081 17325 10115
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12544 10016 12817 10044
rect 10321 10007 10379 10013
rect 12805 10013 12817 10016
rect 12851 10044 12863 10047
rect 12851 10016 12940 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 9582 9976 9588 9988
rect 7852 9948 9588 9976
rect 2648 9936 2654 9948
rect 9582 9936 9588 9948
rect 9640 9976 9646 9988
rect 10336 9976 10364 10007
rect 9640 9948 10364 9976
rect 9640 9936 9646 9948
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 12912 9976 12940 10016
rect 12986 10004 12992 10056
rect 13044 10004 13050 10056
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10044 13875 10047
rect 14366 10044 14372 10056
rect 13863 10016 14372 10044
rect 13863 10013 13875 10016
rect 13817 10007 13875 10013
rect 13832 9976 13860 10007
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 17126 10044 17132 10056
rect 17000 10016 17132 10044
rect 17000 10004 17006 10016
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 17218 10004 17224 10056
rect 17276 10044 17282 10056
rect 17328 10044 17356 10075
rect 17604 10053 17632 10152
rect 17276 10016 17356 10044
rect 17589 10047 17647 10053
rect 17276 10004 17282 10016
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 17954 9976 17960 9988
rect 11756 9948 12848 9976
rect 12912 9948 13860 9976
rect 16224 9948 17960 9976
rect 11756 9936 11762 9948
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6546 9908 6552 9920
rect 6052 9880 6552 9908
rect 6052 9868 6058 9880
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 11790 9908 11796 9920
rect 7800 9880 11796 9908
rect 7800 9868 7806 9880
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 12253 9911 12311 9917
rect 12253 9877 12265 9911
rect 12299 9908 12311 9911
rect 12618 9908 12624 9920
rect 12299 9880 12624 9908
rect 12299 9877 12311 9880
rect 12253 9871 12311 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12820 9908 12848 9948
rect 16224 9908 16252 9948
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 12820 9880 16252 9908
rect 16669 9911 16727 9917
rect 16669 9877 16681 9911
rect 16715 9908 16727 9911
rect 16758 9908 16764 9920
rect 16715 9880 16764 9908
rect 16715 9877 16727 9880
rect 16669 9871 16727 9877
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 16942 9908 16948 9920
rect 16903 9880 16948 9908
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 18340 9908 18368 10220
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 19242 10248 19248 10260
rect 18472 10220 19248 10248
rect 18472 10208 18478 10220
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 20128 10220 20269 10248
rect 20128 10208 20134 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 19144 10183 19202 10189
rect 19144 10149 19156 10183
rect 19190 10180 19202 10183
rect 19334 10180 19340 10192
rect 19190 10152 19340 10180
rect 19190 10149 19202 10152
rect 19144 10143 19202 10149
rect 19334 10140 19340 10152
rect 19392 10180 19398 10192
rect 21266 10180 21272 10192
rect 19392 10152 21272 10180
rect 19392 10140 19398 10152
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 18782 10072 18788 10124
rect 18840 10112 18846 10124
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 18840 10084 18889 10112
rect 18840 10072 18846 10084
rect 18877 10081 18889 10084
rect 18923 10081 18935 10115
rect 18877 10075 18935 10081
rect 20438 9908 20444 9920
rect 18340 9880 20444 9908
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2314 9704 2320 9716
rect 2087 9676 2320 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3016 9676 4200 9704
rect 3016 9664 3022 9676
rect 4172 9636 4200 9676
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 6730 9704 6736 9716
rect 5408 9676 6736 9704
rect 5408 9664 5414 9676
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7616 9676 7972 9704
rect 7616 9664 7622 9676
rect 5721 9639 5779 9645
rect 4172 9608 4476 9636
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 2608 9432 2636 9531
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 3108 9472 3249 9500
rect 3108 9460 3114 9472
rect 3237 9469 3249 9472
rect 3283 9500 3295 9503
rect 4062 9500 4068 9512
rect 3283 9472 4068 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 2608 9404 3280 9432
rect 3252 9376 3280 9404
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 3482 9435 3540 9441
rect 3482 9432 3494 9435
rect 3384 9404 3494 9432
rect 3384 9392 3390 9404
rect 3482 9401 3494 9404
rect 3528 9401 3540 9435
rect 4448 9432 4476 9608
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 6825 9639 6883 9645
rect 5767 9608 6500 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 6362 9568 6368 9580
rect 6275 9540 6368 9568
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6472 9568 6500 9608
rect 6825 9605 6837 9639
rect 6871 9636 6883 9639
rect 7190 9636 7196 9648
rect 6871 9608 7196 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7340 9608 7849 9636
rect 7340 9596 7346 9608
rect 7837 9605 7849 9608
rect 7883 9605 7895 9639
rect 7944 9636 7972 9676
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 9950 9704 9956 9716
rect 8168 9676 9956 9704
rect 8168 9664 8174 9676
rect 9950 9664 9956 9676
rect 10008 9704 10014 9716
rect 10008 9676 10640 9704
rect 10008 9664 10014 9676
rect 8938 9636 8944 9648
rect 7944 9608 8432 9636
rect 8899 9608 8944 9636
rect 7837 9599 7895 9605
rect 6914 9568 6920 9580
rect 6472 9540 6920 9568
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 8404 9577 8432 9608
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8496 9540 8708 9568
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5500 9472 6101 9500
rect 5500 9460 5506 9472
rect 6089 9469 6101 9472
rect 6135 9469 6147 9503
rect 6380 9500 6408 9528
rect 6380 9472 6500 9500
rect 6089 9463 6147 9469
rect 6472 9432 6500 9472
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 7064 9472 7205 9500
rect 7064 9460 7070 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7392 9432 7420 9531
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 8496 9500 8524 9540
rect 7616 9472 8524 9500
rect 7616 9460 7622 9472
rect 4448 9404 6316 9432
rect 6472 9404 7420 9432
rect 3482 9395 3540 9401
rect 2406 9364 2412 9376
rect 2367 9336 2412 9364
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 2556 9336 2601 9364
rect 2556 9324 2562 9336
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 4798 9364 4804 9376
rect 4663 9336 4804 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 4798 9324 4804 9336
rect 4856 9364 4862 9376
rect 5074 9364 5080 9376
rect 4856 9336 5080 9364
rect 4856 9324 4862 9336
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6288 9364 6316 9404
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 8386 9432 8392 9444
rect 7524 9404 8392 9432
rect 7524 9392 7530 9404
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8680 9432 8708 9540
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 9490 9568 9496 9580
rect 9451 9540 9496 9568
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 10505 9571 10563 9577
rect 10505 9537 10517 9571
rect 10551 9537 10563 9571
rect 10612 9568 10640 9676
rect 10686 9664 10692 9716
rect 10744 9664 10750 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 15746 9704 15752 9716
rect 12768 9676 13492 9704
rect 12768 9664 12774 9676
rect 10704 9636 10732 9664
rect 10962 9636 10968 9648
rect 10704 9608 10968 9636
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12492 9608 12537 9636
rect 12492 9596 12498 9608
rect 10686 9568 10692 9580
rect 10612 9540 10692 9568
rect 10505 9531 10563 9537
rect 9324 9500 9352 9528
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9324 9472 9413 9500
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9950 9460 9956 9512
rect 10008 9500 10014 9512
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 10008 9472 10333 9500
rect 10008 9460 10014 9472
rect 10321 9469 10333 9472
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 10520 9432 10548 9531
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 11514 9568 11520 9580
rect 11475 9540 11520 9568
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13464 9568 13492 9676
rect 14844 9676 15752 9704
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 14458 9636 14464 9648
rect 13872 9608 14464 9636
rect 13872 9596 13878 9608
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 14642 9596 14648 9648
rect 14700 9596 14706 9648
rect 13464 9540 13952 9568
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9500 11483 9503
rect 11882 9500 11888 9512
rect 11471 9472 11888 9500
rect 11471 9469 11483 9472
rect 11425 9463 11483 9469
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12676 9472 12817 9500
rect 12676 9460 12682 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13170 9500 13176 9512
rect 12943 9472 13176 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13814 9500 13820 9512
rect 13372 9472 13820 9500
rect 8680 9404 10548 9432
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 13372 9432 13400 9472
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 13924 9509 13952 9540
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 14056 9540 14105 9568
rect 14056 9528 14062 9540
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 14550 9500 14556 9512
rect 13955 9472 14556 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 14660 9509 14688 9596
rect 14844 9577 14872 9676
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 18782 9704 18788 9716
rect 18064 9676 18788 9704
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 16390 9568 16396 9580
rect 16264 9540 16396 9568
rect 16264 9528 16270 9540
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16816 9540 17049 9568
rect 16816 9528 16822 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17494 9568 17500 9580
rect 17455 9540 17500 9568
rect 17037 9531 17095 9537
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9469 14703 9503
rect 14645 9463 14703 9469
rect 15096 9503 15154 9509
rect 15096 9469 15108 9503
rect 15142 9500 15154 9503
rect 16776 9500 16804 9528
rect 15142 9472 16804 9500
rect 16853 9503 16911 9509
rect 15142 9469 15154 9472
rect 15096 9463 15154 9469
rect 16853 9469 16865 9503
rect 16899 9500 16911 9503
rect 16942 9500 16948 9512
rect 16899 9472 16948 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 18064 9509 18092 9676
rect 18782 9664 18788 9676
rect 18840 9704 18846 9716
rect 18840 9676 19288 9704
rect 18840 9664 18846 9676
rect 19260 9648 19288 9676
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 20622 9704 20628 9716
rect 20036 9676 20628 9704
rect 20036 9664 20042 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 19242 9596 19248 9648
rect 19300 9596 19306 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 19429 9639 19487 9645
rect 19429 9636 19441 9639
rect 19392 9608 19441 9636
rect 19392 9596 19398 9608
rect 19429 9605 19441 9608
rect 19475 9605 19487 9639
rect 19429 9599 19487 9605
rect 20990 9568 20996 9580
rect 20951 9540 20996 9568
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17460 9472 18061 9500
rect 17460 9460 17466 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 19150 9500 19156 9512
rect 18049 9463 18107 9469
rect 18248 9472 19156 9500
rect 18248 9432 18276 9472
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 19702 9460 19708 9512
rect 19760 9500 19766 9512
rect 20438 9500 20444 9512
rect 19760 9472 20444 9500
rect 19760 9460 19766 9472
rect 20438 9460 20444 9472
rect 20496 9500 20502 9512
rect 20809 9503 20867 9509
rect 20809 9500 20821 9503
rect 20496 9472 20821 9500
rect 20496 9460 20502 9472
rect 20809 9469 20821 9472
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 11379 9404 13400 9432
rect 13464 9404 18276 9432
rect 18316 9435 18374 9441
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6288 9336 7297 9364
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7432 9336 8217 9364
rect 7432 9324 7438 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8662 9364 8668 9376
rect 8343 9336 8668 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 9309 9367 9367 9373
rect 9309 9333 9321 9367
rect 9355 9364 9367 9367
rect 9766 9364 9772 9376
rect 9355 9336 9772 9364
rect 9355 9333 9367 9336
rect 9309 9327 9367 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10134 9364 10140 9376
rect 9999 9336 10140 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 13464 9373 13492 9404
rect 18316 9401 18328 9435
rect 18362 9432 18374 9435
rect 18782 9432 18788 9444
rect 18362 9404 18788 9432
rect 18362 9401 18374 9404
rect 18316 9395 18374 9401
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 18874 9392 18880 9444
rect 18932 9432 18938 9444
rect 21174 9432 21180 9444
rect 18932 9404 21180 9432
rect 18932 9392 18938 9404
rect 21174 9392 21180 9404
rect 21232 9392 21238 9444
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10459 9336 10977 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10965 9333 10977 9336
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 13449 9367 13507 9373
rect 13449 9333 13461 9367
rect 13495 9333 13507 9367
rect 13814 9364 13820 9376
rect 13775 9336 13820 9364
rect 13449 9327 13507 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 14461 9367 14519 9373
rect 14461 9333 14473 9367
rect 14507 9364 14519 9367
rect 14734 9364 14740 9376
rect 14507 9336 14740 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 16022 9364 16028 9376
rect 15252 9336 16028 9364
rect 15252 9324 15258 9336
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16206 9364 16212 9376
rect 16167 9336 16212 9364
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 16482 9364 16488 9376
rect 16443 9336 16488 9364
rect 16482 9324 16488 9336
rect 16540 9324 16546 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16724 9336 16957 9364
rect 16724 9324 16730 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 16945 9327 17003 9333
rect 18506 9324 18512 9376
rect 18564 9364 18570 9376
rect 19978 9364 19984 9376
rect 18564 9336 19984 9364
rect 18564 9324 18570 9336
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20441 9367 20499 9373
rect 20441 9333 20453 9367
rect 20487 9364 20499 9367
rect 20714 9364 20720 9376
rect 20487 9336 20720 9364
rect 20487 9333 20499 9336
rect 20441 9327 20499 9333
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 20901 9367 20959 9373
rect 20901 9333 20913 9367
rect 20947 9364 20959 9367
rect 21726 9364 21732 9376
rect 20947 9336 21732 9364
rect 20947 9333 20959 9336
rect 20901 9327 20959 9333
rect 21726 9324 21732 9336
rect 21784 9324 21790 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3326 9160 3332 9172
rect 3283 9132 3332 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 4028 9132 4077 9160
rect 4028 9120 4034 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 4571 9132 5089 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 5077 9129 5089 9132
rect 5123 9129 5135 9163
rect 5077 9123 5135 9129
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 5491 9132 6101 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 6089 9129 6101 9132
rect 6135 9129 6147 9163
rect 6089 9123 6147 9129
rect 6457 9163 6515 9169
rect 6457 9129 6469 9163
rect 6503 9160 6515 9163
rect 6638 9160 6644 9172
rect 6503 9132 6644 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 6638 9120 6644 9132
rect 6696 9160 6702 9172
rect 8938 9160 8944 9172
rect 6696 9132 8147 9160
rect 8899 9132 8944 9160
rect 6696 9120 6702 9132
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5040 9064 5396 9092
rect 5040 9052 5046 9064
rect 5368 9036 5396 9064
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 7006 9092 7012 9104
rect 6880 9064 7012 9092
rect 6880 9052 6886 9064
rect 7006 9052 7012 9064
rect 7064 9052 7070 9104
rect 7561 9095 7619 9101
rect 7561 9061 7573 9095
rect 7607 9092 7619 9095
rect 8018 9092 8024 9104
rect 7607 9064 8024 9092
rect 7607 9061 7619 9064
rect 7561 9055 7619 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 1946 9024 1952 9036
rect 1903 8996 1952 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 2124 9027 2182 9033
rect 2124 8993 2136 9027
rect 2170 9024 2182 9027
rect 4433 9027 4491 9033
rect 2170 8996 2912 9024
rect 2170 8993 2182 8996
rect 2124 8987 2182 8993
rect 2884 8956 2912 8996
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 5258 9024 5264 9036
rect 4479 8996 5264 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5350 8984 5356 9036
rect 5408 9024 5414 9036
rect 7374 9024 7380 9036
rect 5408 8996 7380 9024
rect 5408 8984 5414 8996
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 8119 9024 8147 9132
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9033 9163 9091 9169
rect 9033 9129 9045 9163
rect 9079 9160 9091 9163
rect 9677 9163 9735 9169
rect 9079 9132 9536 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 9401 9095 9459 9101
rect 9401 9092 9413 9095
rect 8864 9064 9413 9092
rect 8864 9024 8892 9064
rect 9401 9061 9413 9064
rect 9447 9061 9459 9095
rect 9401 9055 9459 9061
rect 7515 8996 8064 9024
rect 8119 8996 8892 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 3234 8956 3240 8968
rect 2884 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8956 3298 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 3292 8928 4629 8956
rect 3292 8916 3298 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5552 8888 5580 8919
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 6546 8956 6552 8968
rect 5684 8928 5729 8956
rect 6507 8928 6552 8956
rect 5684 8916 5690 8928
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 6822 8956 6828 8968
rect 6779 8928 6828 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 6822 8916 6828 8928
rect 6880 8956 6886 8968
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 6880 8928 7665 8956
rect 6880 8916 6886 8928
rect 7653 8925 7665 8928
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7101 8891 7159 8897
rect 7101 8888 7113 8891
rect 5552 8860 7113 8888
rect 7101 8857 7113 8860
rect 7147 8857 7159 8891
rect 8036 8888 8064 8996
rect 8938 8984 8944 9036
rect 8996 9024 9002 9036
rect 9508 9024 9536 9132
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9723 9132 10160 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 10132 9092 10160 9132
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 11882 9160 11888 9172
rect 10284 9132 11888 9160
rect 10284 9120 10290 9132
rect 11882 9120 11888 9132
rect 11940 9160 11946 9172
rect 12894 9160 12900 9172
rect 11940 9132 12900 9160
rect 11940 9120 11946 9132
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 13136 9132 14657 9160
rect 13136 9120 13142 9132
rect 14645 9129 14657 9132
rect 14691 9160 14703 9163
rect 15194 9160 15200 9172
rect 14691 9132 15200 9160
rect 14691 9129 14703 9132
rect 14645 9123 14703 9129
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15749 9163 15807 9169
rect 15749 9129 15761 9163
rect 15795 9160 15807 9163
rect 16482 9160 16488 9172
rect 15795 9132 16488 9160
rect 15795 9129 15807 9132
rect 15749 9123 15807 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 19242 9160 19248 9172
rect 18196 9132 19248 9160
rect 18196 9120 18202 9132
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 19521 9163 19579 9169
rect 19521 9160 19533 9163
rect 19484 9132 19533 9160
rect 19484 9120 19490 9132
rect 19521 9129 19533 9132
rect 19567 9129 19579 9163
rect 19521 9123 19579 9129
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 21634 9160 21640 9172
rect 20947 9132 21640 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 9640 9064 10088 9092
rect 10132 9064 10916 9092
rect 9640 9052 9646 9064
rect 9674 9024 9680 9036
rect 8996 8996 9168 9024
rect 9508 8996 9680 9024
rect 8996 8984 9002 8996
rect 9140 8965 9168 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10060 9024 10088 9064
rect 10117 9027 10175 9033
rect 10117 9024 10129 9027
rect 10060 8996 10129 9024
rect 10117 8993 10129 8996
rect 10163 8993 10175 9027
rect 10117 8987 10175 8993
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8956 8171 8959
rect 9125 8959 9183 8965
rect 8159 8928 8800 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8573 8891 8631 8897
rect 8036 8860 8524 8888
rect 7101 8851 7159 8857
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 8294 8820 8300 8832
rect 4304 8792 8300 8820
rect 4304 8780 4310 8792
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8496 8820 8524 8860
rect 8573 8857 8585 8891
rect 8619 8888 8631 8891
rect 8662 8888 8668 8900
rect 8619 8860 8668 8888
rect 8619 8857 8631 8860
rect 8573 8851 8631 8857
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 8772 8888 8800 8928
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9456 8928 9873 8956
rect 9456 8916 9462 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 9766 8888 9772 8900
rect 8772 8860 9772 8888
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 10502 8820 10508 8832
rect 8496 8792 10508 8820
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10888 8820 10916 9064
rect 11054 9052 11060 9104
rect 11112 9092 11118 9104
rect 11514 9092 11520 9104
rect 11112 9064 11520 9092
rect 11112 9052 11118 9064
rect 11514 9052 11520 9064
rect 11572 9092 11578 9104
rect 12434 9092 12440 9104
rect 11572 9064 12440 9092
rect 11572 9052 11578 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 12612 9095 12670 9101
rect 12612 9061 12624 9095
rect 12658 9092 12670 9095
rect 13630 9092 13636 9104
rect 12658 9064 13636 9092
rect 12658 9061 12670 9064
rect 12612 9055 12670 9061
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 15212 9064 18460 9092
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 13078 9024 13084 9036
rect 11020 8996 13084 9024
rect 11020 8984 11026 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 13372 8996 14565 9024
rect 13372 8968 13400 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 15212 9024 15240 9064
rect 14553 8987 14611 8993
rect 14752 8996 15240 9024
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 12216 8928 12357 8956
rect 12216 8916 12222 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 13354 8916 13360 8968
rect 13412 8916 13418 8968
rect 11238 8888 11244 8900
rect 11199 8860 11244 8888
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 13722 8888 13728 8900
rect 13635 8860 13728 8888
rect 13722 8848 13728 8860
rect 13780 8888 13786 8900
rect 14752 8888 14780 8996
rect 15286 8984 15292 9036
rect 15344 9024 15350 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15344 8996 15669 9024
rect 15344 8984 15350 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 16666 9024 16672 9036
rect 16627 8996 16672 9024
rect 15657 8987 15715 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 17494 9024 17500 9036
rect 16868 8996 17500 9024
rect 16868 8968 16896 8996
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 17672 9027 17730 9033
rect 17672 8993 17684 9027
rect 17718 9024 17730 9027
rect 18138 9024 18144 9036
rect 17718 8996 18144 9024
rect 17718 8993 17730 8996
rect 17672 8987 17730 8993
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 14829 8959 14887 8965
rect 14829 8925 14841 8959
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 13780 8860 14780 8888
rect 14844 8888 14872 8919
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15252 8928 15853 8956
rect 15252 8916 15258 8928
rect 15841 8925 15853 8928
rect 15887 8956 15899 8959
rect 16206 8956 16212 8968
rect 15887 8928 16212 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 16761 8959 16819 8965
rect 16761 8956 16773 8959
rect 16632 8928 16773 8956
rect 16632 8916 16638 8928
rect 16761 8925 16773 8928
rect 16807 8925 16819 8959
rect 16761 8919 16819 8925
rect 15289 8891 15347 8897
rect 14844 8860 15240 8888
rect 13780 8848 13786 8860
rect 13814 8820 13820 8832
rect 10888 8792 13820 8820
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14185 8823 14243 8829
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 15102 8820 15108 8832
rect 14231 8792 15108 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15212 8820 15240 8860
rect 15289 8857 15301 8891
rect 15335 8888 15347 8891
rect 16114 8888 16120 8900
rect 15335 8860 16120 8888
rect 15335 8857 15347 8860
rect 15289 8851 15347 8857
rect 16114 8848 16120 8860
rect 16172 8848 16178 8900
rect 16390 8888 16396 8900
rect 16224 8860 16396 8888
rect 16224 8832 16252 8860
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 16776 8888 16804 8919
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 17402 8956 17408 8968
rect 16908 8928 16953 8956
rect 17363 8928 17408 8956
rect 16908 8916 16914 8928
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 18432 8956 18460 9064
rect 18506 9052 18512 9104
rect 18564 9092 18570 9104
rect 21266 9092 21272 9104
rect 18564 9064 21272 9092
rect 18564 9052 18570 9064
rect 21266 9052 21272 9064
rect 21324 9052 21330 9104
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 9024 18935 9027
rect 19334 9024 19340 9036
rect 18923 8996 19340 9024
rect 18923 8993 18935 8996
rect 18877 8987 18935 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 9024 19487 9027
rect 19794 9024 19800 9036
rect 19475 8996 19800 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 19613 8959 19671 8965
rect 19613 8956 19625 8959
rect 18432 8928 19625 8956
rect 19613 8925 19625 8928
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 16942 8888 16948 8900
rect 16776 8860 16948 8888
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 18782 8888 18788 8900
rect 18743 8860 18788 8888
rect 18782 8848 18788 8860
rect 18840 8888 18846 8900
rect 19794 8888 19800 8900
rect 18840 8860 19800 8888
rect 18840 8848 18846 8860
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 15378 8820 15384 8832
rect 15212 8792 15384 8820
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 16206 8780 16212 8832
rect 16264 8780 16270 8832
rect 16301 8823 16359 8829
rect 16301 8789 16313 8823
rect 16347 8820 16359 8823
rect 17310 8820 17316 8832
rect 16347 8792 17316 8820
rect 16347 8789 16359 8792
rect 16301 8783 16359 8789
rect 17310 8780 17316 8792
rect 17368 8780 17374 8832
rect 18138 8780 18144 8832
rect 18196 8820 18202 8832
rect 18877 8823 18935 8829
rect 18877 8820 18889 8823
rect 18196 8792 18889 8820
rect 18196 8780 18202 8792
rect 18877 8789 18889 8792
rect 18923 8789 18935 8823
rect 18877 8783 18935 8789
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19061 8823 19119 8829
rect 19061 8820 19073 8823
rect 19024 8792 19073 8820
rect 19024 8780 19030 8792
rect 19061 8789 19073 8792
rect 19107 8789 19119 8823
rect 19061 8783 19119 8789
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 20070 8820 20076 8832
rect 19576 8792 20076 8820
rect 19576 8780 19582 8792
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 3234 8616 3240 8628
rect 3195 8588 3240 8616
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5258 8616 5264 8628
rect 4856 8588 5120 8616
rect 5219 8588 5264 8616
rect 4856 8576 4862 8588
rect 4985 8551 5043 8557
rect 4985 8517 4997 8551
rect 5031 8517 5043 8551
rect 5092 8548 5120 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 7190 8616 7196 8628
rect 6840 8588 7196 8616
rect 6273 8551 6331 8557
rect 6273 8548 6285 8551
rect 5092 8520 6285 8548
rect 4985 8511 5043 8517
rect 6273 8517 6285 8520
rect 6319 8517 6331 8551
rect 6273 8511 6331 8517
rect 5000 8480 5028 8511
rect 5626 8480 5632 8492
rect 5000 8452 5632 8480
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 1946 8412 1952 8424
rect 1903 8384 1952 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 1946 8372 1952 8384
rect 2004 8412 2010 8424
rect 3050 8412 3056 8424
rect 2004 8384 3056 8412
rect 2004 8372 2010 8384
rect 3050 8372 3056 8384
rect 3108 8412 3114 8424
rect 3326 8412 3332 8424
rect 3108 8384 3332 8412
rect 3108 8372 3114 8384
rect 3326 8372 3332 8384
rect 3384 8412 3390 8424
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3384 8384 3617 8412
rect 3384 8372 3390 8384
rect 3605 8381 3617 8384
rect 3651 8381 3663 8415
rect 5000 8412 5028 8452
rect 5626 8440 5632 8452
rect 5684 8480 5690 8492
rect 6840 8489 6868 8588
rect 7190 8576 7196 8588
rect 7248 8616 7254 8628
rect 8294 8616 8300 8628
rect 7248 8588 8300 8616
rect 7248 8576 7254 8588
rect 8294 8576 8300 8588
rect 8352 8616 8358 8628
rect 9398 8616 9404 8628
rect 8352 8588 9404 8616
rect 8352 8576 8358 8588
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 7852 8520 8217 8548
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5684 8452 5825 8480
rect 5684 8440 5690 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 7098 8421 7104 8424
rect 6457 8415 6515 8421
rect 3605 8375 3663 8381
rect 3712 8384 5028 8412
rect 5460 8384 5856 8412
rect 2124 8347 2182 8353
rect 2124 8313 2136 8347
rect 2170 8344 2182 8347
rect 2682 8344 2688 8356
rect 2170 8316 2688 8344
rect 2170 8313 2182 8316
rect 2124 8307 2182 8313
rect 2682 8304 2688 8316
rect 2740 8344 2746 8356
rect 3712 8344 3740 8384
rect 3878 8353 3884 8356
rect 3872 8344 3884 8353
rect 2740 8316 3740 8344
rect 3839 8316 3884 8344
rect 2740 8304 2746 8316
rect 3872 8307 3884 8316
rect 3878 8304 3884 8307
rect 3936 8304 3942 8356
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 5460 8276 5488 8384
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 5592 8316 5733 8344
rect 5592 8304 5598 8316
rect 5721 8313 5733 8316
rect 5767 8313 5779 8347
rect 5721 8307 5779 8313
rect 5626 8276 5632 8288
rect 4120 8248 5488 8276
rect 5587 8248 5632 8276
rect 4120 8236 4126 8248
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 5828 8276 5856 8384
rect 6457 8381 6469 8415
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 7092 8375 7104 8421
rect 7156 8412 7162 8424
rect 7156 8384 7192 8412
rect 6472 8344 6500 8375
rect 7098 8372 7104 8375
rect 7156 8372 7162 8384
rect 7466 8372 7472 8424
rect 7524 8412 7530 8424
rect 7852 8412 7880 8520
rect 8205 8517 8217 8520
rect 8251 8517 8263 8551
rect 8205 8511 8263 8517
rect 8496 8489 8524 8588
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 9640 8588 11529 8616
rect 9640 8576 9646 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12437 8619 12495 8625
rect 12437 8616 12449 8619
rect 12308 8588 12449 8616
rect 12308 8576 12314 8588
rect 12437 8585 12449 8588
rect 12483 8585 12495 8619
rect 12437 8579 12495 8585
rect 14090 8576 14096 8628
rect 14148 8616 14154 8628
rect 16666 8616 16672 8628
rect 14148 8588 16672 8616
rect 14148 8576 14154 8588
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 20622 8616 20628 8628
rect 16776 8588 20628 8616
rect 9416 8548 9444 8576
rect 9861 8551 9919 8557
rect 9416 8520 9536 8548
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 9508 8480 9536 8520
rect 9861 8517 9873 8551
rect 9907 8548 9919 8551
rect 9953 8551 10011 8557
rect 9953 8548 9965 8551
rect 9907 8520 9965 8548
rect 9907 8517 9919 8520
rect 9861 8511 9919 8517
rect 9953 8517 9965 8520
rect 9999 8517 10011 8551
rect 9953 8511 10011 8517
rect 13633 8551 13691 8557
rect 13633 8517 13645 8551
rect 13679 8548 13691 8551
rect 16776 8548 16804 8588
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 13679 8520 16804 8548
rect 13679 8517 13691 8520
rect 13633 8511 13691 8517
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 18196 8520 18245 8548
rect 18196 8508 18202 8520
rect 18233 8517 18245 8520
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 18877 8551 18935 8557
rect 18877 8517 18889 8551
rect 18923 8548 18935 8551
rect 19426 8548 19432 8560
rect 18923 8520 19432 8548
rect 18923 8517 18935 8520
rect 18877 8511 18935 8517
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 20990 8548 20996 8560
rect 19904 8520 20996 8548
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9508 8452 10149 8480
rect 8481 8443 8539 8449
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 11330 8440 11336 8492
rect 11388 8480 11394 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 11388 8452 13001 8480
rect 11388 8440 11394 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 14056 8452 14197 8480
rect 14056 8440 14062 8452
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 15010 8440 15016 8492
rect 15068 8440 15074 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15160 8452 15761 8480
rect 15160 8440 15166 8452
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 16758 8480 16764 8492
rect 15979 8452 16764 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 16908 8452 16953 8480
rect 16908 8440 16914 8452
rect 17034 8440 17040 8492
rect 17092 8480 17098 8492
rect 17092 8452 19012 8480
rect 17092 8440 17098 8452
rect 7524 8384 7880 8412
rect 8748 8415 8806 8421
rect 7524 8372 7530 8384
rect 8748 8381 8760 8415
rect 8794 8412 8806 8415
rect 9490 8412 9496 8424
rect 8794 8384 9496 8412
rect 8794 8381 8806 8384
rect 8748 8375 8806 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 14090 8412 14096 8424
rect 10284 8384 14096 8412
rect 10284 8372 10290 8384
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 8478 8344 8484 8356
rect 6472 8316 8484 8344
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 9953 8347 10011 8353
rect 9953 8344 9965 8347
rect 8996 8316 9965 8344
rect 8996 8304 9002 8316
rect 9953 8313 9965 8316
rect 9999 8344 10011 8347
rect 10382 8347 10440 8353
rect 10382 8344 10394 8347
rect 9999 8316 10394 8344
rect 9999 8313 10011 8316
rect 9953 8307 10011 8313
rect 10382 8313 10394 8316
rect 10428 8313 10440 8347
rect 10382 8307 10440 8313
rect 10594 8304 10600 8356
rect 10652 8344 10658 8356
rect 11698 8344 11704 8356
rect 10652 8316 11704 8344
rect 10652 8304 10658 8316
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 12802 8344 12808 8356
rect 12763 8316 12808 8344
rect 12802 8304 12808 8316
rect 12860 8344 12866 8356
rect 13265 8347 13323 8353
rect 13265 8344 13277 8347
rect 12860 8316 13277 8344
rect 12860 8304 12866 8316
rect 13265 8313 13277 8316
rect 13311 8313 13323 8347
rect 13265 8307 13323 8313
rect 14001 8347 14059 8353
rect 14001 8313 14013 8347
rect 14047 8344 14059 8347
rect 14366 8344 14372 8356
rect 14047 8316 14372 8344
rect 14047 8313 14059 8316
rect 14001 8307 14059 8313
rect 14366 8304 14372 8316
rect 14424 8344 14430 8356
rect 14642 8344 14648 8356
rect 14424 8316 14648 8344
rect 14424 8304 14430 8316
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 11146 8276 11152 8288
rect 5828 8248 11152 8276
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 12897 8279 12955 8285
rect 12897 8276 12909 8279
rect 11296 8248 12909 8276
rect 11296 8236 11302 8248
rect 12897 8245 12909 8248
rect 12943 8276 12955 8279
rect 13906 8276 13912 8288
rect 12943 8248 13912 8276
rect 12943 8245 12955 8248
rect 12897 8239 12955 8245
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 14090 8276 14096 8288
rect 14051 8248 14096 8276
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 15028 8285 15056 8440
rect 15197 8415 15255 8421
rect 15197 8412 15209 8415
rect 15120 8384 15209 8412
rect 15120 8356 15148 8384
rect 15197 8381 15209 8384
rect 15243 8381 15255 8415
rect 15197 8375 15255 8381
rect 15286 8372 15292 8424
rect 15344 8372 15350 8424
rect 15654 8412 15660 8424
rect 15615 8384 15660 8412
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18984 8412 19012 8452
rect 19058 8440 19064 8492
rect 19116 8480 19122 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19116 8452 19349 8480
rect 19116 8440 19122 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 19904 8480 19932 8520
rect 20640 8492 20668 8520
rect 20990 8508 20996 8520
rect 21048 8508 21054 8560
rect 20622 8480 20628 8492
rect 19567 8452 19932 8480
rect 20583 8452 20628 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 18984 8384 20300 8412
rect 15102 8304 15108 8356
rect 15160 8304 15166 8356
rect 15304 8285 15332 8372
rect 16758 8344 16764 8356
rect 16719 8316 16764 8344
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17678 8304 17684 8356
rect 17736 8344 17742 8356
rect 18782 8344 18788 8356
rect 17736 8316 18788 8344
rect 17736 8304 17742 8316
rect 18782 8304 18788 8316
rect 18840 8344 18846 8356
rect 19245 8347 19303 8353
rect 19245 8344 19257 8347
rect 18840 8316 19257 8344
rect 18840 8304 18846 8316
rect 19245 8313 19257 8316
rect 19291 8313 19303 8347
rect 20272 8344 20300 8384
rect 20272 8316 20576 8344
rect 19245 8307 19303 8313
rect 15013 8279 15071 8285
rect 15013 8245 15025 8279
rect 15059 8245 15071 8279
rect 15013 8239 15071 8245
rect 15289 8279 15347 8285
rect 15289 8245 15301 8279
rect 15335 8245 15347 8279
rect 16298 8276 16304 8288
rect 16259 8248 16304 8276
rect 15289 8239 15347 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 16666 8276 16672 8288
rect 16627 8248 16672 8276
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 17586 8236 17592 8288
rect 17644 8276 17650 8288
rect 17770 8276 17776 8288
rect 17644 8248 17776 8276
rect 17644 8236 17650 8248
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 18322 8236 18328 8288
rect 18380 8276 18386 8288
rect 19334 8276 19340 8288
rect 18380 8248 19340 8276
rect 18380 8236 18386 8248
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 20070 8276 20076 8288
rect 20031 8248 20076 8276
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 20346 8236 20352 8288
rect 20404 8276 20410 8288
rect 20548 8285 20576 8316
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 20404 8248 20453 8276
rect 20404 8236 20410 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 20441 8239 20499 8245
rect 20533 8279 20591 8285
rect 20533 8245 20545 8279
rect 20579 8276 20591 8279
rect 21450 8276 21456 8288
rect 20579 8248 21456 8276
rect 20579 8245 20591 8248
rect 20533 8239 20591 8245
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2406 8072 2412 8084
rect 2179 8044 2412 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 4985 8075 5043 8081
rect 4985 8041 4997 8075
rect 5031 8072 5043 8075
rect 5534 8072 5540 8084
rect 5031 8044 5540 8072
rect 5031 8041 5043 8044
rect 4985 8035 5043 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 5684 8044 6285 8072
rect 5684 8032 5690 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 7791 8044 8248 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 1670 7964 1676 8016
rect 1728 8004 1734 8016
rect 2590 8004 2596 8016
rect 1728 7976 2596 8004
rect 1728 7964 1734 7976
rect 2590 7964 2596 7976
rect 2648 8004 2654 8016
rect 5994 8004 6000 8016
rect 2648 7976 6000 8004
rect 2648 7964 2654 7976
rect 5994 7964 6000 7976
rect 6052 7964 6058 8016
rect 6362 7964 6368 8016
rect 6420 8004 6426 8016
rect 6641 8007 6699 8013
rect 6641 8004 6653 8007
rect 6420 7976 6653 8004
rect 6420 7964 6426 7976
rect 6641 7973 6653 7976
rect 6687 8004 6699 8007
rect 7374 8004 7380 8016
rect 6687 7976 7380 8004
rect 6687 7973 6699 7976
rect 6641 7967 6699 7973
rect 7374 7964 7380 7976
rect 7432 7964 7438 8016
rect 8220 8004 8248 8044
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8352 8044 8397 8072
rect 8352 8032 8358 8044
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8720 8044 8953 8072
rect 8720 8032 8726 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 9953 8075 10011 8081
rect 9953 8041 9965 8075
rect 9999 8072 10011 8075
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 9999 8044 11345 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 11333 8041 11345 8044
rect 11379 8041 11391 8075
rect 11333 8035 11391 8041
rect 11425 8075 11483 8081
rect 11425 8041 11437 8075
rect 11471 8072 11483 8075
rect 13170 8072 13176 8084
rect 11471 8044 13176 8072
rect 11471 8041 11483 8044
rect 11425 8035 11483 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 15654 8072 15660 8084
rect 14148 8044 15660 8072
rect 14148 8032 14154 8044
rect 15654 8032 15660 8044
rect 15712 8072 15718 8084
rect 16206 8072 16212 8084
rect 15712 8044 16212 8072
rect 15712 8032 15718 8044
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16724 8044 16957 8072
rect 16724 8032 16730 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 16945 8035 17003 8041
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17092 8044 17325 8072
rect 17092 8032 17098 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 17460 8044 17505 8072
rect 17460 8032 17466 8044
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18417 8075 18475 8081
rect 18417 8072 18429 8075
rect 18380 8044 18429 8072
rect 18380 8032 18386 8044
rect 18417 8041 18429 8044
rect 18463 8041 18475 8075
rect 18417 8035 18475 8041
rect 8220 7976 9720 8004
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 2547 7908 3157 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 3145 7905 3157 7908
rect 3191 7905 3203 7939
rect 5350 7936 5356 7948
rect 5311 7908 5356 7936
rect 3145 7899 3203 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7936 5503 7939
rect 5810 7936 5816 7948
rect 5491 7908 5816 7936
rect 5491 7905 5503 7908
rect 5445 7899 5503 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 6914 7936 6920 7948
rect 6779 7908 6920 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 8202 7936 8208 7948
rect 7699 7908 8208 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 3936 7840 5549 7868
rect 3936 7828 3942 7840
rect 5537 7837 5549 7840
rect 5583 7868 5595 7871
rect 6822 7868 6828 7880
rect 5583 7840 6828 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 7892 7840 7937 7868
rect 7892 7828 7898 7840
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8076 7840 9045 7868
rect 8076 7828 8082 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9582 7868 9588 7880
rect 9263 7840 9588 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9692 7868 9720 7976
rect 9766 7964 9772 8016
rect 9824 8004 9830 8016
rect 10413 8007 10471 8013
rect 10413 8004 10425 8007
rect 9824 7976 10425 8004
rect 9824 7964 9830 7976
rect 10413 7973 10425 7976
rect 10459 7973 10471 8007
rect 14734 8004 14740 8016
rect 10413 7967 10471 7973
rect 12636 7976 14740 8004
rect 12636 7945 12664 7976
rect 14734 7964 14740 7976
rect 14792 7964 14798 8016
rect 15746 8004 15752 8016
rect 14844 7976 15752 8004
rect 10321 7939 10379 7945
rect 10321 7905 10333 7939
rect 10367 7936 10379 7939
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 10367 7908 11989 7936
rect 10367 7905 10379 7908
rect 10321 7899 10379 7905
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 11977 7899 12035 7905
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 12980 7939 13038 7945
rect 12980 7905 12992 7939
rect 13026 7936 13038 7939
rect 13722 7936 13728 7948
rect 13026 7908 13728 7936
rect 13026 7905 13038 7908
rect 12980 7899 13038 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 14366 7936 14372 7948
rect 14327 7908 14372 7936
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 14844 7936 14872 7976
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 19306 8007 19364 8013
rect 19306 8004 19318 8007
rect 18932 7976 19318 8004
rect 18932 7964 18938 7976
rect 19306 7973 19318 7976
rect 19352 7973 19364 8007
rect 19306 7967 19364 7973
rect 19978 7964 19984 8016
rect 20036 7964 20042 8016
rect 15286 7936 15292 7948
rect 14700 7908 14872 7936
rect 15247 7908 15292 7936
rect 14700 7896 14706 7908
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15378 7896 15384 7948
rect 15436 7936 15442 7948
rect 15556 7939 15614 7945
rect 15556 7936 15568 7939
rect 15436 7908 15568 7936
rect 15436 7896 15442 7908
rect 15556 7905 15568 7908
rect 15602 7936 15614 7939
rect 18325 7939 18383 7945
rect 15602 7908 17540 7936
rect 15602 7905 15614 7908
rect 15556 7899 15614 7905
rect 17512 7880 17540 7908
rect 18325 7905 18337 7939
rect 18371 7936 18383 7939
rect 19150 7936 19156 7948
rect 18371 7908 19156 7936
rect 18371 7905 18383 7908
rect 18325 7899 18383 7905
rect 19150 7896 19156 7908
rect 19208 7936 19214 7948
rect 19996 7936 20024 7964
rect 19208 7908 20024 7936
rect 19208 7896 19214 7908
rect 9766 7868 9772 7880
rect 9692 7840 9772 7868
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 10594 7868 10600 7880
rect 10555 7840 10600 7868
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10870 7828 10876 7880
rect 10928 7828 10934 7880
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 11790 7868 11796 7880
rect 11655 7840 11796 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 7190 7800 7196 7812
rect 4028 7772 7196 7800
rect 4028 7760 4034 7772
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 7285 7803 7343 7809
rect 7285 7769 7297 7803
rect 7331 7800 7343 7803
rect 10888 7800 10916 7828
rect 7331 7772 7788 7800
rect 7331 7769 7343 7772
rect 7285 7763 7343 7769
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 7558 7732 7564 7744
rect 6236 7704 7564 7732
rect 6236 7692 6242 7704
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7760 7732 7788 7772
rect 8496 7772 10916 7800
rect 8496 7732 8524 7772
rect 12728 7744 12756 7831
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 17678 7868 17684 7880
rect 17552 7840 17684 7868
rect 17552 7828 17558 7840
rect 17678 7828 17684 7840
rect 17736 7868 17742 7880
rect 18509 7871 18567 7877
rect 17736 7840 18368 7868
rect 17736 7828 17742 7840
rect 18340 7800 18368 7840
rect 18509 7837 18521 7871
rect 18555 7837 18567 7871
rect 19058 7868 19064 7880
rect 19019 7840 19064 7868
rect 18509 7831 18567 7837
rect 18524 7800 18552 7831
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 18340 7772 18552 7800
rect 7760 7704 8524 7732
rect 8573 7735 8631 7741
rect 8573 7701 8585 7735
rect 8619 7732 8631 7735
rect 10870 7732 10876 7744
rect 8619 7704 10876 7732
rect 8619 7701 8631 7704
rect 8573 7695 8631 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 10965 7735 11023 7741
rect 10965 7701 10977 7735
rect 11011 7732 11023 7735
rect 11238 7732 11244 7744
rect 11011 7704 11244 7732
rect 11011 7701 11023 7704
rect 10965 7695 11023 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 12158 7692 12164 7744
rect 12216 7732 12222 7744
rect 12437 7735 12495 7741
rect 12437 7732 12449 7735
rect 12216 7704 12449 7732
rect 12216 7692 12222 7704
rect 12437 7701 12449 7704
rect 12483 7732 12495 7735
rect 12710 7732 12716 7744
rect 12483 7704 12716 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14550 7732 14556 7744
rect 14148 7704 14193 7732
rect 14511 7704 14556 7732
rect 14148 7692 14154 7704
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 16850 7732 16856 7744
rect 16715 7704 16856 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 16850 7692 16856 7704
rect 16908 7732 16914 7744
rect 17586 7732 17592 7744
rect 16908 7704 17592 7732
rect 16908 7692 16914 7704
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 17954 7732 17960 7744
rect 17915 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 20441 7735 20499 7741
rect 20441 7701 20453 7735
rect 20487 7732 20499 7735
rect 20622 7732 20628 7744
rect 20487 7704 20628 7732
rect 20487 7701 20499 7704
rect 20441 7695 20499 7701
rect 20622 7692 20628 7704
rect 20680 7732 20686 7744
rect 21542 7732 21548 7744
rect 20680 7704 21548 7732
rect 20680 7692 20686 7704
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7528 2375 7531
rect 2498 7528 2504 7540
rect 2363 7500 2504 7528
rect 2363 7497 2375 7500
rect 2317 7491 2375 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4120 7500 5764 7528
rect 4120 7488 4126 7500
rect 2682 7420 2688 7472
rect 2740 7460 2746 7472
rect 3510 7460 3516 7472
rect 2740 7432 3516 7460
rect 2740 7420 2746 7432
rect 3510 7420 3516 7432
rect 3568 7420 3574 7472
rect 3694 7420 3700 7472
rect 3752 7460 3758 7472
rect 5736 7460 5764 7500
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 6178 7528 6184 7540
rect 5868 7500 6184 7528
rect 5868 7488 5874 7500
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 8018 7528 8024 7540
rect 7515 7500 8024 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 9122 7528 9128 7540
rect 8628 7500 9128 7528
rect 8628 7488 8634 7500
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 10428 7500 11652 7528
rect 10428 7460 10456 7500
rect 3752 7432 4108 7460
rect 5736 7432 10456 7460
rect 10505 7463 10563 7469
rect 3752 7420 3758 7432
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2648 7364 2881 7392
rect 2648 7352 2654 7364
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 3878 7392 3884 7404
rect 3839 7364 3884 7392
rect 2869 7355 2927 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 3050 7324 3056 7336
rect 1627 7296 3056 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 3476 7296 3709 7324
rect 3476 7284 3482 7296
rect 3697 7293 3709 7296
rect 3743 7293 3755 7327
rect 4080 7324 4108 7432
rect 10505 7429 10517 7463
rect 10551 7460 10563 7463
rect 10686 7460 10692 7472
rect 10551 7432 10692 7460
rect 10551 7429 10563 7432
rect 10505 7423 10563 7429
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 11624 7460 11652 7500
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12308 7500 17724 7528
rect 12308 7488 12314 7500
rect 13446 7460 13452 7472
rect 11624 7432 13452 7460
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 15565 7463 15623 7469
rect 15565 7429 15577 7463
rect 15611 7460 15623 7463
rect 16850 7460 16856 7472
rect 15611 7432 16856 7460
rect 15611 7429 15623 7432
rect 15565 7423 15623 7429
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 4798 7392 4804 7404
rect 4759 7364 4804 7392
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 7742 7392 7748 7404
rect 7208 7364 7748 7392
rect 7208 7324 7236 7364
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8938 7392 8944 7404
rect 8159 7364 8944 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 9122 7324 9128 7336
rect 4080 7296 7236 7324
rect 7300 7296 9128 7324
rect 3697 7287 3755 7293
rect 1857 7259 1915 7265
rect 1857 7225 1869 7259
rect 1903 7256 1915 7259
rect 3142 7256 3148 7268
rect 1903 7228 3148 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 5046 7259 5104 7265
rect 5046 7256 5058 7259
rect 3712 7228 5058 7256
rect 3712 7200 3740 7228
rect 5046 7225 5058 7228
rect 5092 7256 5104 7259
rect 5092 7228 6868 7256
rect 5092 7225 5104 7228
rect 5046 7219 5104 7225
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 3329 7191 3387 7197
rect 3329 7188 3341 7191
rect 2823 7160 3341 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 3329 7157 3341 7160
rect 3375 7157 3387 7191
rect 3329 7151 3387 7157
rect 3694 7148 3700 7200
rect 3752 7148 3758 7200
rect 3789 7191 3847 7197
rect 3789 7157 3801 7191
rect 3835 7188 3847 7191
rect 4154 7188 4160 7200
rect 3835 7160 4160 7188
rect 3835 7157 3847 7160
rect 3789 7151 3847 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 6638 7188 6644 7200
rect 4387 7160 6644 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 6840 7188 6868 7228
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 7300 7256 7328 7296
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9324 7324 9352 7355
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 9548 7364 10241 7392
rect 9548 7352 9554 7364
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12207 7364 13001 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 14516 7364 15700 7392
rect 14516 7352 14522 7364
rect 9582 7324 9588 7336
rect 9324 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 9674 7284 9680 7336
rect 9732 7284 9738 7336
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7324 10103 7327
rect 10502 7324 10508 7336
rect 10091 7296 10508 7324
rect 10091 7293 10103 7296
rect 10045 7287 10103 7293
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 10686 7324 10692 7336
rect 10647 7296 10692 7324
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 12768 7296 13461 7324
rect 12768 7284 12774 7296
rect 13449 7293 13461 7296
rect 13495 7293 13507 7327
rect 13449 7287 13507 7293
rect 13716 7327 13774 7333
rect 13716 7293 13728 7327
rect 13762 7324 13774 7327
rect 15194 7324 15200 7336
rect 13762 7296 15200 7324
rect 13762 7293 13774 7296
rect 13716 7287 13774 7293
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7324 15439 7327
rect 15562 7324 15568 7336
rect 15427 7296 15568 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 15672 7324 15700 7364
rect 16298 7352 16304 7404
rect 16356 7392 16362 7404
rect 16393 7395 16451 7401
rect 16393 7392 16405 7395
rect 16356 7364 16405 7392
rect 16356 7352 16362 7364
rect 16393 7361 16405 7364
rect 16439 7361 16451 7395
rect 16393 7355 16451 7361
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 17586 7392 17592 7404
rect 16540 7364 16585 7392
rect 17547 7364 17592 7392
rect 16540 7352 16546 7364
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17696 7392 17724 7500
rect 18874 7488 18880 7540
rect 18932 7528 18938 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 18932 7500 20085 7528
rect 18932 7488 18938 7500
rect 20073 7497 20085 7500
rect 20119 7497 20131 7531
rect 20073 7491 20131 7497
rect 20254 7488 20260 7540
rect 20312 7528 20318 7540
rect 20349 7531 20407 7537
rect 20349 7528 20361 7531
rect 20312 7500 20361 7528
rect 20312 7488 20318 7500
rect 20349 7497 20361 7500
rect 20395 7497 20407 7531
rect 20349 7491 20407 7497
rect 17696 7364 18828 7392
rect 16206 7324 16212 7336
rect 15672 7296 16212 7324
rect 16206 7284 16212 7296
rect 16264 7324 16270 7336
rect 17310 7324 17316 7336
rect 16264 7296 17172 7324
rect 17271 7296 17316 7324
rect 16264 7284 16270 7296
rect 6972 7228 7328 7256
rect 6972 7216 6978 7228
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 7929 7259 7987 7265
rect 7929 7256 7941 7259
rect 7616 7228 7941 7256
rect 7616 7216 7622 7228
rect 7929 7225 7941 7228
rect 7975 7225 7987 7259
rect 7929 7219 7987 7225
rect 8573 7259 8631 7265
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8619 7228 8800 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 7466 7188 7472 7200
rect 6840 7160 7472 7188
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7837 7191 7895 7197
rect 7837 7157 7849 7191
rect 7883 7188 7895 7191
rect 8294 7188 8300 7200
rect 7883 7160 8300 7188
rect 7883 7157 7895 7160
rect 7837 7151 7895 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 8662 7188 8668 7200
rect 8623 7160 8668 7188
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 8772 7188 8800 7228
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 9033 7259 9091 7265
rect 9033 7256 9045 7259
rect 8904 7228 9045 7256
rect 8904 7216 8910 7228
rect 9033 7225 9045 7228
rect 9079 7225 9091 7259
rect 9692 7256 9720 7284
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9692 7228 10149 7256
rect 9033 7219 9091 7225
rect 10137 7225 10149 7228
rect 10183 7256 10195 7259
rect 10410 7256 10416 7268
rect 10183 7228 10416 7256
rect 10183 7225 10195 7228
rect 10137 7219 10195 7225
rect 10410 7216 10416 7228
rect 10468 7216 10474 7268
rect 10594 7216 10600 7268
rect 10652 7256 10658 7268
rect 10956 7259 11014 7265
rect 10956 7256 10968 7259
rect 10652 7228 10968 7256
rect 10652 7216 10658 7228
rect 10956 7225 10968 7228
rect 11002 7256 11014 7259
rect 13998 7256 14004 7268
rect 11002 7228 14004 7256
rect 11002 7225 11014 7228
rect 10956 7219 11014 7225
rect 13998 7216 14004 7228
rect 14056 7216 14062 7268
rect 16301 7259 16359 7265
rect 16301 7225 16313 7259
rect 16347 7256 16359 7259
rect 17144 7256 17172 7296
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 18064 7256 18092 7287
rect 18506 7284 18512 7336
rect 18564 7324 18570 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18564 7296 18705 7324
rect 18564 7284 18570 7296
rect 18693 7293 18705 7296
rect 18739 7293 18751 7327
rect 18800 7324 18828 7364
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 20254 7392 20260 7404
rect 19852 7364 20260 7392
rect 19852 7352 19858 7364
rect 20254 7352 20260 7364
rect 20312 7392 20318 7404
rect 20901 7395 20959 7401
rect 20901 7392 20913 7395
rect 20312 7364 20913 7392
rect 20312 7352 20318 7364
rect 20901 7361 20913 7364
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 20809 7327 20867 7333
rect 18800 7296 20024 7324
rect 18693 7287 18751 7293
rect 16347 7228 16988 7256
rect 17144 7228 18092 7256
rect 18960 7259 19018 7265
rect 16347 7225 16359 7228
rect 16301 7219 16359 7225
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8772 7160 9137 7188
rect 9125 7157 9137 7160
rect 9171 7188 9183 7191
rect 9398 7188 9404 7200
rect 9171 7160 9404 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7188 9735 7191
rect 10042 7188 10048 7200
rect 9723 7160 10048 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10502 7188 10508 7200
rect 10463 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 11790 7148 11796 7200
rect 11848 7188 11854 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 11848 7160 12081 7188
rect 11848 7148 11854 7160
rect 12069 7157 12081 7160
rect 12115 7188 12127 7191
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 12115 7160 12173 7188
rect 12115 7157 12127 7160
rect 12069 7151 12127 7157
rect 12161 7157 12173 7160
rect 12207 7157 12219 7191
rect 12161 7151 12219 7157
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12676 7160 12817 7188
rect 12676 7148 12682 7160
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 12805 7151 12863 7157
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 14458 7188 14464 7200
rect 12943 7160 14464 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 14829 7191 14887 7197
rect 14829 7188 14841 7191
rect 14792 7160 14841 7188
rect 14792 7148 14798 7160
rect 14829 7157 14841 7160
rect 14875 7157 14887 7191
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 14829 7151 14887 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16960 7197 16988 7228
rect 18960 7225 18972 7259
rect 19006 7256 19018 7259
rect 19886 7256 19892 7268
rect 19006 7228 19892 7256
rect 19006 7225 19018 7228
rect 18960 7219 19018 7225
rect 19886 7216 19892 7228
rect 19944 7216 19950 7268
rect 16945 7191 17003 7197
rect 16945 7157 16957 7191
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 17405 7191 17463 7197
rect 17405 7157 17417 7191
rect 17451 7188 17463 7191
rect 18046 7188 18052 7200
rect 17451 7160 18052 7188
rect 17451 7157 17463 7160
rect 17405 7151 17463 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18233 7191 18291 7197
rect 18233 7157 18245 7191
rect 18279 7188 18291 7191
rect 19058 7188 19064 7200
rect 18279 7160 19064 7188
rect 18279 7157 18291 7160
rect 18233 7151 18291 7157
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 19996 7188 20024 7296
rect 20809 7293 20821 7327
rect 20855 7324 20867 7327
rect 21818 7324 21824 7336
rect 20855 7296 21824 7324
rect 20855 7293 20867 7296
rect 20809 7287 20867 7293
rect 21818 7284 21824 7296
rect 21876 7284 21882 7336
rect 20717 7259 20775 7265
rect 20717 7225 20729 7259
rect 20763 7256 20775 7259
rect 21910 7256 21916 7268
rect 20763 7228 21916 7256
rect 20763 7225 20775 7228
rect 20717 7219 20775 7225
rect 21910 7216 21916 7228
rect 21968 7216 21974 7268
rect 21082 7188 21088 7200
rect 19996 7160 21088 7188
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 3234 6984 3240 6996
rect 1964 6956 3240 6984
rect 1964 6860 1992 6956
rect 3234 6944 3240 6956
rect 3292 6944 3298 6996
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3878 6984 3884 6996
rect 3375 6956 3884 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 5258 6984 5264 6996
rect 4212 6956 5264 6984
rect 4212 6944 4218 6956
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 6178 6984 6184 6996
rect 5776 6956 6184 6984
rect 5776 6944 5782 6956
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 7469 6987 7527 6993
rect 7469 6953 7481 6987
rect 7515 6984 7527 6987
rect 7558 6984 7564 6996
rect 7515 6956 7564 6984
rect 7515 6953 7527 6956
rect 7469 6947 7527 6953
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7837 6987 7895 6993
rect 7837 6953 7849 6987
rect 7883 6984 7895 6987
rect 8662 6984 8668 6996
rect 7883 6956 8668 6984
rect 7883 6953 7895 6956
rect 7837 6947 7895 6953
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 8849 6987 8907 6993
rect 8849 6953 8861 6987
rect 8895 6984 8907 6987
rect 8938 6984 8944 6996
rect 8895 6956 8944 6984
rect 8895 6953 8907 6956
rect 8849 6947 8907 6953
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 9180 6956 10057 6984
rect 9180 6944 9186 6956
rect 10045 6953 10057 6956
rect 10091 6953 10103 6987
rect 10045 6947 10103 6953
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 10468 6956 13676 6984
rect 10468 6944 10474 6956
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 4433 6919 4491 6925
rect 4433 6916 4445 6919
rect 4396 6888 4445 6916
rect 4396 6876 4402 6888
rect 4433 6885 4445 6888
rect 4479 6885 4491 6919
rect 4433 6879 4491 6885
rect 5629 6919 5687 6925
rect 5629 6885 5641 6919
rect 5675 6916 5687 6919
rect 6086 6916 6092 6928
rect 5675 6888 6092 6916
rect 5675 6885 5687 6888
rect 5629 6879 5687 6885
rect 6086 6876 6092 6888
rect 6144 6916 6150 6928
rect 6546 6916 6552 6928
rect 6144 6888 6552 6916
rect 6144 6876 6150 6888
rect 6546 6876 6552 6888
rect 6604 6876 6610 6928
rect 6638 6876 6644 6928
rect 6696 6916 6702 6928
rect 12713 6919 12771 6925
rect 12713 6916 12725 6919
rect 6696 6888 12725 6916
rect 6696 6876 6702 6888
rect 12713 6885 12725 6888
rect 12759 6885 12771 6919
rect 12713 6879 12771 6885
rect 1946 6848 1952 6860
rect 1859 6820 1952 6848
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2216 6851 2274 6857
rect 2216 6817 2228 6851
rect 2262 6848 2274 6851
rect 2774 6848 2780 6860
rect 2262 6820 2780 6848
rect 2262 6817 2274 6820
rect 2216 6811 2274 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3292 6820 4660 6848
rect 3292 6808 3298 6820
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4632 6789 4660 6820
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6052 6820 9996 6848
rect 6052 6808 6058 6820
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4120 6752 4537 6780
rect 4120 6740 4126 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 6328 6752 6373 6780
rect 6328 6740 6334 6752
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6822 6780 6828 6792
rect 6696 6752 6828 6780
rect 6696 6740 6702 6752
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8159 6752 8892 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 2884 6684 5856 6712
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2884 6644 2912 6684
rect 1912 6616 2912 6644
rect 1912 6604 1918 6616
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3568 6616 4077 6644
rect 3568 6604 3574 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 5718 6644 5724 6656
rect 5679 6616 5724 6644
rect 4065 6607 4123 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 5828 6644 5856 6684
rect 6086 6672 6092 6724
rect 6144 6712 6150 6724
rect 7282 6712 7288 6724
rect 6144 6684 7288 6712
rect 6144 6672 6150 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 7944 6712 7972 6743
rect 8481 6715 8539 6721
rect 8481 6712 8493 6715
rect 7944 6684 8493 6712
rect 8481 6681 8493 6684
rect 8527 6681 8539 6715
rect 8864 6712 8892 6752
rect 8938 6740 8944 6792
rect 8996 6780 9002 6792
rect 9122 6780 9128 6792
rect 8996 6752 9041 6780
rect 9083 6752 9128 6780
rect 8996 6740 9002 6752
rect 9122 6740 9128 6752
rect 9180 6780 9186 6792
rect 9582 6780 9588 6792
rect 9180 6752 9588 6780
rect 9180 6740 9186 6752
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9490 6712 9496 6724
rect 8864 6684 9496 6712
rect 8481 6675 8539 6681
rect 9490 6672 9496 6684
rect 9548 6672 9554 6724
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 5828 6616 9689 6644
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 9968 6644 9996 6820
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 10956 6851 11014 6857
rect 10192 6820 10237 6848
rect 10192 6808 10198 6820
rect 10956 6817 10968 6851
rect 11002 6848 11014 6851
rect 11790 6848 11796 6860
rect 11002 6820 11796 6848
rect 11002 6817 11014 6820
rect 10956 6811 11014 6817
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 13648 6857 13676 6956
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 14553 6987 14611 6993
rect 14553 6984 14565 6987
rect 13780 6956 14565 6984
rect 13780 6944 13786 6956
rect 14553 6953 14565 6956
rect 14599 6984 14611 6987
rect 15838 6984 15844 6996
rect 14599 6956 15844 6984
rect 14599 6953 14611 6956
rect 14553 6947 14611 6953
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 16577 6987 16635 6993
rect 16577 6984 16589 6987
rect 15988 6956 16589 6984
rect 15988 6944 15994 6956
rect 16577 6953 16589 6956
rect 16623 6953 16635 6987
rect 16577 6947 16635 6953
rect 16945 6987 17003 6993
rect 16945 6953 16957 6987
rect 16991 6984 17003 6987
rect 18598 6984 18604 6996
rect 16991 6956 18604 6984
rect 16991 6953 17003 6956
rect 16945 6947 17003 6953
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 14645 6919 14703 6925
rect 14645 6885 14657 6919
rect 14691 6916 14703 6919
rect 15746 6916 15752 6928
rect 14691 6888 15752 6916
rect 14691 6885 14703 6888
rect 14645 6879 14703 6885
rect 13633 6851 13691 6857
rect 12584 6820 12940 6848
rect 12584 6808 12590 6820
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 10100 6752 10241 6780
rect 10100 6740 10106 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10686 6780 10692 6792
rect 10647 6752 10692 6780
rect 10229 6743 10287 6749
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 12912 6789 12940 6820
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 14660 6848 14688 6879
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 16114 6916 16120 6928
rect 15856 6888 16120 6916
rect 15590 6851 15648 6857
rect 13679 6820 14688 6848
rect 14752 6820 15516 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 11716 6752 12817 6780
rect 11716 6712 11744 6752
rect 12805 6749 12817 6752
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14752 6780 14780 6820
rect 13964 6752 14780 6780
rect 14829 6783 14887 6789
rect 13964 6740 13970 6752
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 15378 6780 15384 6792
rect 14875 6752 15384 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15488 6780 15516 6820
rect 15590 6817 15602 6851
rect 15636 6848 15648 6851
rect 15856 6848 15884 6888
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 16482 6916 16488 6928
rect 16443 6888 16488 6916
rect 16482 6876 16488 6888
rect 16540 6876 16546 6928
rect 16666 6876 16672 6928
rect 16724 6916 16730 6928
rect 17497 6919 17555 6925
rect 17497 6916 17509 6919
rect 16724 6888 17509 6916
rect 16724 6876 16730 6888
rect 17497 6885 17509 6888
rect 17543 6885 17555 6919
rect 17497 6879 17555 6885
rect 18874 6876 18880 6928
rect 18932 6916 18938 6928
rect 18932 6888 19003 6916
rect 18932 6876 18938 6888
rect 17402 6848 17408 6860
rect 15636 6820 15884 6848
rect 15939 6820 17408 6848
rect 15636 6817 15648 6820
rect 15590 6811 15648 6817
rect 15939 6780 15967 6820
rect 17402 6808 17408 6820
rect 17460 6848 17466 6860
rect 17589 6851 17647 6857
rect 17589 6848 17601 6851
rect 17460 6820 17601 6848
rect 17460 6808 17466 6820
rect 17589 6817 17601 6820
rect 17635 6817 17647 6851
rect 18506 6848 18512 6860
rect 18467 6820 18512 6848
rect 17589 6811 17647 6817
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 18782 6857 18788 6860
rect 18776 6811 18788 6857
rect 18840 6848 18846 6860
rect 18975 6848 19003 6888
rect 20165 6851 20223 6857
rect 20165 6848 20177 6851
rect 18840 6820 18876 6848
rect 18975 6820 20177 6848
rect 18782 6808 18788 6811
rect 18840 6808 18846 6820
rect 20165 6817 20177 6820
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 15488 6752 15967 6780
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 16669 6783 16727 6789
rect 16669 6780 16681 6783
rect 16356 6752 16681 6780
rect 16356 6740 16362 6752
rect 16669 6749 16681 6752
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 17736 6752 17781 6780
rect 17736 6740 17742 6752
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20772 6752 20913 6780
rect 20772 6740 20778 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 11624 6684 11744 6712
rect 11624 6644 11652 6684
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 14185 6715 14243 6721
rect 11940 6684 12204 6712
rect 11940 6672 11946 6684
rect 9968 6616 11652 6644
rect 9677 6607 9735 6613
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 11756 6616 12081 6644
rect 11756 6604 11762 6616
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12176 6644 12204 6684
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 16117 6715 16175 6721
rect 14231 6684 15700 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 15672 6656 15700 6684
rect 16117 6681 16129 6715
rect 16163 6712 16175 6715
rect 16945 6715 17003 6721
rect 16945 6712 16957 6715
rect 16163 6684 16957 6712
rect 16163 6681 16175 6684
rect 16117 6675 16175 6681
rect 16945 6681 16957 6684
rect 16991 6681 17003 6715
rect 16945 6675 17003 6681
rect 17129 6715 17187 6721
rect 17129 6681 17141 6715
rect 17175 6712 17187 6715
rect 17218 6712 17224 6724
rect 17175 6684 17224 6712
rect 17175 6681 17187 6684
rect 17129 6675 17187 6681
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 19886 6712 19892 6724
rect 19847 6684 19892 6712
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 12176 6616 12357 6644
rect 12069 6607 12127 6613
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 12345 6607 12403 6613
rect 13817 6647 13875 6653
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 15378 6644 15384 6656
rect 13863 6616 15384 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 15654 6604 15660 6656
rect 15712 6604 15718 6656
rect 15749 6647 15807 6653
rect 15749 6613 15761 6647
rect 15795 6644 15807 6647
rect 17770 6644 17776 6656
rect 15795 6616 17776 6644
rect 15795 6613 15807 6616
rect 15749 6607 15807 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18690 6644 18696 6656
rect 18104 6616 18696 6644
rect 18104 6604 18110 6616
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6644 20407 6647
rect 20898 6644 20904 6656
rect 20395 6616 20904 6644
rect 20395 6613 20407 6616
rect 20349 6607 20407 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3050 6440 3056 6452
rect 2832 6412 2877 6440
rect 3011 6412 3056 6440
rect 2832 6400 2838 6412
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 5810 6440 5816 6452
rect 4304 6412 5816 6440
rect 4304 6400 4310 6412
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6546 6400 6552 6452
rect 6604 6440 6610 6452
rect 8202 6440 8208 6452
rect 6604 6412 8208 6440
rect 6604 6400 6610 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 8352 6412 9597 6440
rect 8352 6400 8358 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 10410 6440 10416 6452
rect 9732 6412 10416 6440
rect 9732 6400 9738 6412
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6440 11115 6443
rect 15470 6440 15476 6452
rect 11103 6412 15476 6440
rect 11103 6409 11115 6412
rect 11057 6403 11115 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 16025 6443 16083 6449
rect 16025 6409 16037 6443
rect 16071 6440 16083 6443
rect 16482 6440 16488 6452
rect 16071 6412 16488 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 17678 6440 17684 6452
rect 16632 6412 17684 6440
rect 16632 6400 16638 6412
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 19061 6443 19119 6449
rect 19061 6409 19073 6443
rect 19107 6440 19119 6443
rect 20073 6443 20131 6449
rect 19107 6412 20024 6440
rect 19107 6409 19119 6412
rect 19061 6403 19119 6409
rect 2792 6372 2820 6400
rect 5445 6375 5503 6381
rect 2792 6344 3648 6372
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 3620 6313 3648 6344
rect 5445 6341 5457 6375
rect 5491 6372 5503 6375
rect 9309 6375 9367 6381
rect 5491 6344 7512 6372
rect 5491 6341 5503 6344
rect 5445 6335 5503 6341
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 1946 6236 1952 6248
rect 1443 6208 1952 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 3384 6208 4077 6236
rect 3384 6196 3390 6208
rect 4065 6205 4077 6208
rect 4111 6236 4123 6239
rect 4706 6236 4712 6248
rect 4111 6208 4712 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 5460 6236 5488 6335
rect 5810 6264 5816 6316
rect 5868 6304 5874 6316
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 5868 6276 6101 6304
rect 5868 6264 5874 6276
rect 6089 6273 6101 6276
rect 6135 6304 6147 6307
rect 6270 6304 6276 6316
rect 6135 6276 6276 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 6880 6276 7389 6304
rect 6880 6264 6886 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7484 6304 7512 6344
rect 9309 6341 9321 6375
rect 9355 6372 9367 6375
rect 9490 6372 9496 6384
rect 9355 6344 9496 6372
rect 9355 6341 9367 6344
rect 9309 6335 9367 6341
rect 9490 6332 9496 6344
rect 9548 6372 9554 6384
rect 9548 6344 10180 6372
rect 9548 6332 9554 6344
rect 10152 6313 10180 6344
rect 10686 6332 10692 6384
rect 10744 6372 10750 6384
rect 14277 6375 14335 6381
rect 10744 6344 12756 6372
rect 10744 6332 10750 6344
rect 10137 6307 10195 6313
rect 7484 6276 8064 6304
rect 7377 6267 7435 6273
rect 5994 6236 6000 6248
rect 4856 6208 5488 6236
rect 5955 6208 6000 6236
rect 4856 6196 4862 6208
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6205 7987 6239
rect 8036 6236 8064 6276
rect 10137 6273 10149 6307
rect 10183 6273 10195 6307
rect 11606 6304 11612 6316
rect 11567 6276 11612 6304
rect 10137 6267 10195 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 12728 6248 12756 6344
rect 14277 6341 14289 6375
rect 14323 6372 14335 6375
rect 15194 6372 15200 6384
rect 14323 6344 15200 6372
rect 14323 6341 14335 6344
rect 14277 6335 14335 6341
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 17586 6372 17592 6384
rect 15672 6344 17592 6372
rect 15672 6316 15700 6344
rect 17586 6332 17592 6344
rect 17644 6332 17650 6384
rect 18049 6375 18107 6381
rect 18049 6341 18061 6375
rect 18095 6372 18107 6375
rect 19996 6372 20024 6412
rect 20073 6409 20085 6443
rect 20119 6440 20131 6443
rect 20162 6440 20168 6452
rect 20119 6412 20168 6440
rect 20119 6409 20131 6412
rect 20073 6403 20131 6409
rect 20162 6400 20168 6412
rect 20220 6400 20226 6452
rect 20990 6372 20996 6384
rect 18095 6344 19564 6372
rect 19996 6344 20996 6372
rect 18095 6341 18107 6344
rect 18049 6335 18107 6341
rect 15654 6304 15660 6316
rect 15567 6276 15660 6304
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16172 6276 16528 6304
rect 16172 6264 16178 6276
rect 10042 6236 10048 6248
rect 8036 6208 10048 6236
rect 7929 6199 7987 6205
rect 1664 6171 1722 6177
rect 1664 6137 1676 6171
rect 1710 6168 1722 6171
rect 2314 6168 2320 6180
rect 1710 6140 2320 6168
rect 1710 6137 1722 6140
rect 1664 6131 1722 6137
rect 2314 6128 2320 6140
rect 2372 6128 2378 6180
rect 3878 6128 3884 6180
rect 3936 6168 3942 6180
rect 4246 6168 4252 6180
rect 3936 6140 4252 6168
rect 3936 6128 3942 6140
rect 4246 6128 4252 6140
rect 4304 6177 4310 6180
rect 4304 6171 4368 6177
rect 4304 6137 4322 6171
rect 4356 6137 4368 6171
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 4304 6131 4368 6137
rect 4448 6140 7297 6168
rect 4304 6128 4310 6131
rect 3418 6100 3424 6112
rect 3379 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4448 6100 4476 6140
rect 7285 6137 7297 6140
rect 7331 6137 7343 6171
rect 7285 6131 7343 6137
rect 5534 6100 5540 6112
rect 4028 6072 4476 6100
rect 5495 6072 5540 6100
rect 4028 6060 4034 6072
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6362 6100 6368 6112
rect 6323 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6696 6072 6837 6100
rect 6696 6060 6702 6072
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7742 6100 7748 6112
rect 7248 6072 7748 6100
rect 7248 6060 7254 6072
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 7944 6100 7972 6199
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 11238 6196 11244 6248
rect 11296 6236 11302 6248
rect 11425 6239 11483 6245
rect 11425 6236 11437 6239
rect 11296 6208 11437 6236
rect 11296 6196 11302 6208
rect 11425 6205 11437 6208
rect 11471 6205 11483 6239
rect 11425 6199 11483 6205
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 12434 6236 12440 6248
rect 11563 6208 12440 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 12897 6239 12955 6245
rect 12897 6236 12909 6239
rect 12768 6208 12909 6236
rect 12768 6196 12774 6208
rect 12897 6205 12909 6208
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 13164 6239 13222 6245
rect 13164 6205 13176 6239
rect 13210 6236 13222 6239
rect 14734 6236 14740 6248
rect 13210 6208 14740 6236
rect 13210 6205 13222 6208
rect 13164 6199 13222 6205
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6236 15531 6239
rect 15562 6236 15568 6248
rect 15519 6208 15568 6236
rect 15519 6205 15531 6208
rect 15473 6199 15531 6205
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 16390 6236 16396 6248
rect 16351 6208 16396 6236
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16500 6236 16528 6276
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 18693 6307 18751 6313
rect 16632 6276 16677 6304
rect 16632 6264 16638 6276
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 18782 6304 18788 6316
rect 18739 6276 18788 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 18782 6264 18788 6276
rect 18840 6304 18846 6316
rect 19334 6304 19340 6316
rect 18840 6276 19340 6304
rect 18840 6264 18846 6276
rect 19334 6264 19340 6276
rect 19392 6264 19398 6316
rect 19536 6313 19564 6344
rect 20990 6332 20996 6344
rect 21048 6332 21054 6384
rect 19521 6307 19579 6313
rect 19521 6273 19533 6307
rect 19567 6273 19579 6307
rect 19521 6267 19579 6273
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6304 19763 6307
rect 19886 6304 19892 6316
rect 19751 6276 19892 6304
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 20254 6264 20260 6316
rect 20312 6304 20318 6316
rect 20717 6307 20775 6313
rect 20717 6304 20729 6307
rect 20312 6276 20729 6304
rect 20312 6264 20318 6276
rect 20717 6273 20729 6276
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 17218 6236 17224 6248
rect 16500 6208 17224 6236
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 17402 6236 17408 6248
rect 17363 6208 17408 6236
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 19610 6196 19616 6248
rect 19668 6236 19674 6248
rect 20441 6239 20499 6245
rect 20441 6236 20453 6239
rect 19668 6208 20453 6236
rect 19668 6196 19674 6208
rect 20441 6205 20453 6208
rect 20487 6205 20499 6239
rect 20441 6199 20499 6205
rect 20530 6196 20536 6248
rect 20588 6236 20594 6248
rect 21085 6239 21143 6245
rect 20588 6208 20633 6236
rect 20588 6196 20594 6208
rect 21085 6205 21097 6239
rect 21131 6236 21143 6239
rect 21174 6236 21180 6248
rect 21131 6208 21180 6236
rect 21131 6205 21143 6208
rect 21085 6199 21143 6205
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 8202 6177 8208 6180
rect 8196 6168 8208 6177
rect 8163 6140 8208 6168
rect 8196 6131 8208 6140
rect 8202 6128 8208 6131
rect 8260 6128 8266 6180
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8352 6140 8524 6168
rect 8352 6128 8358 6140
rect 8386 6100 8392 6112
rect 7944 6072 8392 6100
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8496 6100 8524 6140
rect 8938 6128 8944 6180
rect 8996 6168 9002 6180
rect 18417 6171 18475 6177
rect 8996 6140 11284 6168
rect 8996 6128 9002 6140
rect 11256 6112 11284 6140
rect 15028 6140 16436 6168
rect 9582 6100 9588 6112
rect 8496 6072 9588 6100
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 9953 6103 10011 6109
rect 9953 6100 9965 6103
rect 9732 6072 9965 6100
rect 9732 6060 9738 6072
rect 9953 6069 9965 6072
rect 9999 6069 10011 6103
rect 9953 6063 10011 6069
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10597 6103 10655 6109
rect 10100 6072 10145 6100
rect 10100 6060 10106 6072
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 10778 6100 10784 6112
rect 10643 6072 10784 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11238 6060 11244 6112
rect 11296 6060 11302 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12158 6100 12164 6112
rect 11848 6072 12164 6100
rect 11848 6060 11854 6072
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 15028 6109 15056 6140
rect 15013 6103 15071 6109
rect 15013 6069 15025 6103
rect 15059 6069 15071 6103
rect 15013 6063 15071 6069
rect 15381 6103 15439 6109
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 15562 6100 15568 6112
rect 15427 6072 15568 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 15562 6060 15568 6072
rect 15620 6100 15626 6112
rect 16022 6100 16028 6112
rect 15620 6072 16028 6100
rect 15620 6060 15626 6072
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16408 6100 16436 6140
rect 18417 6137 18429 6171
rect 18463 6168 18475 6171
rect 18598 6168 18604 6180
rect 18463 6140 18604 6168
rect 18463 6137 18475 6140
rect 18417 6131 18475 6137
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 18782 6128 18788 6180
rect 18840 6168 18846 6180
rect 18840 6140 21312 6168
rect 18840 6128 18846 6140
rect 16485 6103 16543 6109
rect 16485 6100 16497 6103
rect 16408 6072 16497 6100
rect 16485 6069 16497 6072
rect 16531 6069 16543 6103
rect 16485 6063 16543 6069
rect 17589 6103 17647 6109
rect 17589 6069 17601 6103
rect 17635 6100 17647 6103
rect 18230 6100 18236 6112
rect 17635 6072 18236 6100
rect 17635 6069 17647 6072
rect 17589 6063 17647 6069
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 18690 6100 18696 6112
rect 18555 6072 18696 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 19426 6100 19432 6112
rect 19387 6072 19432 6100
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 21284 6109 21312 6140
rect 21269 6103 21327 6109
rect 21269 6069 21281 6103
rect 21315 6069 21327 6103
rect 21269 6063 21327 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 3234 5896 3240 5908
rect 2372 5868 3240 5896
rect 2372 5856 2378 5868
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 4062 5896 4068 5908
rect 4023 5868 4068 5896
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 5534 5896 5540 5908
rect 4479 5868 5540 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 5629 5899 5687 5905
rect 5629 5865 5641 5899
rect 5675 5896 5687 5899
rect 6086 5896 6092 5908
rect 5675 5868 6092 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 6457 5899 6515 5905
rect 6457 5896 6469 5899
rect 6420 5868 6469 5896
rect 6420 5856 6426 5868
rect 6457 5865 6469 5868
rect 6503 5865 6515 5899
rect 6457 5859 6515 5865
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 6730 5896 6736 5908
rect 6595 5868 6736 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7098 5856 7104 5908
rect 7156 5896 7162 5908
rect 7653 5899 7711 5905
rect 7653 5896 7665 5899
rect 7156 5868 7665 5896
rect 7156 5856 7162 5868
rect 7653 5865 7665 5868
rect 7699 5865 7711 5899
rect 7653 5859 7711 5865
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 10042 5896 10048 5908
rect 8619 5868 10048 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 11146 5896 11152 5908
rect 10468 5868 11152 5896
rect 10468 5856 10474 5868
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 11716 5868 15792 5896
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5828 4583 5831
rect 5718 5828 5724 5840
rect 4571 5800 5724 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 8294 5828 8300 5840
rect 6012 5800 8300 5828
rect 6012 5772 6040 5800
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 8941 5831 8999 5837
rect 8941 5797 8953 5831
rect 8987 5797 8999 5831
rect 10220 5831 10278 5837
rect 8941 5791 8999 5797
rect 9416 5800 9996 5828
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 1946 5760 1952 5772
rect 1903 5732 1952 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 2124 5763 2182 5769
rect 2124 5729 2136 5763
rect 2170 5760 2182 5763
rect 2590 5760 2596 5772
rect 2170 5732 2596 5760
rect 2170 5729 2182 5732
rect 2124 5723 2182 5729
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 5994 5760 6000 5772
rect 5583 5732 6000 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 7800 5732 7845 5760
rect 7800 5720 7806 5732
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 8947 5760 8975 5791
rect 8720 5732 8975 5760
rect 9033 5763 9091 5769
rect 8720 5720 8726 5732
rect 9033 5729 9045 5763
rect 9079 5760 9091 5763
rect 9306 5760 9312 5772
rect 9079 5732 9312 5760
rect 9079 5729 9091 5732
rect 9033 5723 9091 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4304 5664 4629 5692
rect 4304 5652 4310 5664
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 5810 5692 5816 5704
rect 5771 5664 5816 5692
rect 4617 5655 4675 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 6733 5655 6791 5661
rect 7760 5664 7849 5692
rect 6748 5624 6776 5655
rect 6822 5624 6828 5636
rect 6735 5596 6828 5624
rect 6822 5584 6828 5596
rect 6880 5624 6886 5636
rect 7760 5624 7788 5664
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 9122 5692 9128 5704
rect 8352 5664 9128 5692
rect 8352 5652 8358 5664
rect 9122 5652 9128 5664
rect 9180 5692 9186 5704
rect 9180 5664 9273 5692
rect 9180 5652 9186 5664
rect 6880 5596 7788 5624
rect 6880 5584 6886 5596
rect 7760 5568 7788 5596
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9416 5624 9444 5800
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9968 5769 9996 5800
rect 10220 5797 10232 5831
rect 10266 5828 10278 5831
rect 11606 5828 11612 5840
rect 10266 5800 11612 5828
rect 10266 5797 10278 5800
rect 10220 5791 10278 5797
rect 11606 5788 11612 5800
rect 11664 5788 11670 5840
rect 9953 5763 10011 5769
rect 9548 5732 9812 5760
rect 9548 5720 9554 5732
rect 9784 5692 9812 5732
rect 9953 5729 9965 5763
rect 9999 5729 10011 5763
rect 11716 5760 11744 5868
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 14185 5831 14243 5837
rect 14185 5828 14197 5831
rect 13872 5800 14197 5828
rect 13872 5788 13878 5800
rect 14185 5797 14197 5800
rect 14231 5797 14243 5831
rect 14185 5791 14243 5797
rect 14274 5788 14280 5840
rect 14332 5788 14338 5840
rect 15654 5837 15660 5840
rect 15648 5828 15660 5837
rect 15615 5800 15660 5828
rect 15648 5791 15660 5800
rect 15654 5788 15660 5791
rect 15712 5788 15718 5840
rect 15764 5828 15792 5868
rect 16390 5856 16396 5908
rect 16448 5896 16454 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 16448 5868 17049 5896
rect 16448 5856 16454 5868
rect 17037 5865 17049 5868
rect 17083 5865 17095 5899
rect 17037 5859 17095 5865
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 18288 5868 19288 5896
rect 18288 5856 18294 5868
rect 17494 5828 17500 5840
rect 15764 5800 17500 5828
rect 17494 5788 17500 5800
rect 17552 5788 17558 5840
rect 18776 5831 18834 5837
rect 18776 5797 18788 5831
rect 18822 5828 18834 5831
rect 18874 5828 18880 5840
rect 18822 5800 18880 5828
rect 18822 5797 18834 5800
rect 18776 5791 18834 5797
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 19260 5828 19288 5868
rect 19334 5856 19340 5908
rect 19392 5896 19398 5908
rect 19702 5896 19708 5908
rect 19392 5868 19708 5896
rect 19392 5856 19398 5868
rect 19702 5856 19708 5868
rect 19760 5896 19766 5908
rect 19889 5899 19947 5905
rect 19889 5896 19901 5899
rect 19760 5868 19901 5896
rect 19760 5856 19766 5868
rect 19889 5865 19901 5868
rect 19935 5865 19947 5899
rect 19889 5859 19947 5865
rect 19610 5828 19616 5840
rect 19260 5800 19616 5828
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 9953 5723 10011 5729
rect 10051 5732 11744 5760
rect 10051 5692 10079 5732
rect 11790 5720 11796 5772
rect 11848 5760 11854 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11848 5732 12081 5760
rect 11848 5720 11854 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 12161 5763 12219 5769
rect 12161 5729 12173 5763
rect 12207 5760 12219 5763
rect 12434 5760 12440 5772
rect 12207 5732 12440 5760
rect 12207 5729 12219 5732
rect 12161 5723 12219 5729
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 13078 5760 13084 5772
rect 13039 5732 13084 5760
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 13998 5760 14004 5772
rect 13280 5732 14004 5760
rect 9784 5664 10079 5692
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5692 12403 5695
rect 13170 5692 13176 5704
rect 12391 5664 13032 5692
rect 13131 5664 13176 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 8444 5596 9444 5624
rect 11701 5627 11759 5633
rect 8444 5584 8450 5596
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 12066 5624 12072 5636
rect 11747 5596 12072 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 12360 5596 12725 5624
rect 5166 5556 5172 5568
rect 5127 5528 5172 5556
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 6086 5556 6092 5568
rect 6047 5528 6092 5556
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 7190 5556 7196 5568
rect 7151 5528 7196 5556
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 7340 5528 7385 5556
rect 7340 5516 7346 5528
rect 7742 5516 7748 5568
rect 7800 5516 7806 5568
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 9582 5556 9588 5568
rect 7984 5528 9588 5556
rect 7984 5516 7990 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 10376 5528 11345 5556
rect 10376 5516 10382 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12360 5556 12388 5596
rect 12713 5593 12725 5596
rect 12759 5593 12771 5627
rect 13004 5624 13032 5664
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13280 5624 13308 5732
rect 13998 5720 14004 5732
rect 14056 5720 14062 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5760 14151 5763
rect 14292 5760 14320 5788
rect 14139 5732 14320 5760
rect 14139 5729 14151 5732
rect 14093 5723 14151 5729
rect 14642 5720 14648 5772
rect 14700 5760 14706 5772
rect 14918 5760 14924 5772
rect 14700 5732 14924 5760
rect 14700 5720 14706 5732
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 15528 5732 16865 5760
rect 15528 5720 15534 5732
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 17405 5763 17463 5769
rect 17405 5729 17417 5763
rect 17451 5760 17463 5763
rect 18049 5763 18107 5769
rect 18049 5760 18061 5763
rect 17451 5732 18061 5760
rect 17451 5729 17463 5732
rect 17405 5723 17463 5729
rect 18049 5729 18061 5732
rect 18095 5729 18107 5763
rect 18506 5760 18512 5772
rect 18467 5732 18512 5760
rect 18049 5723 18107 5729
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 20257 5763 20315 5769
rect 20257 5729 20269 5763
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5760 20959 5763
rect 21082 5760 21088 5772
rect 20947 5732 21088 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 14734 5692 14740 5704
rect 14323 5664 14357 5692
rect 14695 5664 14740 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 13004 5596 13308 5624
rect 13372 5624 13400 5655
rect 14292 5624 14320 5655
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 15381 5655 15439 5661
rect 14642 5624 14648 5636
rect 13372 5596 14648 5624
rect 12713 5587 12771 5593
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 11848 5528 12388 5556
rect 11848 5516 11854 5528
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 12492 5528 13737 5556
rect 12492 5516 12498 5528
rect 13725 5525 13737 5528
rect 13771 5525 13783 5559
rect 15396 5556 15424 5655
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 17644 5664 17689 5692
rect 17644 5652 17650 5664
rect 17862 5652 17868 5704
rect 17920 5692 17926 5704
rect 18524 5692 18552 5720
rect 17920 5664 18552 5692
rect 20272 5692 20300 5723
rect 21082 5720 21088 5732
rect 21140 5720 21146 5772
rect 21174 5692 21180 5704
rect 20272 5664 21180 5692
rect 17920 5652 17926 5664
rect 21174 5652 21180 5664
rect 21232 5652 21238 5704
rect 20441 5627 20499 5633
rect 20441 5593 20453 5627
rect 20487 5624 20499 5627
rect 21358 5624 21364 5636
rect 20487 5596 21364 5624
rect 20487 5593 20499 5596
rect 20441 5587 20499 5593
rect 21358 5584 21364 5596
rect 21416 5584 21422 5636
rect 15654 5556 15660 5568
rect 15396 5528 15660 5556
rect 13725 5519 13783 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 15746 5516 15752 5568
rect 15804 5556 15810 5568
rect 16390 5556 16396 5568
rect 15804 5528 16396 5556
rect 15804 5516 15810 5528
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 16482 5516 16488 5568
rect 16540 5556 16546 5568
rect 16761 5559 16819 5565
rect 16761 5556 16773 5559
rect 16540 5528 16773 5556
rect 16540 5516 16546 5528
rect 16761 5525 16773 5528
rect 16807 5525 16819 5559
rect 16761 5519 16819 5525
rect 16853 5559 16911 5565
rect 16853 5525 16865 5559
rect 16899 5556 16911 5559
rect 20990 5556 20996 5568
rect 16899 5528 20996 5556
rect 16899 5525 16911 5528
rect 16853 5519 16911 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 21085 5559 21143 5565
rect 21085 5525 21097 5559
rect 21131 5556 21143 5559
rect 21818 5556 21824 5568
rect 21131 5528 21824 5556
rect 21131 5525 21143 5528
rect 21085 5519 21143 5525
rect 21818 5516 21824 5528
rect 21876 5516 21882 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 3418 5352 3424 5364
rect 1995 5324 3424 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 8202 5352 8208 5364
rect 7524 5324 7788 5352
rect 8163 5324 8208 5352
rect 7524 5312 7530 5324
rect 7760 5284 7788 5324
rect 8202 5312 8208 5324
rect 8260 5352 8266 5364
rect 8294 5352 8300 5364
rect 8260 5324 8300 5352
rect 8260 5312 8266 5324
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 9030 5312 9036 5364
rect 9088 5312 9094 5364
rect 9306 5312 9312 5364
rect 9364 5352 9370 5364
rect 11977 5355 12035 5361
rect 9364 5324 11928 5352
rect 9364 5312 9370 5324
rect 8481 5287 8539 5293
rect 7760 5256 8340 5284
rect 8312 5228 8340 5256
rect 8481 5253 8493 5287
rect 8527 5253 8539 5287
rect 8481 5247 8539 5253
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 2501 5219 2559 5225
rect 2501 5216 2513 5219
rect 2372 5188 2513 5216
rect 2372 5176 2378 5188
rect 2501 5185 2513 5188
rect 2547 5185 2559 5219
rect 2501 5179 2559 5185
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 6273 5219 6331 5225
rect 6273 5185 6285 5219
rect 6319 5216 6331 5219
rect 6319 5188 6960 5216
rect 6319 5185 6331 5188
rect 6273 5179 6331 5185
rect 3160 5148 3188 5179
rect 3234 5148 3240 5160
rect 3160 5120 3240 5148
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 3412 5151 3470 5157
rect 3412 5117 3424 5151
rect 3458 5148 3470 5151
rect 4154 5148 4160 5160
rect 3458 5120 4160 5148
rect 3458 5117 3470 5120
rect 3412 5111 3470 5117
rect 4154 5108 4160 5120
rect 4212 5148 4218 5160
rect 5810 5148 5816 5160
rect 4212 5120 5816 5148
rect 4212 5108 4218 5120
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 6086 5148 6092 5160
rect 6047 5120 6092 5148
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6638 5148 6644 5160
rect 6227 5120 6644 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 6932 5148 6960 5188
rect 8294 5176 8300 5228
rect 8352 5176 8358 5228
rect 8496 5216 8524 5247
rect 9048 5216 9076 5312
rect 11790 5284 11796 5296
rect 11164 5256 11796 5284
rect 8496 5188 9076 5216
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9180 5188 9225 5216
rect 9180 5176 9186 5188
rect 9582 5176 9588 5228
rect 9640 5216 9646 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9640 5188 10241 5216
rect 9640 5176 9646 5188
rect 10229 5185 10241 5188
rect 10275 5216 10287 5219
rect 10318 5216 10324 5228
rect 10275 5188 10324 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 11164 5225 11192 5256
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 11900 5284 11928 5324
rect 11977 5321 11989 5355
rect 12023 5352 12035 5355
rect 15930 5352 15936 5364
rect 12023 5324 15936 5352
rect 12023 5321 12035 5324
rect 11977 5315 12035 5321
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 16356 5324 17049 5352
rect 16356 5312 16362 5324
rect 17037 5321 17049 5324
rect 17083 5321 17095 5355
rect 17037 5315 17095 5321
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 17494 5352 17500 5364
rect 17276 5324 17500 5352
rect 17276 5312 17282 5324
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 19153 5355 19211 5361
rect 19153 5321 19165 5355
rect 19199 5352 19211 5355
rect 19426 5352 19432 5364
rect 19199 5324 19432 5352
rect 19199 5321 19211 5324
rect 19153 5315 19211 5321
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 20162 5352 20168 5364
rect 20123 5324 20168 5352
rect 20162 5312 20168 5324
rect 20220 5352 20226 5364
rect 20220 5324 20852 5352
rect 20220 5312 20226 5324
rect 13078 5284 13084 5296
rect 11900 5256 13084 5284
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 14093 5287 14151 5293
rect 14093 5253 14105 5287
rect 14139 5284 14151 5287
rect 14277 5287 14335 5293
rect 14277 5284 14289 5287
rect 14139 5256 14289 5284
rect 14139 5253 14151 5256
rect 14093 5247 14151 5253
rect 14277 5253 14289 5256
rect 14323 5253 14335 5287
rect 14277 5247 14335 5253
rect 14826 5244 14832 5296
rect 14884 5284 14890 5296
rect 15470 5284 15476 5296
rect 14884 5256 15476 5284
rect 14884 5244 14890 5256
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 17589 5287 17647 5293
rect 17589 5253 17601 5287
rect 17635 5284 17647 5287
rect 20438 5284 20444 5296
rect 17635 5256 20444 5284
rect 17635 5253 17647 5256
rect 17589 5247 17647 5253
rect 20438 5244 20444 5256
rect 20496 5244 20502 5296
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 12066 5216 12072 5228
rect 11379 5188 12072 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 13538 5216 13544 5228
rect 12207 5188 13544 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 13817 5219 13875 5225
rect 13817 5216 13829 5219
rect 13688 5188 13829 5216
rect 13688 5176 13694 5188
rect 13817 5185 13829 5188
rect 13863 5185 13875 5219
rect 13817 5179 13875 5185
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15194 5216 15200 5228
rect 14967 5188 15200 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 15194 5176 15200 5188
rect 15252 5216 15258 5228
rect 18785 5219 18843 5225
rect 15252 5188 15424 5216
rect 15252 5176 15258 5188
rect 8849 5151 8907 5157
rect 6932 5120 7788 5148
rect 6825 5111 6883 5117
rect 2130 5040 2136 5092
rect 2188 5080 2194 5092
rect 2317 5083 2375 5089
rect 2317 5080 2329 5083
rect 2188 5052 2329 5080
rect 2188 5040 2194 5052
rect 2317 5049 2329 5052
rect 2363 5049 2375 5083
rect 2317 5043 2375 5049
rect 3142 5040 3148 5092
rect 3200 5080 3206 5092
rect 3602 5080 3608 5092
rect 3200 5052 3608 5080
rect 3200 5040 3206 5052
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 2406 5012 2412 5024
rect 2367 4984 2412 5012
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 4246 5012 4252 5024
rect 2648 4984 4252 5012
rect 2648 4972 2654 4984
rect 4246 4972 4252 4984
rect 4304 5012 4310 5024
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4304 4984 4537 5012
rect 4304 4972 4310 4984
rect 4525 4981 4537 4984
rect 4571 4981 4583 5015
rect 5718 5012 5724 5024
rect 5679 4984 5724 5012
rect 4525 4975 4583 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6840 5012 6868 5111
rect 7760 5092 7788 5120
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9490 5148 9496 5160
rect 8895 5120 9496 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 11054 5148 11060 5160
rect 10192 5120 11060 5148
rect 10192 5108 10198 5120
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 11790 5148 11796 5160
rect 11751 5120 11796 5148
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5148 12771 5151
rect 13725 5151 13783 5157
rect 12759 5120 13584 5148
rect 12759 5117 12771 5120
rect 12713 5111 12771 5117
rect 7098 5089 7104 5092
rect 7092 5080 7104 5089
rect 7059 5052 7104 5080
rect 7092 5043 7104 5052
rect 7098 5040 7104 5043
rect 7156 5040 7162 5092
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 7248 5052 7604 5080
rect 7248 5040 7254 5052
rect 7466 5012 7472 5024
rect 6840 4984 7472 5012
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 7576 5012 7604 5052
rect 7742 5040 7748 5092
rect 7800 5040 7806 5092
rect 9306 5080 9312 5092
rect 8404 5052 9312 5080
rect 8404 5012 8432 5052
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 10045 5083 10103 5089
rect 10045 5049 10057 5083
rect 10091 5080 10103 5083
rect 13354 5080 13360 5092
rect 10091 5052 13360 5080
rect 10091 5049 10103 5052
rect 10045 5043 10103 5049
rect 13354 5040 13360 5052
rect 13412 5040 13418 5092
rect 7576 4984 8432 5012
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 8996 4984 9041 5012
rect 8996 4972 9002 4984
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 9677 5015 9735 5021
rect 9677 5012 9689 5015
rect 9180 4984 9689 5012
rect 9180 4972 9186 4984
rect 9677 4981 9689 4984
rect 9723 4981 9735 5015
rect 9677 4975 9735 4981
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10410 5012 10416 5024
rect 10183 4984 10416 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10686 5012 10692 5024
rect 10647 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 11057 5015 11115 5021
rect 11057 4981 11069 5015
rect 11103 5012 11115 5015
rect 11330 5012 11336 5024
rect 11103 4984 11336 5012
rect 11103 4981 11115 4984
rect 11057 4975 11115 4981
rect 11330 4972 11336 4984
rect 11388 5012 11394 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 11388 4984 12173 5012
rect 11388 4972 11394 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12161 4975 12219 4981
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12676 4984 12909 5012
rect 12676 4972 12682 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 13078 4972 13084 5024
rect 13136 5012 13142 5024
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 13136 4984 13277 5012
rect 13136 4972 13142 4984
rect 13265 4981 13277 4984
rect 13311 4981 13323 5015
rect 13556 5012 13584 5120
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 14645 5151 14703 5157
rect 13771 5120 14596 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 13633 5083 13691 5089
rect 13633 5049 13645 5083
rect 13679 5080 13691 5083
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 13679 5052 14105 5080
rect 13679 5049 13691 5052
rect 13633 5043 13691 5049
rect 14093 5049 14105 5052
rect 14139 5049 14151 5083
rect 14568 5080 14596 5120
rect 14645 5117 14657 5151
rect 14691 5148 14703 5151
rect 14734 5148 14740 5160
rect 14691 5120 14740 5148
rect 14691 5117 14703 5120
rect 14645 5111 14703 5117
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 15286 5080 15292 5092
rect 14568 5052 15292 5080
rect 14093 5043 14151 5049
rect 15286 5040 15292 5052
rect 15344 5040 15350 5092
rect 15396 5080 15424 5188
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 19702 5216 19708 5228
rect 19663 5188 19708 5216
rect 18785 5179 18843 5185
rect 15654 5148 15660 5160
rect 15615 5120 15660 5148
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 15924 5151 15982 5157
rect 15924 5117 15936 5151
rect 15970 5148 15982 5151
rect 16482 5148 16488 5160
rect 15970 5120 16488 5148
rect 15970 5117 15982 5120
rect 15924 5111 15982 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 16666 5108 16672 5160
rect 16724 5148 16730 5160
rect 17405 5151 17463 5157
rect 17405 5148 17417 5151
rect 16724 5120 17417 5148
rect 16724 5108 16730 5120
rect 17405 5117 17417 5120
rect 17451 5117 17463 5151
rect 18506 5148 18512 5160
rect 18467 5120 18512 5148
rect 17405 5111 17463 5117
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 18800 5148 18828 5179
rect 19702 5176 19708 5188
rect 19760 5176 19766 5228
rect 20824 5225 20852 5324
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5185 20867 5219
rect 20990 5216 20996 5228
rect 20951 5188 20996 5216
rect 20809 5179 20867 5185
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 19334 5148 19340 5160
rect 18800 5120 19340 5148
rect 19334 5108 19340 5120
rect 19392 5148 19398 5160
rect 20162 5148 20168 5160
rect 19392 5120 20168 5148
rect 19392 5108 19398 5120
rect 20162 5108 20168 5120
rect 20220 5108 20226 5160
rect 20714 5148 20720 5160
rect 20675 5120 20720 5148
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 16022 5080 16028 5092
rect 15396 5052 16028 5080
rect 16022 5040 16028 5052
rect 16080 5040 16086 5092
rect 17954 5040 17960 5092
rect 18012 5080 18018 5092
rect 18601 5083 18659 5089
rect 18601 5080 18613 5083
rect 18012 5052 18613 5080
rect 18012 5040 18018 5052
rect 18601 5049 18613 5052
rect 18647 5049 18659 5083
rect 18601 5043 18659 5049
rect 19521 5083 19579 5089
rect 19521 5049 19533 5083
rect 19567 5080 19579 5083
rect 19567 5052 20392 5080
rect 19567 5049 19579 5052
rect 19521 5043 19579 5049
rect 13814 5012 13820 5024
rect 13556 4984 13820 5012
rect 13265 4975 13323 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14737 5015 14795 5021
rect 14737 5012 14749 5015
rect 14240 4984 14749 5012
rect 14240 4972 14246 4984
rect 14737 4981 14749 4984
rect 14783 4981 14795 5015
rect 14737 4975 14795 4981
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 16482 5012 16488 5024
rect 15528 4984 16488 5012
rect 15528 4972 15534 4984
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 18414 5012 18420 5024
rect 18187 4984 18420 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 19610 4972 19616 5024
rect 19668 5012 19674 5024
rect 20364 5021 20392 5052
rect 20349 5015 20407 5021
rect 19668 4984 19713 5012
rect 19668 4972 19674 4984
rect 20349 4981 20361 5015
rect 20395 4981 20407 5015
rect 20349 4975 20407 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2130 4808 2136 4820
rect 2091 4780 2136 4808
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 5166 4808 5172 4820
rect 4847 4780 5172 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 7340 4780 7573 4808
rect 7340 4768 7346 4780
rect 7561 4777 7573 4780
rect 7607 4777 7619 4811
rect 7561 4771 7619 4777
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 9030 4808 9036 4820
rect 7699 4780 9036 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9950 4808 9956 4820
rect 9723 4780 9956 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 11149 4811 11207 4817
rect 11149 4808 11161 4811
rect 10744 4780 11161 4808
rect 10744 4768 10750 4780
rect 11149 4777 11161 4780
rect 11195 4777 11207 4811
rect 11149 4771 11207 4777
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 15562 4808 15568 4820
rect 13504 4780 15568 4808
rect 13504 4768 13510 4780
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 17405 4811 17463 4817
rect 17405 4808 17417 4811
rect 15712 4780 17417 4808
rect 15712 4768 15718 4780
rect 2593 4743 2651 4749
rect 2593 4740 2605 4743
rect 2424 4712 2605 4740
rect 1762 4496 1768 4548
rect 1820 4536 1826 4548
rect 2424 4536 2452 4712
rect 2593 4709 2605 4712
rect 2639 4709 2651 4743
rect 2593 4703 2651 4709
rect 4709 4743 4767 4749
rect 4709 4709 4721 4743
rect 4755 4740 4767 4743
rect 9122 4740 9128 4752
rect 4755 4712 9128 4740
rect 4755 4709 4767 4712
rect 4709 4703 4767 4709
rect 9122 4700 9128 4712
rect 9180 4700 9186 4752
rect 10042 4740 10048 4752
rect 9955 4712 10048 4740
rect 10042 4700 10048 4712
rect 10100 4740 10106 4752
rect 10962 4740 10968 4752
rect 10100 4712 10968 4740
rect 10100 4700 10106 4712
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 14553 4743 14611 4749
rect 14553 4740 14565 4743
rect 12176 4712 14565 4740
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 3145 4675 3203 4681
rect 3145 4672 3157 4675
rect 2547 4644 3157 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 3145 4641 3157 4644
rect 3191 4641 3203 4675
rect 3145 4635 3203 4641
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 5793 4675 5851 4681
rect 5793 4672 5805 4675
rect 5684 4644 5805 4672
rect 5684 4632 5690 4644
rect 5793 4641 5805 4644
rect 5839 4641 5851 4675
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 5793 4635 5851 4641
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 10134 4672 10140 4684
rect 10095 4644 10140 4672
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 11054 4672 11060 4684
rect 11015 4644 11060 4672
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11330 4632 11336 4684
rect 11388 4672 11394 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 11388 4644 12081 4672
rect 11388 4632 11394 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 2682 4604 2688 4616
rect 2643 4576 2688 4604
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 4304 4576 4905 4604
rect 4304 4564 4310 4576
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 5350 4604 5356 4616
rect 5224 4576 5356 4604
rect 5224 4564 5230 4576
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 7742 4604 7748 4616
rect 6564 4576 7236 4604
rect 7703 4576 7748 4604
rect 2958 4536 2964 4548
rect 1820 4508 2964 4536
rect 1820 4496 1826 4508
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 4062 4428 4068 4480
rect 4120 4468 4126 4480
rect 6564 4468 6592 4576
rect 6917 4539 6975 4545
rect 6917 4505 6929 4539
rect 6963 4536 6975 4539
rect 7098 4536 7104 4548
rect 6963 4508 7104 4536
rect 6963 4505 6975 4508
rect 6917 4499 6975 4505
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 7208 4536 7236 4576
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 8478 4564 8484 4616
rect 8536 4604 8542 4616
rect 8662 4604 8668 4616
rect 8536 4576 8668 4604
rect 8536 4564 8542 4576
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 8846 4604 8852 4616
rect 8807 4576 8852 4604
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 10226 4604 10232 4616
rect 10187 4576 10232 4604
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11204 4576 11253 4604
rect 11204 4564 11210 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 9582 4536 9588 4548
rect 7208 4508 9588 4536
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 9950 4496 9956 4548
rect 10008 4536 10014 4548
rect 12176 4536 12204 4712
rect 14553 4709 14565 4712
rect 14599 4709 14611 4743
rect 14553 4703 14611 4709
rect 12888 4675 12946 4681
rect 12888 4641 12900 4675
rect 12934 4672 12946 4675
rect 12934 4644 13860 4672
rect 12934 4641 12946 4644
rect 12888 4635 12946 4641
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 12584 4576 12633 4604
rect 12584 4564 12590 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 13832 4604 13860 4644
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 13964 4644 14289 4672
rect 13964 4632 13970 4644
rect 14277 4641 14289 4644
rect 14323 4641 14335 4675
rect 14277 4635 14335 4641
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15746 4672 15752 4684
rect 15335 4644 15752 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 15856 4681 15884 4780
rect 17405 4777 17417 4780
rect 17451 4808 17463 4811
rect 17862 4808 17868 4820
rect 17451 4780 17868 4808
rect 17451 4777 17463 4780
rect 17405 4771 17463 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 19429 4811 19487 4817
rect 19429 4777 19441 4811
rect 19475 4808 19487 4811
rect 19610 4808 19616 4820
rect 19475 4780 19616 4808
rect 19475 4777 19487 4780
rect 19429 4771 19487 4777
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 16108 4743 16166 4749
rect 16108 4709 16120 4743
rect 16154 4740 16166 4743
rect 16298 4740 16304 4752
rect 16154 4712 16304 4740
rect 16154 4709 16166 4712
rect 16108 4703 16166 4709
rect 16298 4700 16304 4712
rect 16356 4700 16362 4752
rect 18414 4700 18420 4752
rect 18472 4740 18478 4752
rect 19889 4743 19947 4749
rect 19889 4740 19901 4743
rect 18472 4712 19901 4740
rect 18472 4700 18478 4712
rect 19889 4709 19901 4712
rect 19935 4709 19947 4743
rect 19889 4703 19947 4709
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4641 15899 4675
rect 17764 4675 17822 4681
rect 17764 4672 17776 4675
rect 15841 4635 15899 4641
rect 17236 4644 17776 4672
rect 15194 4604 15200 4616
rect 13832 4576 15200 4604
rect 12621 4567 12679 4573
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 17236 4548 17264 4644
rect 17764 4641 17776 4644
rect 17810 4672 17822 4675
rect 19334 4672 19340 4684
rect 17810 4644 19340 4672
rect 17810 4641 17822 4644
rect 17764 4635 17822 4641
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 19794 4672 19800 4684
rect 19755 4644 19800 4672
rect 19794 4632 19800 4644
rect 19852 4632 19858 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 21266 4672 21272 4684
rect 20947 4644 21272 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 17451 4576 17509 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 17497 4573 17509 4576
rect 17543 4573 17555 4607
rect 20073 4607 20131 4613
rect 20073 4604 20085 4607
rect 17497 4567 17555 4573
rect 18892 4576 20085 4604
rect 18892 4548 18920 4576
rect 20073 4573 20085 4576
rect 20119 4604 20131 4607
rect 20990 4604 20996 4616
rect 20119 4576 20996 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 10008 4508 12204 4536
rect 10008 4496 10014 4508
rect 14090 4496 14096 4548
rect 14148 4536 14154 4548
rect 15562 4536 15568 4548
rect 14148 4508 15568 4536
rect 14148 4496 14154 4508
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 17218 4536 17224 4548
rect 17131 4508 17224 4536
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 18874 4536 18880 4548
rect 18787 4508 18880 4536
rect 18874 4496 18880 4508
rect 18932 4496 18938 4548
rect 7190 4468 7196 4480
rect 4120 4440 6592 4468
rect 7151 4440 7196 4468
rect 4120 4428 4126 4440
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7650 4428 7656 4480
rect 7708 4468 7714 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 7708 4440 8217 4468
rect 7708 4428 7714 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 10689 4471 10747 4477
rect 10689 4468 10701 4471
rect 8352 4440 10701 4468
rect 8352 4428 8358 4440
rect 10689 4437 10701 4440
rect 10735 4437 10747 4471
rect 10689 4431 10747 4437
rect 12253 4471 12311 4477
rect 12253 4437 12265 4471
rect 12299 4468 12311 4471
rect 13538 4468 13544 4480
rect 12299 4440 13544 4468
rect 12299 4437 12311 4440
rect 12253 4431 12311 4437
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 14001 4471 14059 4477
rect 14001 4468 14013 4471
rect 13688 4440 14013 4468
rect 13688 4428 13694 4440
rect 14001 4437 14013 4440
rect 14047 4437 14059 4471
rect 14001 4431 14059 4437
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14826 4468 14832 4480
rect 14240 4440 14832 4468
rect 14240 4428 14246 4440
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 19334 4468 19340 4480
rect 15519 4440 19340 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 22738 4468 22744 4480
rect 21131 4440 22744 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 22738 4428 22744 4440
rect 22796 4428 22802 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 2406 4264 2412 4276
rect 2367 4236 2412 4264
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 7742 4264 7748 4276
rect 6380 4236 7748 4264
rect 2682 4156 2688 4208
rect 2740 4196 2746 4208
rect 2740 4168 3004 4196
rect 2740 4156 2746 4168
rect 2976 4137 3004 4168
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 3786 4088 3792 4140
rect 3844 4128 3850 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3844 4100 3893 4128
rect 3844 4088 3850 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4154 4128 4160 4140
rect 4111 4100 4160 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2866 4060 2872 4072
rect 2823 4032 2872 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3234 4020 3240 4072
rect 3292 4060 3298 4072
rect 4982 4060 4988 4072
rect 3292 4032 4988 4060
rect 3292 4020 3298 4032
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 5252 4063 5310 4069
rect 5252 4029 5264 4063
rect 5298 4060 5310 4063
rect 6380 4060 6408 4236
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 8846 4224 8852 4276
rect 8904 4224 8910 4276
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9493 4267 9551 4273
rect 9493 4264 9505 4267
rect 8996 4236 9505 4264
rect 8996 4224 9002 4236
rect 9493 4233 9505 4236
rect 9539 4233 9551 4267
rect 9493 4227 9551 4233
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 13446 4264 13452 4276
rect 9640 4236 13452 4264
rect 9640 4224 9646 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 13722 4264 13728 4276
rect 13556 4236 13728 4264
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 8864 4196 8892 4224
rect 9030 4196 9036 4208
rect 6788 4168 7420 4196
rect 8864 4168 9036 4196
rect 6788 4156 6794 4168
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7392 4137 7420 4168
rect 9030 4156 9036 4168
rect 9088 4196 9094 4208
rect 9217 4199 9275 4205
rect 9217 4196 9229 4199
rect 9088 4168 9229 4196
rect 9088 4156 9094 4168
rect 9217 4165 9229 4168
rect 9263 4165 9275 4199
rect 9217 4159 9275 4165
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 10321 4199 10379 4205
rect 9364 4168 10088 4196
rect 9364 4156 9370 4168
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 7248 4100 7297 4128
rect 7248 4088 7254 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7484 4100 7972 4128
rect 7484 4060 7512 4100
rect 5298 4032 6408 4060
rect 6472 4032 7512 4060
rect 7837 4063 7895 4069
rect 5298 4029 5310 4032
rect 5252 4023 5310 4029
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 4154 3992 4160 4004
rect 3835 3964 4160 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 4154 3952 4160 3964
rect 4212 3992 4218 4004
rect 5442 3992 5448 4004
rect 4212 3964 5448 3992
rect 4212 3952 4218 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 6472 3992 6500 4032
rect 7837 4029 7849 4063
rect 7883 4029 7895 4063
rect 7944 4060 7972 4100
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 9858 4128 9864 4140
rect 8904 4100 9864 4128
rect 8904 4088 8910 4100
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10060 4137 10088 4168
rect 10321 4165 10333 4199
rect 10367 4196 10379 4199
rect 10502 4196 10508 4208
rect 10367 4168 10508 4196
rect 10367 4165 10379 4168
rect 10321 4159 10379 4165
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 13556 4196 13584 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14642 4264 14648 4276
rect 14240 4236 14648 4264
rect 14240 4224 14246 4236
rect 14642 4224 14648 4236
rect 14700 4264 14706 4276
rect 15102 4264 15108 4276
rect 14700 4236 15108 4264
rect 14700 4224 14706 4236
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 15749 4267 15807 4273
rect 15749 4264 15761 4267
rect 15212 4236 15761 4264
rect 13280 4168 13584 4196
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 11146 4128 11152 4140
rect 11107 4100 11152 4128
rect 10045 4091 10103 4097
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 11790 4128 11796 4140
rect 11751 4100 11796 4128
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 13280 4137 13308 4168
rect 13630 4156 13636 4208
rect 13688 4196 13694 4208
rect 13688 4168 14320 4196
rect 13688 4156 13694 4168
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14292 4137 14320 4168
rect 14734 4156 14740 4208
rect 14792 4196 14798 4208
rect 15212 4196 15240 4236
rect 15749 4233 15761 4236
rect 15795 4233 15807 4267
rect 15749 4227 15807 4233
rect 15838 4224 15844 4276
rect 15896 4264 15902 4276
rect 19886 4264 19892 4276
rect 15896 4236 19892 4264
rect 15896 4224 15902 4236
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 14792 4168 15240 4196
rect 14792 4156 14798 4168
rect 15562 4156 15568 4208
rect 15620 4196 15626 4208
rect 15620 4168 16344 4196
rect 15620 4156 15626 4168
rect 14185 4131 14243 4137
rect 14185 4128 14197 4131
rect 14148 4100 14197 4128
rect 14148 4088 14154 4100
rect 14185 4097 14197 4100
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4097 14335 4131
rect 15102 4128 15108 4140
rect 15063 4100 15108 4128
rect 14277 4091 14335 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 16316 4137 16344 4168
rect 16390 4156 16396 4208
rect 16448 4196 16454 4208
rect 17862 4196 17868 4208
rect 16448 4168 17868 4196
rect 16448 4156 16454 4168
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 20254 4156 20260 4208
rect 20312 4196 20318 4208
rect 20312 4168 21036 4196
rect 20312 4156 20318 4168
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16942 4088 16948 4140
rect 17000 4128 17006 4140
rect 17126 4128 17132 4140
rect 17000 4100 17132 4128
rect 17000 4088 17006 4100
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17276 4100 17509 4128
rect 17276 4088 17282 4100
rect 17497 4097 17509 4100
rect 17543 4128 17555 4131
rect 17586 4128 17592 4140
rect 17543 4100 17592 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 18969 4131 19027 4137
rect 18969 4128 18981 4131
rect 18932 4100 18981 4128
rect 18932 4088 18938 4100
rect 18969 4097 18981 4100
rect 19015 4097 19027 4131
rect 18969 4091 19027 4097
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20162 4128 20168 4140
rect 20119 4100 20168 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 21008 4137 21036 4168
rect 20901 4131 20959 4137
rect 20901 4128 20913 4131
rect 20864 4100 20913 4128
rect 20864 4088 20870 4100
rect 20901 4097 20913 4100
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4097 21051 4131
rect 20993 4091 21051 4097
rect 7944 4032 9444 4060
rect 7837 4023 7895 4029
rect 7374 3992 7380 4004
rect 5552 3964 6500 3992
rect 6840 3964 7380 3992
rect 2869 3927 2927 3933
rect 2869 3893 2881 3927
rect 2915 3924 2927 3927
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 2915 3896 3433 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 3421 3893 3433 3896
rect 3467 3893 3479 3927
rect 3421 3887 3479 3893
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 5552 3924 5580 3964
rect 3660 3896 5580 3924
rect 3660 3884 3666 3896
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5684 3896 6377 3924
rect 5684 3884 5690 3896
rect 6365 3893 6377 3896
rect 6411 3924 6423 3927
rect 6730 3924 6736 3936
rect 6411 3896 6736 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 6840 3933 6868 3964
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 7852 3992 7880 4023
rect 7524 3964 7880 3992
rect 8104 3995 8162 4001
rect 7524 3952 7530 3964
rect 8104 3961 8116 3995
rect 8150 3992 8162 3995
rect 9306 3992 9312 4004
rect 8150 3964 9312 3992
rect 8150 3961 8162 3964
rect 8104 3955 8162 3961
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 9416 3992 9444 4032
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9824 4032 9965 4060
rect 9824 4020 9830 4032
rect 9953 4029 9965 4032
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 10928 4032 11621 4060
rect 10928 4020 10934 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11900 4060 11928 4088
rect 13078 4060 13084 4072
rect 11609 4023 11667 4029
rect 11716 4032 11928 4060
rect 13039 4032 13084 4060
rect 11716 3992 11744 4032
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 13228 4032 14596 4060
rect 13228 4020 13234 4032
rect 9416 3964 11744 3992
rect 11882 3952 11888 4004
rect 11940 3992 11946 4004
rect 14568 3992 14596 4032
rect 17310 4020 17316 4072
rect 17368 4060 17374 4072
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 17368 4032 17785 4060
rect 17368 4020 17374 4032
rect 17773 4029 17785 4032
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 19797 4063 19855 4069
rect 19797 4060 19809 4063
rect 18104 4032 19809 4060
rect 18104 4020 18110 4032
rect 19797 4029 19809 4032
rect 19843 4029 19855 4063
rect 19797 4023 19855 4029
rect 14918 3992 14924 4004
rect 11940 3964 14228 3992
rect 14568 3964 14688 3992
rect 14879 3964 14924 3992
rect 11940 3952 11946 3964
rect 6825 3927 6883 3933
rect 6825 3893 6837 3927
rect 6871 3893 6883 3927
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 6825 3887 6883 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 9907 3896 10333 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 10321 3887 10379 3893
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10870 3924 10876 3936
rect 10831 3896 10876 3924
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11238 3924 11244 3936
rect 11011 3896 11244 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 12710 3924 12716 3936
rect 12671 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 13173 3927 13231 3933
rect 13173 3893 13185 3927
rect 13219 3924 13231 3927
rect 13725 3927 13783 3933
rect 13725 3924 13737 3927
rect 13219 3896 13737 3924
rect 13219 3893 13231 3896
rect 13173 3887 13231 3893
rect 13725 3893 13737 3896
rect 13771 3893 13783 3927
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 13725 3887 13783 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14200 3924 14228 3964
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 14200 3896 14565 3924
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 14660 3924 14688 3964
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 15010 3952 15016 4004
rect 15068 3992 15074 4004
rect 15068 3964 15113 3992
rect 15068 3952 15074 3964
rect 15194 3952 15200 4004
rect 15252 3992 15258 4004
rect 15565 3995 15623 4001
rect 15565 3992 15577 3995
rect 15252 3964 15577 3992
rect 15252 3952 15258 3964
rect 15565 3961 15577 3964
rect 15611 3992 15623 3995
rect 16117 3995 16175 4001
rect 16117 3992 16129 3995
rect 15611 3964 16129 3992
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 16117 3961 16129 3964
rect 16163 3961 16175 3995
rect 18785 3995 18843 4001
rect 18785 3992 18797 3995
rect 16117 3955 16175 3961
rect 16960 3964 18797 3992
rect 16960 3933 16988 3964
rect 18785 3961 18797 3964
rect 18831 3961 18843 3995
rect 19812 3992 19840 4023
rect 20990 3992 20996 4004
rect 19812 3964 20996 3992
rect 18785 3955 18843 3961
rect 20990 3952 20996 3964
rect 21048 3952 21054 4004
rect 16209 3927 16267 3933
rect 16209 3924 16221 3927
rect 14660 3896 16221 3924
rect 14553 3887 14611 3893
rect 16209 3893 16221 3896
rect 16255 3893 16267 3927
rect 16209 3887 16267 3893
rect 16945 3927 17003 3933
rect 16945 3893 16957 3927
rect 16991 3893 17003 3927
rect 17310 3924 17316 3936
rect 17271 3896 17316 3924
rect 16945 3887 17003 3893
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17405 3927 17463 3933
rect 17405 3893 17417 3927
rect 17451 3924 17463 3927
rect 17773 3927 17831 3933
rect 17773 3924 17785 3927
rect 17451 3896 17785 3924
rect 17451 3893 17463 3896
rect 17405 3887 17463 3893
rect 17773 3893 17785 3896
rect 17819 3924 17831 3927
rect 18230 3924 18236 3936
rect 17819 3896 18236 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18417 3927 18475 3933
rect 18417 3893 18429 3927
rect 18463 3924 18475 3927
rect 18598 3924 18604 3936
rect 18463 3896 18604 3924
rect 18463 3893 18475 3896
rect 18417 3887 18475 3893
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 18877 3927 18935 3933
rect 18877 3893 18889 3927
rect 18923 3924 18935 3927
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 18923 3896 19441 3924
rect 18923 3893 18935 3896
rect 18877 3887 18935 3893
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19429 3887 19487 3893
rect 19794 3884 19800 3936
rect 19852 3924 19858 3936
rect 19889 3927 19947 3933
rect 19889 3924 19901 3927
rect 19852 3896 19901 3924
rect 19852 3884 19858 3896
rect 19889 3893 19901 3896
rect 19935 3893 19947 3927
rect 19889 3887 19947 3893
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20036 3896 20453 3924
rect 20036 3884 20042 3896
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20806 3924 20812 3936
rect 20767 3896 20812 3924
rect 20441 3887 20499 3893
rect 20806 3884 20812 3896
rect 20864 3884 20870 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5718 3720 5724 3732
rect 5215 3692 5724 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6086 3720 6092 3732
rect 6012 3692 6092 3720
rect 2317 3655 2375 3661
rect 2317 3621 2329 3655
rect 2363 3652 2375 3655
rect 2869 3655 2927 3661
rect 2869 3652 2881 3655
rect 2363 3624 2881 3652
rect 2363 3621 2375 3624
rect 2317 3615 2375 3621
rect 2869 3621 2881 3624
rect 2915 3621 2927 3655
rect 2869 3615 2927 3621
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 3234 3584 3240 3596
rect 2455 3556 3240 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 3329 3587 3387 3593
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 3602 3584 3608 3596
rect 3375 3556 3608 3584
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5534 3584 5540 3596
rect 5040 3556 5540 3584
rect 5040 3544 5046 3556
rect 5534 3544 5540 3556
rect 5592 3584 5598 3596
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 5592 3556 5825 3584
rect 5592 3544 5598 3556
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 6012 3584 6040 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 6880 3692 10824 3720
rect 6880 3680 6886 3692
rect 6178 3612 6184 3664
rect 6236 3652 6242 3664
rect 10502 3652 10508 3664
rect 6236 3624 10508 3652
rect 6236 3612 6242 3624
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 10796 3652 10824 3692
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11425 3723 11483 3729
rect 11425 3720 11437 3723
rect 10928 3692 11437 3720
rect 10928 3680 10934 3692
rect 11425 3689 11437 3692
rect 11471 3689 11483 3723
rect 11882 3720 11888 3732
rect 11843 3692 11888 3720
rect 11425 3683 11483 3689
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 13170 3720 13176 3732
rect 12636 3692 13176 3720
rect 12636 3652 12664 3692
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 13722 3720 13728 3732
rect 13320 3692 13728 3720
rect 13320 3680 13326 3692
rect 13722 3680 13728 3692
rect 13780 3720 13786 3732
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 13780 3692 14197 3720
rect 13780 3680 13786 3692
rect 14185 3689 14197 3692
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 14274 3680 14280 3732
rect 14332 3720 14338 3732
rect 15286 3720 15292 3732
rect 14332 3692 14596 3720
rect 15247 3692 15292 3720
rect 14332 3680 14338 3692
rect 10796 3624 12664 3652
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 14568 3652 14596 3692
rect 15286 3680 15292 3692
rect 15344 3680 15350 3732
rect 15654 3720 15660 3732
rect 15615 3692 15660 3720
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 17034 3720 17040 3732
rect 16632 3692 16896 3720
rect 16995 3692 17040 3720
rect 16632 3680 16638 3692
rect 16758 3652 16764 3664
rect 12768 3624 14504 3652
rect 14568 3624 16764 3652
rect 12768 3612 12774 3624
rect 6069 3587 6127 3593
rect 6069 3584 6081 3587
rect 6012 3556 6081 3584
rect 5813 3547 5871 3553
rect 6069 3553 6081 3556
rect 6115 3553 6127 3587
rect 6069 3547 6127 3553
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 8185 3587 8243 3593
rect 8185 3584 8197 3587
rect 7340 3556 8197 3584
rect 7340 3544 7346 3556
rect 8185 3553 8197 3556
rect 8231 3584 8243 3587
rect 9858 3584 9864 3596
rect 8231 3556 9864 3584
rect 8231 3553 8243 3556
rect 8185 3547 8243 3553
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 10036 3587 10094 3593
rect 10036 3553 10048 3587
rect 10082 3584 10094 3587
rect 11793 3587 11851 3593
rect 10082 3556 11376 3584
rect 10082 3553 10094 3556
rect 10036 3547 10094 3553
rect 2590 3516 2596 3528
rect 2551 3488 2596 3516
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3016 3488 3433 3516
rect 3016 3476 3022 3488
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3970 3516 3976 3528
rect 3559 3488 3976 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 5258 3516 5264 3528
rect 5219 3488 5264 3516
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5626 3516 5632 3528
rect 5491 3488 5632 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7926 3516 7932 3528
rect 7524 3488 7932 3516
rect 7524 3476 7530 3488
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 9766 3516 9772 3528
rect 9727 3488 9772 3516
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 11348 3516 11376 3556
rect 11793 3553 11805 3587
rect 11839 3584 11851 3587
rect 12618 3584 12624 3596
rect 11839 3556 12624 3584
rect 11839 3553 11851 3556
rect 11793 3547 11851 3553
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 13072 3587 13130 3593
rect 13072 3553 13084 3587
rect 13118 3584 13130 3587
rect 13630 3584 13636 3596
rect 13118 3556 13636 3584
rect 13118 3553 13130 3556
rect 13072 3547 13130 3553
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 14476 3593 14504 3624
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 16868 3652 16896 3692
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 18509 3723 18567 3729
rect 17420 3692 18000 3720
rect 16945 3655 17003 3661
rect 16945 3652 16957 3655
rect 16868 3624 16957 3652
rect 16945 3621 16957 3624
rect 16991 3621 17003 3655
rect 17420 3652 17448 3692
rect 16945 3615 17003 3621
rect 17052 3624 17448 3652
rect 14461 3587 14519 3593
rect 14461 3553 14473 3587
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 17052 3584 17080 3624
rect 17494 3612 17500 3664
rect 17552 3652 17558 3664
rect 17865 3655 17923 3661
rect 17865 3652 17877 3655
rect 17552 3624 17877 3652
rect 17552 3612 17558 3624
rect 17865 3621 17877 3624
rect 17911 3621 17923 3655
rect 17972 3652 18000 3692
rect 18509 3689 18521 3723
rect 18555 3720 18567 3723
rect 18690 3720 18696 3732
rect 18555 3692 18696 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 18877 3723 18935 3729
rect 18877 3689 18889 3723
rect 18923 3720 18935 3723
rect 19521 3723 19579 3729
rect 19521 3720 19533 3723
rect 18923 3692 19533 3720
rect 18923 3689 18935 3692
rect 18877 3683 18935 3689
rect 19521 3689 19533 3692
rect 19567 3689 19579 3723
rect 19521 3683 19579 3689
rect 19981 3655 20039 3661
rect 19981 3652 19993 3655
rect 17972 3624 19993 3652
rect 17865 3615 17923 3621
rect 19981 3621 19993 3624
rect 20027 3621 20039 3655
rect 21174 3652 21180 3664
rect 21135 3624 21180 3652
rect 19981 3615 20039 3621
rect 21174 3612 21180 3624
rect 21232 3612 21238 3664
rect 16724 3556 17080 3584
rect 17589 3587 17647 3593
rect 16724 3544 16730 3556
rect 17589 3553 17601 3587
rect 17635 3584 17647 3587
rect 17678 3584 17684 3596
rect 17635 3556 17684 3584
rect 17635 3553 17647 3556
rect 17589 3547 17647 3553
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 18874 3544 18880 3596
rect 18932 3584 18938 3596
rect 19889 3587 19947 3593
rect 18932 3556 19104 3584
rect 18932 3544 18938 3556
rect 12066 3516 12072 3528
rect 11348 3488 12072 3516
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 12802 3516 12808 3528
rect 12584 3488 12808 3516
rect 12584 3476 12590 3488
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 13872 3488 14657 3516
rect 13872 3476 13878 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 15746 3516 15752 3528
rect 15707 3488 15752 3516
rect 14645 3479 14703 3485
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16022 3516 16028 3528
rect 15979 3488 16028 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 17221 3519 17279 3525
rect 17221 3485 17233 3519
rect 17267 3516 17279 3519
rect 17494 3516 17500 3528
rect 17267 3488 17500 3516
rect 17267 3485 17279 3488
rect 17221 3479 17279 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 19076 3525 19104 3556
rect 19889 3553 19901 3587
rect 19935 3584 19947 3587
rect 20346 3584 20352 3596
rect 19935 3556 20352 3584
rect 19935 3553 19947 3556
rect 19889 3547 19947 3553
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 21082 3584 21088 3596
rect 20947 3556 21088 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 18969 3519 19027 3525
rect 18969 3485 18981 3519
rect 19015 3485 19027 3519
rect 18969 3479 19027 3485
rect 19061 3519 19119 3525
rect 19061 3485 19073 3519
rect 19107 3485 19119 3519
rect 20162 3516 20168 3528
rect 20123 3488 20168 3516
rect 19061 3479 19119 3485
rect 1946 3448 1952 3460
rect 1907 3420 1952 3448
rect 1946 3408 1952 3420
rect 2004 3408 2010 3460
rect 2869 3451 2927 3457
rect 2869 3417 2881 3451
rect 2915 3448 2927 3451
rect 9306 3448 9312 3460
rect 2915 3420 5856 3448
rect 2915 3417 2927 3420
rect 2869 3411 2927 3417
rect 2961 3383 3019 3389
rect 2961 3349 2973 3383
rect 3007 3380 3019 3383
rect 3050 3380 3056 3392
rect 3007 3352 3056 3380
rect 3007 3349 3019 3352
rect 2961 3343 3019 3349
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 5718 3380 5724 3392
rect 4847 3352 5724 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 5828 3380 5856 3420
rect 6748 3420 7880 3448
rect 9267 3420 9312 3448
rect 6748 3380 6776 3420
rect 5828 3352 6776 3380
rect 7193 3383 7251 3389
rect 7193 3349 7205 3383
rect 7239 3380 7251 3383
rect 7282 3380 7288 3392
rect 7239 3352 7288 3380
rect 7239 3349 7251 3352
rect 7193 3343 7251 3349
rect 7282 3340 7288 3352
rect 7340 3380 7346 3392
rect 7742 3380 7748 3392
rect 7340 3352 7748 3380
rect 7340 3340 7346 3352
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 7852 3380 7880 3420
rect 9306 3408 9312 3420
rect 9364 3408 9370 3460
rect 15194 3408 15200 3460
rect 15252 3448 15258 3460
rect 16206 3448 16212 3460
rect 15252 3420 16212 3448
rect 15252 3408 15258 3420
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 16577 3451 16635 3457
rect 16577 3417 16589 3451
rect 16623 3448 16635 3451
rect 18984 3448 19012 3479
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 16623 3420 19012 3448
rect 16623 3417 16635 3420
rect 16577 3411 16635 3417
rect 8294 3380 8300 3392
rect 7852 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 11146 3380 11152 3392
rect 11107 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 13170 3380 13176 3392
rect 11756 3352 13176 3380
rect 11756 3340 11762 3352
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 17218 3380 17224 3392
rect 13596 3352 17224 3380
rect 13596 3340 13602 3352
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3050 3136 3056 3188
rect 3108 3176 3114 3188
rect 3108 3148 4936 3176
rect 3108 3136 3114 3148
rect 4908 3108 4936 3148
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5316 3148 5641 3176
rect 5316 3136 5322 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 6914 3176 6920 3188
rect 5629 3139 5687 3145
rect 5736 3148 6920 3176
rect 5736 3108 5764 3148
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7190 3176 7196 3188
rect 7151 3148 7196 3176
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 9766 3176 9772 3188
rect 7984 3148 9772 3176
rect 7984 3136 7990 3148
rect 7282 3108 7288 3120
rect 4908 3080 5764 3108
rect 6196 3080 7288 3108
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3694 3040 3700 3052
rect 3651 3012 3700 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 6196 3049 6224 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3009 6239 3043
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 6181 3003 6239 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8570 3040 8576 3052
rect 7800 3012 7845 3040
rect 8496 3012 8576 3040
rect 7800 3000 7806 3012
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 3973 2975 4031 2981
rect 3476 2944 3521 2972
rect 3476 2932 3482 2944
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4982 2972 4988 2984
rect 4019 2944 4988 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 8496 2972 8524 3012
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 8680 3049 8708 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9916 3148 10057 3176
rect 9916 3136 9922 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 11885 3179 11943 3185
rect 10045 3139 10103 3145
rect 10428 3148 11836 3176
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 10428 2972 10456 3148
rect 11808 3108 11836 3148
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12066 3176 12072 3188
rect 11931 3148 12072 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12360 3148 14044 3176
rect 12360 3108 12388 3148
rect 11808 3080 12388 3108
rect 14016 3040 14044 3148
rect 14090 3136 14096 3188
rect 14148 3176 14154 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 14148 3148 15301 3176
rect 14148 3136 14154 3148
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 15289 3139 15347 3145
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 16485 3179 16543 3185
rect 16485 3176 16497 3179
rect 15804 3148 16497 3176
rect 15804 3136 15810 3148
rect 16485 3145 16497 3148
rect 16531 3145 16543 3179
rect 16485 3139 16543 3145
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 18690 3176 18696 3188
rect 17184 3148 18696 3176
rect 17184 3136 17190 3148
rect 18690 3136 18696 3148
rect 18748 3136 18754 3188
rect 20441 3179 20499 3185
rect 20441 3145 20453 3179
rect 20487 3176 20499 3179
rect 20806 3176 20812 3188
rect 20487 3148 20812 3176
rect 20487 3145 20499 3148
rect 20441 3139 20499 3145
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 14458 3108 14464 3120
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 16298 3108 16304 3120
rect 16259 3080 16304 3108
rect 16298 3068 16304 3080
rect 16356 3108 16362 3120
rect 16356 3080 16436 3108
rect 16356 3068 16362 3080
rect 15105 3043 15163 3049
rect 14016 3012 14780 3040
rect 5368 2944 8524 2972
rect 8588 2944 10456 2972
rect 10505 2975 10563 2981
rect 1946 2864 1952 2916
rect 2004 2904 2010 2916
rect 4246 2913 4252 2916
rect 2004 2876 4016 2904
rect 2004 2864 2010 2876
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 3329 2839 3387 2845
rect 3329 2836 3341 2839
rect 3292 2808 3341 2836
rect 3292 2796 3298 2808
rect 3329 2805 3341 2808
rect 3375 2836 3387 2839
rect 3510 2836 3516 2848
rect 3375 2808 3516 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 3988 2836 4016 2876
rect 4240 2867 4252 2913
rect 4304 2904 4310 2916
rect 4304 2876 4340 2904
rect 4246 2864 4252 2867
rect 4304 2864 4310 2876
rect 5258 2836 5264 2848
rect 3988 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5368 2845 5396 2944
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 6089 2907 6147 2913
rect 6089 2904 6101 2907
rect 5592 2876 6101 2904
rect 5592 2864 5598 2876
rect 6089 2873 6101 2876
rect 6135 2873 6147 2907
rect 6089 2867 6147 2873
rect 7561 2907 7619 2913
rect 7561 2873 7573 2907
rect 7607 2904 7619 2907
rect 8202 2904 8208 2916
rect 7607 2876 8208 2904
rect 7607 2873 7619 2876
rect 7561 2867 7619 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 5353 2839 5411 2845
rect 5353 2805 5365 2839
rect 5399 2805 5411 2839
rect 5994 2836 6000 2848
rect 5955 2808 6000 2836
rect 5353 2799 5411 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 8588 2836 8616 2944
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 12802 2972 12808 2984
rect 10551 2944 12808 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 8932 2907 8990 2913
rect 8932 2873 8944 2907
rect 8978 2904 8990 2907
rect 10772 2907 10830 2913
rect 8978 2876 10732 2904
rect 8978 2873 8990 2876
rect 8932 2867 8990 2873
rect 6328 2808 8616 2836
rect 6328 2796 6334 2808
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 10042 2836 10048 2848
rect 9640 2808 10048 2836
rect 9640 2796 9646 2808
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10704 2836 10732 2876
rect 10772 2873 10784 2907
rect 10818 2904 10830 2907
rect 11606 2904 11612 2916
rect 10818 2876 11612 2904
rect 10818 2873 10830 2876
rect 10772 2867 10830 2873
rect 11606 2864 11612 2876
rect 11664 2864 11670 2916
rect 13072 2907 13130 2913
rect 13072 2873 13084 2907
rect 13118 2904 13130 2907
rect 13262 2904 13268 2916
rect 13118 2876 13268 2904
rect 13118 2873 13130 2876
rect 13072 2867 13130 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 14752 2904 14780 3012
rect 15105 3009 15117 3043
rect 15151 3040 15163 3043
rect 15562 3040 15568 3052
rect 15151 3012 15568 3040
rect 15151 3009 15163 3012
rect 15105 3003 15163 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16022 3040 16028 3052
rect 15979 3012 16028 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 15657 2975 15715 2981
rect 14884 2944 14929 2972
rect 14884 2932 14890 2944
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 16298 2972 16304 2984
rect 15703 2944 16304 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 16408 2972 16436 3080
rect 18322 3068 18328 3120
rect 18380 3108 18386 3120
rect 18877 3111 18935 3117
rect 18877 3108 18889 3111
rect 18380 3080 18889 3108
rect 18380 3068 18386 3080
rect 18877 3077 18889 3080
rect 18923 3077 18935 3111
rect 18877 3071 18935 3077
rect 19429 3111 19487 3117
rect 19429 3077 19441 3111
rect 19475 3108 19487 3111
rect 20622 3108 20628 3120
rect 19475 3080 20628 3108
rect 19475 3077 19487 3080
rect 19429 3071 19487 3077
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16540 3012 17049 3040
rect 16540 3000 16546 3012
rect 17037 3009 17049 3012
rect 17083 3040 17095 3043
rect 17126 3040 17132 3052
rect 17083 3012 17132 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 18414 3000 18420 3052
rect 18472 3000 18478 3052
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 18564 3012 18613 3040
rect 18564 3000 18570 3012
rect 18601 3009 18613 3012
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 19518 3000 19524 3052
rect 19576 3040 19582 3052
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19576 3012 19901 3040
rect 19576 3000 19582 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3040 20039 3043
rect 20254 3040 20260 3052
rect 20027 3012 20260 3040
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 20254 3000 20260 3012
rect 20312 3000 20318 3052
rect 21085 3043 21143 3049
rect 21085 3009 21097 3043
rect 21131 3040 21143 3043
rect 21542 3040 21548 3052
rect 21131 3012 21548 3040
rect 21131 3009 21143 3012
rect 21085 3003 21143 3009
rect 21542 3000 21548 3012
rect 21600 3000 21606 3052
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16408 2944 16865 2972
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 17957 2975 18015 2981
rect 17957 2941 17969 2975
rect 18003 2972 18015 2975
rect 18003 2944 18184 2972
rect 18003 2941 18015 2944
rect 17957 2935 18015 2941
rect 15749 2907 15807 2913
rect 14752 2876 15332 2904
rect 11146 2836 11152 2848
rect 10704 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 14182 2836 14188 2848
rect 14143 2808 14188 2836
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 14921 2839 14979 2845
rect 14921 2805 14933 2839
rect 14967 2836 14979 2839
rect 15194 2836 15200 2848
rect 14967 2808 15200 2836
rect 14967 2805 14979 2808
rect 14921 2799 14979 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15304 2836 15332 2876
rect 15749 2873 15761 2907
rect 15795 2904 15807 2907
rect 15795 2876 18092 2904
rect 15795 2873 15807 2876
rect 15749 2867 15807 2873
rect 18064 2845 18092 2876
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 15304 2808 16957 2836
rect 16945 2805 16957 2808
rect 16991 2836 17003 2839
rect 17865 2839 17923 2845
rect 17865 2836 17877 2839
rect 16991 2808 17877 2836
rect 16991 2805 17003 2808
rect 16945 2799 17003 2805
rect 17865 2805 17877 2808
rect 17911 2805 17923 2839
rect 17865 2799 17923 2805
rect 18049 2839 18107 2845
rect 18049 2805 18061 2839
rect 18095 2805 18107 2839
rect 18156 2836 18184 2944
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 18432 2972 18460 3000
rect 19797 2975 19855 2981
rect 18432 2944 18552 2972
rect 18340 2904 18368 2932
rect 18524 2913 18552 2944
rect 19797 2941 19809 2975
rect 19843 2972 19855 2975
rect 20070 2972 20076 2984
rect 19843 2944 20076 2972
rect 19843 2941 19855 2944
rect 19797 2935 19855 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 18340 2876 18429 2904
rect 18417 2873 18429 2876
rect 18463 2873 18475 2907
rect 18417 2867 18475 2873
rect 18509 2907 18567 2913
rect 18509 2873 18521 2907
rect 18555 2873 18567 2907
rect 18509 2867 18567 2873
rect 19518 2864 19524 2916
rect 19576 2904 19582 2916
rect 19702 2904 19708 2916
rect 19576 2876 19708 2904
rect 19576 2864 19582 2876
rect 19702 2864 19708 2876
rect 19760 2864 19766 2916
rect 20809 2907 20867 2913
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 21082 2904 21088 2916
rect 20855 2876 21088 2904
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 21082 2864 21088 2876
rect 21140 2864 21146 2916
rect 19426 2836 19432 2848
rect 18156 2808 19432 2836
rect 18049 2799 18107 2805
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 20622 2836 20628 2848
rect 19852 2808 20628 2836
rect 19852 2796 19858 2808
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 20901 2839 20959 2845
rect 20901 2805 20913 2839
rect 20947 2836 20959 2839
rect 20990 2836 20996 2848
rect 20947 2808 20996 2836
rect 20947 2805 20959 2808
rect 20901 2799 20959 2805
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 5534 2632 5540 2644
rect 4847 2604 5540 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 5994 2632 6000 2644
rect 5859 2604 6000 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6270 2632 6276 2644
rect 6231 2604 6276 2632
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8202 2632 8208 2644
rect 7975 2604 8208 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11425 2635 11483 2641
rect 11425 2632 11437 2635
rect 11296 2604 11437 2632
rect 11296 2592 11302 2604
rect 11425 2601 11437 2604
rect 11471 2601 11483 2635
rect 11425 2595 11483 2601
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 12986 2632 12992 2644
rect 11931 2604 12848 2632
rect 12947 2604 12992 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 3326 2524 3332 2576
rect 3384 2564 3390 2576
rect 3384 2536 5580 2564
rect 3384 2524 3390 2536
rect 2406 2456 2412 2508
rect 2464 2496 2470 2508
rect 5169 2499 5227 2505
rect 5169 2496 5181 2499
rect 2464 2468 5181 2496
rect 2464 2456 2470 2468
rect 5169 2465 5181 2468
rect 5215 2496 5227 2499
rect 5350 2496 5356 2508
rect 5215 2468 5356 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 5552 2496 5580 2536
rect 5718 2524 5724 2576
rect 5776 2564 5782 2576
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 5776 2536 7297 2564
rect 5776 2524 5782 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 10778 2564 10784 2576
rect 10739 2536 10784 2564
rect 7285 2527 7343 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 11606 2524 11612 2576
rect 11664 2564 11670 2576
rect 12820 2564 12848 2604
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 13633 2635 13691 2641
rect 13633 2601 13645 2635
rect 13679 2601 13691 2635
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13633 2595 13691 2601
rect 13648 2564 13676 2595
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 14792 2604 15485 2632
rect 14792 2592 14798 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 16298 2592 16304 2644
rect 16356 2632 16362 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 16356 2604 16497 2632
rect 16356 2592 16362 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 18325 2635 18383 2641
rect 18325 2632 18337 2635
rect 16485 2595 16543 2601
rect 16684 2604 18337 2632
rect 11664 2536 12756 2564
rect 12820 2536 13676 2564
rect 11664 2524 11670 2536
rect 6178 2496 6184 2508
rect 5552 2468 6184 2496
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 8260 2468 8309 2496
rect 8260 2456 8266 2468
rect 8297 2465 8309 2468
rect 8343 2465 8355 2499
rect 8297 2459 8355 2465
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2465 9183 2499
rect 9858 2496 9864 2508
rect 9819 2468 9864 2496
rect 9125 2459 9183 2465
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5902 2428 5908 2440
rect 5491 2400 5908 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5902 2388 5908 2400
rect 5960 2428 5966 2440
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 5960 2400 6469 2428
rect 5960 2388 5966 2400
rect 6457 2397 6469 2400
rect 6503 2397 6515 2431
rect 6457 2391 6515 2397
rect 6472 2360 6500 2391
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7156 2400 7481 2428
rect 7156 2388 7162 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 7469 2391 7527 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9030 2428 9036 2440
rect 8619 2400 9036 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8588 2360 8616 2391
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9140 2428 9168 2459
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 12434 2496 12440 2508
rect 11839 2468 12440 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 12728 2496 12756 2536
rect 14366 2524 14372 2576
rect 14424 2564 14430 2576
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 14424 2536 14933 2564
rect 14424 2524 14430 2536
rect 14921 2533 14933 2536
rect 14967 2533 14979 2567
rect 14921 2527 14979 2533
rect 15841 2567 15899 2573
rect 15841 2533 15853 2567
rect 15887 2564 15899 2567
rect 16684 2564 16712 2604
rect 18325 2601 18337 2604
rect 18371 2601 18383 2635
rect 18690 2632 18696 2644
rect 18651 2604 18696 2632
rect 18325 2595 18383 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 18782 2592 18788 2644
rect 18840 2632 18846 2644
rect 19705 2635 19763 2641
rect 18840 2604 18885 2632
rect 18840 2592 18846 2604
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 20070 2632 20076 2644
rect 19751 2604 20076 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 15887 2536 16712 2564
rect 15887 2533 15899 2536
rect 15841 2527 15899 2533
rect 17402 2524 17408 2576
rect 17460 2564 17466 2576
rect 17773 2567 17831 2573
rect 17773 2564 17785 2567
rect 17460 2536 17785 2564
rect 17460 2524 17466 2536
rect 17773 2533 17785 2536
rect 17819 2533 17831 2567
rect 17773 2527 17831 2533
rect 17862 2524 17868 2576
rect 17920 2564 17926 2576
rect 19797 2567 19855 2573
rect 19797 2564 19809 2567
rect 17920 2536 19809 2564
rect 17920 2524 17926 2536
rect 19797 2533 19809 2536
rect 19843 2533 19855 2567
rect 19797 2527 19855 2533
rect 12728 2468 13216 2496
rect 9950 2428 9956 2440
rect 9140 2400 9956 2428
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 12066 2428 12072 2440
rect 11103 2400 12072 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13188 2437 13216 2468
rect 13998 2456 14004 2508
rect 14056 2496 14062 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 14056 2468 14105 2496
rect 14056 2456 14062 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14642 2496 14648 2508
rect 14603 2468 14648 2496
rect 14093 2459 14151 2465
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2496 15991 2499
rect 16853 2499 16911 2505
rect 16853 2496 16865 2499
rect 15979 2468 16712 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12952 2400 13093 2428
rect 12952 2388 12958 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 14182 2428 14188 2440
rect 13219 2400 14188 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 6472 2332 8616 2360
rect 9309 2363 9367 2369
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 12618 2360 12624 2372
rect 9355 2332 11192 2360
rect 12579 2332 12624 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6822 2292 6828 2304
rect 6236 2264 6828 2292
rect 6236 2252 6242 2264
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 6917 2295 6975 2301
rect 6917 2261 6929 2295
rect 6963 2292 6975 2295
rect 9674 2292 9680 2304
rect 6963 2264 9680 2292
rect 6963 2261 6975 2264
rect 6917 2255 6975 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10413 2295 10471 2301
rect 10413 2261 10425 2295
rect 10459 2292 10471 2295
rect 11054 2292 11060 2304
rect 10459 2264 11060 2292
rect 10459 2261 10471 2264
rect 10413 2255 10471 2261
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 11164 2292 11192 2332
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 16684 2360 16712 2468
rect 16776 2468 16865 2496
rect 16776 2440 16804 2468
rect 16853 2465 16865 2468
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17126 2496 17132 2508
rect 16991 2468 17132 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 17497 2499 17555 2505
rect 17497 2465 17509 2499
rect 17543 2496 17555 2499
rect 18966 2496 18972 2508
rect 17543 2468 18972 2496
rect 17543 2465 17555 2468
rect 17497 2459 17555 2465
rect 18966 2456 18972 2468
rect 19024 2456 19030 2508
rect 19242 2456 19248 2508
rect 19300 2496 19306 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 19300 2468 20545 2496
rect 19300 2456 19306 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 16758 2388 16764 2440
rect 16816 2388 16822 2440
rect 17034 2428 17040 2440
rect 16995 2400 17040 2428
rect 17034 2388 17040 2400
rect 17092 2428 17098 2440
rect 18506 2428 18512 2440
rect 17092 2400 18512 2428
rect 17092 2388 17098 2400
rect 18506 2388 18512 2400
rect 18564 2428 18570 2440
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 18564 2400 18889 2428
rect 18564 2388 18570 2400
rect 18877 2397 18889 2400
rect 18923 2428 18935 2431
rect 19889 2431 19947 2437
rect 19889 2428 19901 2431
rect 18923 2400 19901 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19889 2397 19901 2400
rect 19935 2397 19947 2431
rect 19889 2391 19947 2397
rect 19337 2363 19395 2369
rect 19337 2360 19349 2363
rect 16684 2332 19349 2360
rect 19337 2329 19349 2332
rect 19383 2329 19395 2363
rect 19337 2323 19395 2329
rect 15010 2292 15016 2304
rect 11164 2264 15016 2292
rect 15010 2252 15016 2264
rect 15068 2252 15074 2304
rect 20717 2295 20775 2301
rect 20717 2261 20729 2295
rect 20763 2292 20775 2295
rect 22278 2292 22284 2304
rect 20763 2264 22284 2292
rect 20763 2261 20775 2264
rect 20717 2255 20775 2261
rect 22278 2252 22284 2264
rect 22336 2252 22342 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 1486 2048 1492 2100
rect 1544 2088 1550 2100
rect 8202 2088 8208 2100
rect 1544 2060 8208 2088
rect 1544 2048 1550 2060
rect 8202 2048 8208 2060
rect 8260 2048 8266 2100
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 13906 2088 13912 2100
rect 9732 2060 13912 2088
rect 9732 2048 9738 2060
rect 13906 2048 13912 2060
rect 13964 2048 13970 2100
rect 8220 2020 8248 2048
rect 12158 2020 12164 2032
rect 8220 1992 12164 2020
rect 12158 1980 12164 1992
rect 12216 2020 12222 2032
rect 12894 2020 12900 2032
rect 12216 1992 12900 2020
rect 12216 1980 12222 1992
rect 12894 1980 12900 1992
rect 12952 1980 12958 2032
rect 5350 1912 5356 1964
rect 5408 1952 5414 1964
rect 12986 1952 12992 1964
rect 5408 1924 12992 1952
rect 5408 1912 5414 1924
rect 12986 1912 12992 1924
rect 13044 1912 13050 1964
rect 8386 1844 8392 1896
rect 8444 1884 8450 1896
rect 17126 1884 17132 1896
rect 8444 1856 17132 1884
rect 8444 1844 8450 1856
rect 17126 1844 17132 1856
rect 17184 1844 17190 1896
rect 198 1776 204 1828
rect 256 1816 262 1828
rect 8478 1816 8484 1828
rect 256 1788 8484 1816
rect 256 1776 262 1788
rect 8478 1776 8484 1788
rect 8536 1816 8542 1828
rect 11146 1816 11152 1828
rect 8536 1788 11152 1816
rect 8536 1776 8542 1788
rect 11146 1776 11152 1788
rect 11204 1776 11210 1828
rect 5258 1708 5264 1760
rect 5316 1748 5322 1760
rect 9766 1748 9772 1760
rect 5316 1720 9772 1748
rect 5316 1708 5322 1720
rect 9766 1708 9772 1720
rect 9824 1748 9830 1760
rect 16758 1748 16764 1760
rect 9824 1720 16764 1748
rect 9824 1708 9830 1720
rect 16758 1708 16764 1720
rect 16816 1708 16822 1760
rect 1026 1368 1032 1420
rect 1084 1408 1090 1420
rect 8386 1408 8392 1420
rect 1084 1380 8392 1408
rect 1084 1368 1090 1380
rect 8386 1368 8392 1380
rect 8444 1368 8450 1420
rect 3142 1300 3148 1352
rect 3200 1340 3206 1352
rect 5166 1340 5172 1352
rect 3200 1312 5172 1340
rect 3200 1300 3206 1312
rect 5166 1300 5172 1312
rect 5224 1300 5230 1352
rect 10042 1232 10048 1284
rect 10100 1272 10106 1284
rect 16390 1272 16396 1284
rect 10100 1244 16396 1272
rect 10100 1232 10106 1244
rect 16390 1232 16396 1244
rect 16448 1232 16454 1284
rect 13078 552 13084 604
rect 13136 592 13142 604
rect 14090 592 14096 604
rect 13136 564 14096 592
rect 13136 552 13142 564
rect 14090 552 14096 564
rect 14148 552 14154 604
rect 19334 552 19340 604
rect 19392 592 19398 604
rect 19978 592 19984 604
rect 19392 564 19984 592
rect 19392 552 19398 564
rect 19978 552 19984 564
rect 20036 552 20042 604
<< via1 >>
rect 9864 20748 9916 20800
rect 13544 20748 13596 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 2780 20544 2832 20596
rect 3700 20544 3752 20596
rect 15016 20587 15068 20596
rect 9956 20476 10008 20528
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 3332 20340 3384 20392
rect 3792 20340 3844 20392
rect 8208 20408 8260 20460
rect 9312 20408 9364 20460
rect 7380 20340 7432 20392
rect 10600 20476 10652 20528
rect 11060 20476 11112 20528
rect 10416 20408 10468 20460
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 15016 20553 15025 20587
rect 15025 20553 15059 20587
rect 15059 20553 15068 20587
rect 15016 20544 15068 20553
rect 15936 20587 15988 20596
rect 15936 20553 15945 20587
rect 15945 20553 15979 20587
rect 15979 20553 15988 20587
rect 15936 20544 15988 20553
rect 16948 20544 17000 20596
rect 20260 20544 20312 20596
rect 20628 20544 20680 20596
rect 14280 20476 14332 20528
rect 22192 20476 22244 20528
rect 2780 20272 2832 20324
rect 7196 20272 7248 20324
rect 5264 20204 5316 20256
rect 6000 20204 6052 20256
rect 6276 20247 6328 20256
rect 6276 20213 6285 20247
rect 6285 20213 6319 20247
rect 6319 20213 6328 20247
rect 6276 20204 6328 20213
rect 6920 20204 6972 20256
rect 8300 20204 8352 20256
rect 9404 20272 9456 20324
rect 10692 20340 10744 20392
rect 13360 20408 13412 20460
rect 14648 20340 14700 20392
rect 15200 20340 15252 20392
rect 16396 20340 16448 20392
rect 19524 20340 19576 20392
rect 20076 20340 20128 20392
rect 20168 20340 20220 20392
rect 13912 20315 13964 20324
rect 13912 20281 13921 20315
rect 13921 20281 13955 20315
rect 13955 20281 13964 20315
rect 13912 20272 13964 20281
rect 8852 20247 8904 20256
rect 8852 20213 8861 20247
rect 8861 20213 8895 20247
rect 8895 20213 8904 20247
rect 8852 20204 8904 20213
rect 11336 20247 11388 20256
rect 11336 20213 11345 20247
rect 11345 20213 11379 20247
rect 11379 20213 11388 20247
rect 11336 20204 11388 20213
rect 11704 20204 11756 20256
rect 12992 20247 13044 20256
rect 12992 20213 13001 20247
rect 13001 20213 13035 20247
rect 13035 20213 13044 20247
rect 12992 20204 13044 20213
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1860 20000 1912 20052
rect 3056 20043 3108 20052
rect 3056 20009 3065 20043
rect 3065 20009 3099 20043
rect 3099 20009 3108 20043
rect 3056 20000 3108 20009
rect 3792 20000 3844 20052
rect 7380 20043 7432 20052
rect 5264 19932 5316 19984
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 2780 19864 2832 19916
rect 7380 20009 7389 20043
rect 7389 20009 7423 20043
rect 7423 20009 7432 20043
rect 7380 20000 7432 20009
rect 8208 20000 8260 20052
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 11336 20000 11388 20052
rect 14740 20000 14792 20052
rect 15476 20000 15528 20052
rect 17408 20000 17460 20052
rect 17868 20000 17920 20052
rect 19800 20000 19852 20052
rect 19892 20043 19944 20052
rect 19892 20009 19901 20043
rect 19901 20009 19935 20043
rect 19935 20009 19944 20043
rect 20444 20043 20496 20052
rect 19892 20000 19944 20009
rect 20444 20009 20453 20043
rect 20453 20009 20487 20043
rect 20487 20009 20496 20043
rect 20444 20000 20496 20009
rect 21088 20043 21140 20052
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 6368 19932 6420 19984
rect 9312 19932 9364 19984
rect 10600 19975 10652 19984
rect 10600 19941 10634 19975
rect 10634 19941 10652 19975
rect 10600 19932 10652 19941
rect 10968 19932 11020 19984
rect 14188 19932 14240 19984
rect 6644 19864 6696 19916
rect 9036 19864 9088 19916
rect 3700 19796 3752 19848
rect 3792 19796 3844 19848
rect 7656 19839 7708 19848
rect 7656 19805 7665 19839
rect 7665 19805 7699 19839
rect 7699 19805 7708 19839
rect 7656 19796 7708 19805
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 2872 19660 2924 19712
rect 4068 19660 4120 19712
rect 5816 19660 5868 19712
rect 12256 19660 12308 19712
rect 12348 19660 12400 19712
rect 17040 19932 17092 19984
rect 15384 19864 15436 19916
rect 15568 19907 15620 19916
rect 15568 19873 15577 19907
rect 15577 19873 15611 19907
rect 15611 19873 15620 19907
rect 15568 19864 15620 19873
rect 16580 19864 16632 19916
rect 19156 19907 19208 19916
rect 19156 19873 19165 19907
rect 19165 19873 19199 19907
rect 19199 19873 19208 19907
rect 19156 19864 19208 19873
rect 20260 19907 20312 19916
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 20812 19864 20864 19916
rect 14464 19728 14516 19780
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 14004 19660 14056 19712
rect 20444 19796 20496 19848
rect 17960 19728 18012 19780
rect 20720 19728 20772 19780
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 6276 19456 6328 19508
rect 664 19252 716 19304
rect 2596 19252 2648 19304
rect 3516 19320 3568 19372
rect 4068 19320 4120 19372
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 2872 19184 2924 19236
rect 4528 19184 4580 19236
rect 4804 19252 4856 19304
rect 5172 19252 5224 19304
rect 6460 19388 6512 19440
rect 6828 19388 6880 19440
rect 8300 19456 8352 19508
rect 9956 19456 10008 19508
rect 11060 19456 11112 19508
rect 11980 19456 12032 19508
rect 13820 19499 13872 19508
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 20996 19499 21048 19508
rect 13820 19456 13872 19465
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 6644 19252 6696 19304
rect 11428 19388 11480 19440
rect 9312 19320 9364 19372
rect 12348 19388 12400 19440
rect 20996 19465 21005 19499
rect 21005 19465 21039 19499
rect 21039 19465 21048 19499
rect 20996 19456 21048 19465
rect 16304 19320 16356 19372
rect 6920 19184 6972 19236
rect 7564 19184 7616 19236
rect 8116 19184 8168 19236
rect 2596 19159 2648 19168
rect 2596 19125 2605 19159
rect 2605 19125 2639 19159
rect 2639 19125 2648 19159
rect 2596 19116 2648 19125
rect 3148 19116 3200 19168
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 3884 19116 3936 19168
rect 4804 19116 4856 19168
rect 5816 19116 5868 19168
rect 7748 19116 7800 19168
rect 9220 19252 9272 19304
rect 9496 19252 9548 19304
rect 10416 19252 10468 19304
rect 12532 19252 12584 19304
rect 11152 19184 11204 19236
rect 14740 19252 14792 19304
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 16120 19252 16172 19304
rect 16580 19252 16632 19304
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 8668 19116 8720 19168
rect 11244 19116 11296 19168
rect 11796 19116 11848 19168
rect 14280 19184 14332 19236
rect 16028 19184 16080 19236
rect 18236 19252 18288 19304
rect 19800 19252 19852 19304
rect 20260 19295 20312 19304
rect 20260 19261 20269 19295
rect 20269 19261 20303 19295
rect 20303 19261 20312 19295
rect 20260 19252 20312 19261
rect 12808 19116 12860 19168
rect 13452 19116 13504 19168
rect 14372 19116 14424 19168
rect 16488 19116 16540 19168
rect 18144 19116 18196 19168
rect 18880 19116 18932 19168
rect 19432 19116 19484 19168
rect 20720 19252 20772 19304
rect 21272 19184 21324 19236
rect 20536 19116 20588 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1860 18955 1912 18964
rect 1860 18921 1869 18955
rect 1869 18921 1903 18955
rect 1903 18921 1912 18955
rect 1860 18912 1912 18921
rect 1768 18844 1820 18896
rect 3240 18912 3292 18964
rect 3608 18912 3660 18964
rect 6000 18912 6052 18964
rect 7012 18912 7064 18964
rect 4620 18844 4672 18896
rect 8852 18844 8904 18896
rect 12164 18844 12216 18896
rect 1676 18819 1728 18828
rect 1676 18785 1685 18819
rect 1685 18785 1719 18819
rect 1719 18785 1728 18819
rect 1676 18776 1728 18785
rect 2044 18776 2096 18828
rect 3884 18776 3936 18828
rect 4068 18776 4120 18828
rect 5540 18776 5592 18828
rect 6828 18776 6880 18828
rect 1584 18708 1636 18760
rect 1124 18640 1176 18692
rect 3516 18640 3568 18692
rect 3700 18708 3752 18760
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 6368 18751 6420 18760
rect 6368 18717 6377 18751
rect 6377 18717 6411 18751
rect 6411 18717 6420 18751
rect 6368 18708 6420 18717
rect 8208 18776 8260 18828
rect 7380 18751 7432 18760
rect 7380 18717 7389 18751
rect 7389 18717 7423 18751
rect 7423 18717 7432 18751
rect 7380 18708 7432 18717
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 7932 18751 7984 18760
rect 7932 18717 7941 18751
rect 7941 18717 7975 18751
rect 7975 18717 7984 18751
rect 7932 18708 7984 18717
rect 9588 18776 9640 18828
rect 10876 18776 10928 18828
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 13912 18912 13964 18964
rect 14372 18955 14424 18964
rect 14372 18921 14381 18955
rect 14381 18921 14415 18955
rect 14415 18921 14424 18955
rect 14372 18912 14424 18921
rect 15384 18912 15436 18964
rect 18236 18912 18288 18964
rect 19340 18912 19392 18964
rect 21088 18955 21140 18964
rect 21088 18921 21097 18955
rect 21097 18921 21131 18955
rect 21131 18921 21140 18955
rect 21088 18912 21140 18921
rect 13820 18844 13872 18896
rect 14004 18844 14056 18896
rect 15292 18844 15344 18896
rect 18696 18844 18748 18896
rect 19432 18844 19484 18896
rect 22652 18844 22704 18896
rect 12808 18776 12860 18828
rect 14372 18776 14424 18828
rect 19708 18819 19760 18828
rect 19708 18785 19717 18819
rect 19717 18785 19751 18819
rect 19751 18785 19760 18819
rect 19708 18776 19760 18785
rect 19892 18776 19944 18828
rect 20628 18776 20680 18828
rect 9312 18708 9364 18760
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 10968 18708 11020 18760
rect 11152 18708 11204 18760
rect 11980 18708 12032 18760
rect 12256 18751 12308 18760
rect 12256 18717 12265 18751
rect 12265 18717 12299 18751
rect 12299 18717 12308 18751
rect 12256 18708 12308 18717
rect 13544 18708 13596 18760
rect 8668 18640 8720 18692
rect 8760 18640 8812 18692
rect 9864 18640 9916 18692
rect 10692 18683 10744 18692
rect 10692 18649 10701 18683
rect 10701 18649 10735 18683
rect 10735 18649 10744 18683
rect 10692 18640 10744 18649
rect 15568 18640 15620 18692
rect 4344 18572 4396 18624
rect 4988 18572 5040 18624
rect 6092 18572 6144 18624
rect 6736 18615 6788 18624
rect 6736 18581 6745 18615
rect 6745 18581 6779 18615
rect 6779 18581 6788 18615
rect 6736 18572 6788 18581
rect 7196 18572 7248 18624
rect 8208 18572 8260 18624
rect 8300 18572 8352 18624
rect 9128 18572 9180 18624
rect 11704 18572 11756 18624
rect 14096 18572 14148 18624
rect 14280 18572 14332 18624
rect 20812 18708 20864 18760
rect 21732 18640 21784 18692
rect 18144 18572 18196 18624
rect 19984 18572 20036 18624
rect 20260 18572 20312 18624
rect 20352 18572 20404 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2780 18368 2832 18420
rect 4804 18368 4856 18420
rect 5540 18411 5592 18420
rect 5540 18377 5549 18411
rect 5549 18377 5583 18411
rect 5583 18377 5592 18411
rect 5540 18368 5592 18377
rect 6828 18411 6880 18420
rect 6828 18377 6837 18411
rect 6837 18377 6871 18411
rect 6871 18377 6880 18411
rect 6828 18368 6880 18377
rect 7748 18368 7800 18420
rect 8392 18368 8444 18420
rect 2596 18232 2648 18284
rect 3700 18232 3752 18284
rect 5356 18300 5408 18352
rect 9128 18368 9180 18420
rect 10140 18368 10192 18420
rect 11060 18411 11112 18420
rect 11060 18377 11069 18411
rect 11069 18377 11103 18411
rect 11103 18377 11112 18411
rect 11060 18368 11112 18377
rect 12808 18368 12860 18420
rect 12992 18368 13044 18420
rect 14556 18368 14608 18420
rect 14832 18368 14884 18420
rect 19524 18368 19576 18420
rect 21272 18411 21324 18420
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 5632 18232 5684 18284
rect 7564 18232 7616 18284
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 2872 18096 2924 18148
rect 5172 18164 5224 18216
rect 7932 18164 7984 18216
rect 8300 18207 8352 18216
rect 8300 18173 8309 18207
rect 8309 18173 8343 18207
rect 8343 18173 8352 18207
rect 8300 18164 8352 18173
rect 11152 18300 11204 18352
rect 18144 18300 18196 18352
rect 11060 18232 11112 18284
rect 13820 18232 13872 18284
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 14188 18275 14240 18284
rect 14188 18241 14197 18275
rect 14197 18241 14231 18275
rect 14231 18241 14240 18275
rect 14188 18232 14240 18241
rect 16672 18232 16724 18284
rect 17776 18232 17828 18284
rect 18328 18232 18380 18284
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 19800 18275 19852 18284
rect 19800 18241 19809 18275
rect 19809 18241 19843 18275
rect 19843 18241 19852 18275
rect 19800 18232 19852 18241
rect 20628 18275 20680 18284
rect 20628 18241 20637 18275
rect 20637 18241 20671 18275
rect 20671 18241 20680 18275
rect 20628 18232 20680 18241
rect 4160 18139 4212 18148
rect 4160 18105 4194 18139
rect 4194 18105 4212 18139
rect 4160 18096 4212 18105
rect 4436 18096 4488 18148
rect 7472 18096 7524 18148
rect 8484 18096 8536 18148
rect 11336 18096 11388 18148
rect 11704 18096 11756 18148
rect 12624 18096 12676 18148
rect 13820 18096 13872 18148
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 5540 18028 5592 18080
rect 7012 18028 7064 18080
rect 8392 18071 8444 18080
rect 8392 18037 8401 18071
rect 8401 18037 8435 18071
rect 8435 18037 8444 18071
rect 8392 18028 8444 18037
rect 10416 18071 10468 18080
rect 10416 18037 10425 18071
rect 10425 18037 10459 18071
rect 10459 18037 10468 18071
rect 10416 18028 10468 18037
rect 10508 18071 10560 18080
rect 10508 18037 10517 18071
rect 10517 18037 10551 18071
rect 10551 18037 10560 18071
rect 10508 18028 10560 18037
rect 10692 18028 10744 18080
rect 13360 18028 13412 18080
rect 17960 18164 18012 18216
rect 18696 18164 18748 18216
rect 19340 18164 19392 18216
rect 18144 18096 18196 18148
rect 19248 18096 19300 18148
rect 16580 18028 16632 18080
rect 16764 18071 16816 18080
rect 16764 18037 16773 18071
rect 16773 18037 16807 18071
rect 16807 18037 16816 18071
rect 16764 18028 16816 18037
rect 19064 18028 19116 18080
rect 19800 18028 19852 18080
rect 20076 18028 20128 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 3240 17824 3292 17876
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 1768 17756 1820 17808
rect 4344 17824 4396 17876
rect 7380 17824 7432 17876
rect 7748 17824 7800 17876
rect 11152 17824 11204 17876
rect 11336 17867 11388 17876
rect 11336 17833 11345 17867
rect 11345 17833 11379 17867
rect 11379 17833 11388 17867
rect 11336 17824 11388 17833
rect 11888 17824 11940 17876
rect 12624 17824 12676 17876
rect 13360 17824 13412 17876
rect 13820 17867 13872 17876
rect 13820 17833 13829 17867
rect 13829 17833 13863 17867
rect 13863 17833 13872 17867
rect 13820 17824 13872 17833
rect 16764 17824 16816 17876
rect 20260 17824 20312 17876
rect 21088 17867 21140 17876
rect 21088 17833 21097 17867
rect 21097 17833 21131 17867
rect 21131 17833 21140 17867
rect 21088 17824 21140 17833
rect 22008 17867 22060 17876
rect 22008 17833 22017 17867
rect 22017 17833 22051 17867
rect 22051 17833 22060 17867
rect 22008 17824 22060 17833
rect 2136 17688 2188 17740
rect 4804 17756 4856 17808
rect 5632 17799 5684 17808
rect 5632 17765 5666 17799
rect 5666 17765 5684 17799
rect 5632 17756 5684 17765
rect 5724 17756 5776 17808
rect 10508 17756 10560 17808
rect 8668 17688 8720 17740
rect 8852 17731 8904 17740
rect 8852 17697 8861 17731
rect 8861 17697 8895 17731
rect 8895 17697 8904 17731
rect 8852 17688 8904 17697
rect 9220 17688 9272 17740
rect 9404 17688 9456 17740
rect 11060 17688 11112 17740
rect 13176 17756 13228 17808
rect 16580 17756 16632 17808
rect 19248 17756 19300 17808
rect 2228 17620 2280 17672
rect 3516 17663 3568 17672
rect 3516 17629 3525 17663
rect 3525 17629 3559 17663
rect 3559 17629 3568 17663
rect 3516 17620 3568 17629
rect 4160 17620 4212 17672
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 7472 17620 7524 17672
rect 9128 17663 9180 17672
rect 1768 17552 1820 17604
rect 3700 17552 3752 17604
rect 4436 17552 4488 17604
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 9496 17620 9548 17672
rect 10692 17620 10744 17672
rect 13636 17688 13688 17740
rect 14096 17688 14148 17740
rect 12532 17620 12584 17672
rect 6828 17484 6880 17536
rect 8300 17484 8352 17536
rect 9312 17552 9364 17604
rect 13820 17620 13872 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16304 17620 16356 17672
rect 16580 17620 16632 17672
rect 17316 17688 17368 17740
rect 17132 17620 17184 17672
rect 17224 17620 17276 17672
rect 17684 17620 17736 17672
rect 18696 17620 18748 17672
rect 19156 17620 19208 17672
rect 20076 17756 20128 17808
rect 21640 17756 21692 17808
rect 20904 17731 20956 17740
rect 20904 17697 20913 17731
rect 20913 17697 20947 17731
rect 20947 17697 20956 17731
rect 20904 17688 20956 17697
rect 18420 17552 18472 17604
rect 11060 17484 11112 17536
rect 11152 17484 11204 17536
rect 17408 17484 17460 17536
rect 18880 17484 18932 17536
rect 19340 17552 19392 17604
rect 20168 17620 20220 17672
rect 20536 17620 20588 17672
rect 21824 17552 21876 17604
rect 19616 17484 19668 17536
rect 20168 17484 20220 17536
rect 20444 17484 20496 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1492 17280 1544 17332
rect 3056 17280 3108 17332
rect 3884 17280 3936 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 5540 17280 5592 17332
rect 5724 17323 5776 17332
rect 5724 17289 5733 17323
rect 5733 17289 5767 17323
rect 5767 17289 5776 17323
rect 5724 17280 5776 17289
rect 9404 17323 9456 17332
rect 3792 17144 3844 17196
rect 5172 17144 5224 17196
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 3608 17076 3660 17128
rect 7380 17144 7432 17196
rect 7564 17187 7616 17196
rect 7564 17153 7573 17187
rect 7573 17153 7607 17187
rect 7607 17153 7616 17187
rect 7564 17144 7616 17153
rect 7656 17144 7708 17196
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 11060 17280 11112 17332
rect 12256 17280 12308 17332
rect 9220 17212 9272 17264
rect 12164 17212 12216 17264
rect 6828 17076 6880 17128
rect 3148 17008 3200 17060
rect 5172 17008 5224 17060
rect 5264 17008 5316 17060
rect 6644 17008 6696 17060
rect 6920 17008 6972 17060
rect 8576 17076 8628 17128
rect 11060 17119 11112 17128
rect 11060 17085 11069 17119
rect 11069 17085 11103 17119
rect 11103 17085 11112 17119
rect 11060 17076 11112 17085
rect 11428 17144 11480 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 11796 17144 11848 17196
rect 15476 17280 15528 17332
rect 15844 17280 15896 17332
rect 16580 17280 16632 17332
rect 18788 17280 18840 17332
rect 15660 17144 15712 17196
rect 16396 17187 16448 17196
rect 16396 17153 16405 17187
rect 16405 17153 16439 17187
rect 16439 17153 16448 17187
rect 16396 17144 16448 17153
rect 17592 17212 17644 17264
rect 19708 17280 19760 17332
rect 19156 17212 19208 17264
rect 20628 17212 20680 17264
rect 12348 17076 12400 17128
rect 13544 17076 13596 17128
rect 13820 17076 13872 17128
rect 12808 17008 12860 17060
rect 16948 17076 17000 17128
rect 18604 17076 18656 17128
rect 19156 17076 19208 17128
rect 20536 17144 20588 17196
rect 20076 17076 20128 17128
rect 14740 17008 14792 17060
rect 2964 16940 3016 16992
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 7380 16983 7432 16992
rect 4896 16940 4948 16949
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 9680 16983 9732 16992
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 11336 16940 11388 16992
rect 11888 16940 11940 16992
rect 13912 16940 13964 16992
rect 17500 17008 17552 17060
rect 18052 17008 18104 17060
rect 16580 16940 16632 16992
rect 17132 16940 17184 16992
rect 17960 16940 18012 16992
rect 18788 16983 18840 16992
rect 18788 16949 18797 16983
rect 18797 16949 18831 16983
rect 18831 16949 18840 16983
rect 18788 16940 18840 16949
rect 21916 17008 21968 17060
rect 19800 16983 19852 16992
rect 19800 16949 19809 16983
rect 19809 16949 19843 16983
rect 19843 16949 19852 16983
rect 19800 16940 19852 16949
rect 20536 16940 20588 16992
rect 20812 16983 20864 16992
rect 20812 16949 20821 16983
rect 20821 16949 20855 16983
rect 20855 16949 20864 16983
rect 20812 16940 20864 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 2504 16736 2556 16788
rect 2964 16779 3016 16788
rect 2964 16745 2973 16779
rect 2973 16745 3007 16779
rect 3007 16745 3016 16779
rect 2964 16736 3016 16745
rect 4896 16736 4948 16788
rect 6644 16779 6696 16788
rect 6644 16745 6653 16779
rect 6653 16745 6687 16779
rect 6687 16745 6696 16779
rect 6644 16736 6696 16745
rect 7380 16736 7432 16788
rect 9956 16736 10008 16788
rect 10416 16736 10468 16788
rect 204 16668 256 16720
rect 2872 16668 2924 16720
rect 3240 16668 3292 16720
rect 5172 16668 5224 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 4068 16600 4120 16652
rect 4160 16600 4212 16652
rect 5540 16600 5592 16652
rect 2596 16575 2648 16584
rect 2596 16541 2605 16575
rect 2605 16541 2639 16575
rect 2639 16541 2648 16575
rect 2596 16532 2648 16541
rect 3148 16532 3200 16584
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 4804 16532 4856 16584
rect 4988 16532 5040 16584
rect 5356 16532 5408 16584
rect 7656 16600 7708 16652
rect 8576 16668 8628 16720
rect 8668 16668 8720 16720
rect 2320 16464 2372 16516
rect 7104 16532 7156 16584
rect 9220 16532 9272 16584
rect 12440 16668 12492 16720
rect 14280 16736 14332 16788
rect 14556 16736 14608 16788
rect 15568 16736 15620 16788
rect 15844 16736 15896 16788
rect 16028 16736 16080 16788
rect 16304 16779 16356 16788
rect 16304 16745 16313 16779
rect 16313 16745 16347 16779
rect 16347 16745 16356 16779
rect 16304 16736 16356 16745
rect 16580 16736 16632 16788
rect 17316 16779 17368 16788
rect 17316 16745 17325 16779
rect 17325 16745 17359 16779
rect 17359 16745 17368 16779
rect 17316 16736 17368 16745
rect 17408 16736 17460 16788
rect 18144 16736 18196 16788
rect 20720 16736 20772 16788
rect 14004 16668 14056 16720
rect 17868 16668 17920 16720
rect 19524 16668 19576 16720
rect 19984 16668 20036 16720
rect 10968 16532 11020 16584
rect 11336 16532 11388 16584
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 1952 16439 2004 16448
rect 1952 16405 1961 16439
rect 1961 16405 1995 16439
rect 1995 16405 2004 16439
rect 1952 16396 2004 16405
rect 2872 16396 2924 16448
rect 4988 16396 5040 16448
rect 6184 16439 6236 16448
rect 6184 16405 6193 16439
rect 6193 16405 6227 16439
rect 6227 16405 6236 16439
rect 6184 16396 6236 16405
rect 7380 16464 7432 16516
rect 11704 16464 11756 16516
rect 9312 16396 9364 16448
rect 10692 16396 10744 16448
rect 13912 16600 13964 16652
rect 12072 16532 12124 16584
rect 16580 16600 16632 16652
rect 16764 16600 16816 16652
rect 17316 16600 17368 16652
rect 19248 16600 19300 16652
rect 19432 16600 19484 16652
rect 21180 16600 21232 16652
rect 12256 16464 12308 16516
rect 12992 16396 13044 16448
rect 15660 16532 15712 16584
rect 14740 16464 14792 16516
rect 17592 16532 17644 16584
rect 17960 16532 18012 16584
rect 18604 16532 18656 16584
rect 16028 16464 16080 16516
rect 19340 16464 19392 16516
rect 13360 16396 13412 16448
rect 13820 16396 13872 16448
rect 14188 16396 14240 16448
rect 15200 16396 15252 16448
rect 15660 16396 15712 16448
rect 16488 16396 16540 16448
rect 20812 16396 20864 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1492 16124 1544 16176
rect 4160 16192 4212 16244
rect 4804 16192 4856 16244
rect 6828 16192 6880 16244
rect 7656 16192 7708 16244
rect 8392 16192 8444 16244
rect 8944 16192 8996 16244
rect 11152 16192 11204 16244
rect 8576 16124 8628 16176
rect 9864 16124 9916 16176
rect 12716 16192 12768 16244
rect 13912 16192 13964 16244
rect 14096 16235 14148 16244
rect 14096 16201 14105 16235
rect 14105 16201 14139 16235
rect 14139 16201 14148 16235
rect 14096 16192 14148 16201
rect 11888 16124 11940 16176
rect 2780 15920 2832 15972
rect 2964 16056 3016 16108
rect 6368 16099 6420 16108
rect 3056 15988 3108 16040
rect 6368 16065 6377 16099
rect 6377 16065 6411 16099
rect 6411 16065 6420 16099
rect 6368 16056 6420 16065
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 9588 16056 9640 16108
rect 5724 15988 5776 16040
rect 6184 15988 6236 16040
rect 7564 15988 7616 16040
rect 3516 15920 3568 15972
rect 2504 15895 2556 15904
rect 2504 15861 2513 15895
rect 2513 15861 2547 15895
rect 2547 15861 2556 15895
rect 2504 15852 2556 15861
rect 6828 15920 6880 15972
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 6000 15852 6052 15904
rect 6276 15852 6328 15904
rect 9496 15988 9548 16040
rect 11152 16031 11204 16040
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 14740 16099 14792 16108
rect 14740 16065 14749 16099
rect 14749 16065 14783 16099
rect 14783 16065 14792 16099
rect 14740 16056 14792 16065
rect 7932 15920 7984 15972
rect 8668 15895 8720 15904
rect 8668 15861 8677 15895
rect 8677 15861 8711 15895
rect 8711 15861 8720 15895
rect 8668 15852 8720 15861
rect 9772 15895 9824 15904
rect 9772 15861 9781 15895
rect 9781 15861 9815 15895
rect 9815 15861 9824 15895
rect 9772 15852 9824 15861
rect 10416 15920 10468 15972
rect 10600 15852 10652 15904
rect 11152 15852 11204 15904
rect 11520 15988 11572 16040
rect 12348 15988 12400 16040
rect 16672 16124 16724 16176
rect 16948 16124 17000 16176
rect 19892 16124 19944 16176
rect 20260 16192 20312 16244
rect 16396 16056 16448 16108
rect 18512 16056 18564 16108
rect 19248 16056 19300 16108
rect 19708 16056 19760 16108
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 20628 16056 20680 16108
rect 15200 16031 15252 16040
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15476 16031 15528 16040
rect 15200 15988 15252 15997
rect 15476 15997 15510 16031
rect 15510 15997 15528 16031
rect 15476 15988 15528 15997
rect 16580 15988 16632 16040
rect 19340 15988 19392 16040
rect 20720 16031 20772 16040
rect 20720 15997 20729 16031
rect 20729 15997 20763 16031
rect 20763 15997 20772 16031
rect 20720 15988 20772 15997
rect 12716 15963 12768 15972
rect 12716 15929 12750 15963
rect 12750 15929 12768 15963
rect 12716 15920 12768 15929
rect 13360 15920 13412 15972
rect 18144 15920 18196 15972
rect 16488 15852 16540 15904
rect 16672 15852 16724 15904
rect 17132 15852 17184 15904
rect 17776 15852 17828 15904
rect 18052 15895 18104 15904
rect 18052 15861 18061 15895
rect 18061 15861 18095 15895
rect 18095 15861 18104 15895
rect 18052 15852 18104 15861
rect 19708 15895 19760 15904
rect 19708 15861 19717 15895
rect 19717 15861 19751 15895
rect 19751 15861 19760 15895
rect 19708 15852 19760 15861
rect 19800 15895 19852 15904
rect 19800 15861 19809 15895
rect 19809 15861 19843 15895
rect 19843 15861 19852 15895
rect 19800 15852 19852 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 3148 15648 3200 15700
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 4804 15648 4856 15700
rect 1400 15580 1452 15632
rect 2780 15580 2832 15632
rect 7564 15648 7616 15700
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 10600 15691 10652 15700
rect 9036 15623 9088 15632
rect 9036 15589 9045 15623
rect 9045 15589 9079 15623
rect 9079 15589 9088 15623
rect 9036 15580 9088 15589
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 10692 15691 10744 15700
rect 10692 15657 10701 15691
rect 10701 15657 10735 15691
rect 10735 15657 10744 15691
rect 10692 15648 10744 15657
rect 12624 15648 12676 15700
rect 16764 15648 16816 15700
rect 18052 15648 18104 15700
rect 18788 15648 18840 15700
rect 20444 15691 20496 15700
rect 14280 15623 14332 15632
rect 14280 15589 14289 15623
rect 14289 15589 14323 15623
rect 14323 15589 14332 15623
rect 14280 15580 14332 15589
rect 1492 15555 1544 15564
rect 1492 15521 1501 15555
rect 1501 15521 1535 15555
rect 1535 15521 1544 15555
rect 1492 15512 1544 15521
rect 2872 15512 2924 15564
rect 4896 15512 4948 15564
rect 5540 15512 5592 15564
rect 6920 15512 6972 15564
rect 2136 15444 2188 15496
rect 3516 15487 3568 15496
rect 3516 15453 3525 15487
rect 3525 15453 3559 15487
rect 3559 15453 3568 15487
rect 3516 15444 3568 15453
rect 3792 15444 3844 15496
rect 5448 15487 5500 15496
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 9680 15512 9732 15564
rect 10416 15512 10468 15564
rect 11336 15512 11388 15564
rect 12256 15512 12308 15564
rect 13268 15555 13320 15564
rect 13268 15521 13277 15555
rect 13277 15521 13311 15555
rect 13311 15521 13320 15555
rect 13268 15512 13320 15521
rect 16212 15580 16264 15632
rect 18512 15580 18564 15632
rect 19156 15580 19208 15632
rect 19248 15580 19300 15632
rect 2504 15308 2556 15360
rect 2964 15308 3016 15360
rect 6460 15376 6512 15428
rect 8944 15444 8996 15496
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 12624 15444 12676 15496
rect 12256 15376 12308 15428
rect 8208 15308 8260 15360
rect 9036 15308 9088 15360
rect 12716 15308 12768 15360
rect 15844 15444 15896 15496
rect 16304 15512 16356 15564
rect 18604 15555 18656 15564
rect 18604 15521 18613 15555
rect 18613 15521 18647 15555
rect 18647 15521 18656 15555
rect 18604 15512 18656 15521
rect 18696 15512 18748 15564
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 20168 15444 20220 15496
rect 14372 15376 14424 15428
rect 20812 15444 20864 15496
rect 15200 15308 15252 15360
rect 15476 15308 15528 15360
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 17776 15308 17828 15360
rect 19248 15351 19300 15360
rect 19248 15317 19257 15351
rect 19257 15317 19291 15351
rect 19291 15317 19300 15351
rect 19248 15308 19300 15317
rect 21180 15308 21232 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1860 15147 1912 15156
rect 1860 15113 1869 15147
rect 1869 15113 1903 15147
rect 1903 15113 1912 15147
rect 1860 15104 1912 15113
rect 3240 15147 3292 15156
rect 3240 15113 3249 15147
rect 3249 15113 3283 15147
rect 3283 15113 3292 15147
rect 3240 15104 3292 15113
rect 3424 15104 3476 15156
rect 3976 15104 4028 15156
rect 6276 15104 6328 15156
rect 6644 15104 6696 15156
rect 6920 15104 6972 15156
rect 7104 15104 7156 15156
rect 7840 15104 7892 15156
rect 10048 15104 10100 15156
rect 12256 15104 12308 15156
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 13360 15104 13412 15156
rect 14096 15147 14148 15156
rect 14096 15113 14105 15147
rect 14105 15113 14139 15147
rect 14139 15113 14148 15147
rect 14096 15104 14148 15113
rect 14280 15104 14332 15156
rect 15384 15104 15436 15156
rect 17960 15104 18012 15156
rect 19156 15104 19208 15156
rect 20996 15147 21048 15156
rect 20996 15113 21005 15147
rect 21005 15113 21039 15147
rect 21039 15113 21048 15147
rect 20996 15104 21048 15113
rect 3792 15011 3844 15020
rect 3792 14977 3801 15011
rect 3801 14977 3835 15011
rect 3835 14977 3844 15011
rect 3792 14968 3844 14977
rect 6828 15036 6880 15088
rect 7564 15036 7616 15088
rect 7656 15036 7708 15088
rect 10140 15079 10192 15088
rect 10140 15045 10149 15079
rect 10149 15045 10183 15079
rect 10183 15045 10192 15079
rect 10140 15036 10192 15045
rect 11520 15036 11572 15088
rect 5632 14968 5684 15020
rect 5724 15011 5776 15020
rect 5724 14977 5733 15011
rect 5733 14977 5767 15011
rect 5767 14977 5776 15011
rect 5724 14968 5776 14977
rect 6276 14968 6328 15020
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 8760 14968 8812 15020
rect 9588 14968 9640 15020
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 12440 14968 12492 15020
rect 14648 15011 14700 15020
rect 14648 14977 14657 15011
rect 14657 14977 14691 15011
rect 14691 14977 14700 15011
rect 14648 14968 14700 14977
rect 5264 14900 5316 14952
rect 6460 14943 6512 14952
rect 1768 14832 1820 14884
rect 6460 14909 6469 14943
rect 6469 14909 6503 14943
rect 6503 14909 6512 14943
rect 6460 14900 6512 14909
rect 3332 14764 3384 14816
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 5816 14832 5868 14884
rect 6000 14832 6052 14884
rect 8024 14900 8076 14952
rect 8300 14943 8352 14952
rect 8300 14909 8309 14943
rect 8309 14909 8343 14943
rect 8343 14909 8352 14943
rect 8300 14900 8352 14909
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 10416 14900 10468 14952
rect 10784 14943 10836 14952
rect 10784 14909 10818 14943
rect 10818 14909 10836 14943
rect 10784 14900 10836 14909
rect 12624 14900 12676 14952
rect 13728 14900 13780 14952
rect 15292 14943 15344 14952
rect 15292 14909 15301 14943
rect 15301 14909 15335 14943
rect 15335 14909 15344 14943
rect 15292 14900 15344 14909
rect 4068 14764 4120 14816
rect 4344 14764 4396 14816
rect 5080 14764 5132 14816
rect 5172 14764 5224 14816
rect 5448 14764 5500 14816
rect 6368 14764 6420 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 8484 14764 8536 14816
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 9496 14807 9548 14816
rect 9496 14773 9505 14807
rect 9505 14773 9539 14807
rect 9539 14773 9548 14807
rect 9496 14764 9548 14773
rect 15108 14832 15160 14884
rect 20168 15036 20220 15088
rect 17408 14968 17460 15020
rect 20352 15011 20404 15020
rect 15476 14900 15528 14952
rect 17776 14900 17828 14952
rect 20352 14977 20361 15011
rect 20361 14977 20395 15011
rect 20395 14977 20404 15011
rect 20352 14968 20404 14977
rect 16948 14832 17000 14884
rect 20260 14900 20312 14952
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 12532 14764 12584 14816
rect 13912 14764 13964 14816
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 14464 14764 14516 14773
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 14740 14764 14792 14816
rect 16304 14764 16356 14816
rect 16488 14764 16540 14816
rect 18696 14832 18748 14884
rect 17408 14764 17460 14816
rect 20168 14764 20220 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 3516 14603 3568 14612
rect 3516 14569 3525 14603
rect 3525 14569 3559 14603
rect 3559 14569 3568 14603
rect 3516 14560 3568 14569
rect 4252 14560 4304 14612
rect 3976 14492 4028 14544
rect 5724 14560 5776 14612
rect 5540 14492 5592 14544
rect 6828 14560 6880 14612
rect 8760 14560 8812 14612
rect 8852 14560 8904 14612
rect 9588 14560 9640 14612
rect 11520 14560 11572 14612
rect 12716 14560 12768 14612
rect 10048 14492 10100 14544
rect 10968 14492 11020 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 2412 14424 2464 14476
rect 3332 14288 3384 14340
rect 2044 14220 2096 14272
rect 3056 14220 3108 14272
rect 6920 14424 6972 14476
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 7104 14424 7156 14433
rect 9680 14424 9732 14476
rect 10140 14467 10192 14476
rect 10140 14433 10149 14467
rect 10149 14433 10183 14467
rect 10183 14433 10192 14467
rect 10140 14424 10192 14433
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 8944 14356 8996 14408
rect 10784 14424 10836 14476
rect 12164 14467 12216 14476
rect 12164 14433 12173 14467
rect 12173 14433 12207 14467
rect 12207 14433 12216 14467
rect 12164 14424 12216 14433
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 6552 14288 6604 14340
rect 9496 14288 9548 14340
rect 11704 14288 11756 14340
rect 4804 14220 4856 14272
rect 5448 14263 5500 14272
rect 5448 14229 5457 14263
rect 5457 14229 5491 14263
rect 5491 14229 5500 14263
rect 5448 14220 5500 14229
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 5816 14220 5868 14272
rect 8852 14220 8904 14272
rect 8944 14220 8996 14272
rect 13636 14492 13688 14544
rect 14280 14492 14332 14544
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 18604 14560 18656 14612
rect 19248 14603 19300 14612
rect 19248 14569 19257 14603
rect 19257 14569 19291 14603
rect 19291 14569 19300 14603
rect 19248 14560 19300 14569
rect 19340 14560 19392 14612
rect 20168 14560 20220 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 14832 14492 14884 14544
rect 15476 14492 15528 14544
rect 15660 14535 15712 14544
rect 15660 14501 15669 14535
rect 15669 14501 15703 14535
rect 15703 14501 15712 14535
rect 15660 14492 15712 14501
rect 15844 14492 15896 14544
rect 14372 14424 14424 14433
rect 16580 14424 16632 14476
rect 18052 14424 18104 14476
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 16304 14356 16356 14408
rect 17040 14356 17092 14408
rect 20720 14424 20772 14476
rect 18604 14356 18656 14408
rect 13912 14288 13964 14340
rect 15936 14288 15988 14340
rect 19156 14288 19208 14340
rect 20076 14356 20128 14408
rect 20352 14399 20404 14408
rect 20352 14365 20361 14399
rect 20361 14365 20395 14399
rect 20395 14365 20404 14399
rect 20352 14356 20404 14365
rect 13820 14220 13872 14272
rect 14004 14263 14056 14272
rect 14004 14229 14013 14263
rect 14013 14229 14047 14263
rect 14047 14229 14056 14263
rect 14004 14220 14056 14229
rect 14556 14220 14608 14272
rect 16764 14220 16816 14272
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 4252 14016 4304 14068
rect 5632 14016 5684 14068
rect 6460 14059 6512 14068
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 6460 14025 6469 14059
rect 6469 14025 6503 14059
rect 6503 14025 6512 14059
rect 6460 14016 6512 14025
rect 8392 14016 8444 14068
rect 13728 14016 13780 14068
rect 15200 14016 15252 14068
rect 15844 14016 15896 14068
rect 16764 14016 16816 14068
rect 18696 14016 18748 14068
rect 9404 13948 9456 14000
rect 2964 13812 3016 13864
rect 3608 13812 3660 13864
rect 4252 13812 4304 13864
rect 4988 13855 5040 13864
rect 4988 13821 5022 13855
rect 5022 13821 5040 13855
rect 3148 13744 3200 13796
rect 3700 13744 3752 13796
rect 4988 13812 5040 13821
rect 5448 13812 5500 13864
rect 7012 13812 7064 13864
rect 9588 13880 9640 13932
rect 9956 13880 10008 13932
rect 10324 13948 10376 14000
rect 12532 13948 12584 14000
rect 12716 13948 12768 14000
rect 13268 13948 13320 14000
rect 14556 13948 14608 14000
rect 16304 13948 16356 14000
rect 19708 14016 19760 14068
rect 10784 13923 10836 13932
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 10784 13880 10836 13889
rect 12624 13880 12676 13932
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 20352 13948 20404 14000
rect 20444 13880 20496 13932
rect 4804 13744 4856 13796
rect 6368 13744 6420 13796
rect 9128 13812 9180 13864
rect 12348 13812 12400 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 14740 13812 14792 13864
rect 14832 13812 14884 13864
rect 15936 13812 15988 13864
rect 20260 13812 20312 13864
rect 21180 13812 21232 13864
rect 7656 13744 7708 13796
rect 8392 13744 8444 13796
rect 9312 13744 9364 13796
rect 2136 13676 2188 13728
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 8944 13676 8996 13728
rect 9772 13744 9824 13796
rect 11428 13744 11480 13796
rect 12992 13744 13044 13796
rect 14188 13744 14240 13796
rect 14648 13744 14700 13796
rect 18604 13744 18656 13796
rect 19340 13744 19392 13796
rect 19892 13744 19944 13796
rect 20812 13744 20864 13796
rect 16488 13676 16540 13728
rect 16948 13676 17000 13728
rect 20168 13676 20220 13728
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 4344 13515 4396 13524
rect 4344 13481 4353 13515
rect 4353 13481 4387 13515
rect 4387 13481 4396 13515
rect 4344 13472 4396 13481
rect 5080 13472 5132 13524
rect 5724 13472 5776 13524
rect 6184 13472 6236 13524
rect 7104 13472 7156 13524
rect 7564 13472 7616 13524
rect 8300 13472 8352 13524
rect 8852 13515 8904 13524
rect 8852 13481 8861 13515
rect 8861 13481 8895 13515
rect 8895 13481 8904 13515
rect 8852 13472 8904 13481
rect 2044 13336 2096 13388
rect 2504 13404 2556 13456
rect 3056 13404 3108 13456
rect 5816 13404 5868 13456
rect 6460 13404 6512 13456
rect 6828 13404 6880 13456
rect 2596 13379 2648 13388
rect 2596 13345 2630 13379
rect 2630 13345 2648 13379
rect 2596 13336 2648 13345
rect 4160 13336 4212 13388
rect 7656 13404 7708 13456
rect 1400 13268 1452 13320
rect 3884 13268 3936 13320
rect 4344 13268 4396 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 4988 13311 5040 13320
rect 4988 13277 4997 13311
rect 4997 13277 5031 13311
rect 5031 13277 5040 13311
rect 4988 13268 5040 13277
rect 8852 13336 8904 13388
rect 9220 13472 9272 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 9956 13472 10008 13524
rect 10600 13472 10652 13524
rect 10784 13472 10836 13524
rect 12072 13472 12124 13524
rect 12256 13472 12308 13524
rect 6000 13268 6052 13320
rect 3700 13243 3752 13252
rect 3700 13209 3709 13243
rect 3709 13209 3743 13243
rect 3743 13209 3752 13243
rect 7380 13268 7432 13320
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 8208 13268 8260 13320
rect 10324 13404 10376 13456
rect 11428 13447 11480 13456
rect 11428 13413 11437 13447
rect 11437 13413 11471 13447
rect 11471 13413 11480 13447
rect 11428 13404 11480 13413
rect 11520 13447 11572 13456
rect 11520 13413 11529 13447
rect 11529 13413 11563 13447
rect 11563 13413 11572 13447
rect 11520 13404 11572 13413
rect 9404 13336 9456 13388
rect 9956 13336 10008 13388
rect 11152 13336 11204 13388
rect 13636 13447 13688 13456
rect 13636 13413 13670 13447
rect 13670 13413 13688 13447
rect 13636 13404 13688 13413
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 11060 13268 11112 13320
rect 11428 13268 11480 13320
rect 3700 13200 3752 13209
rect 3516 13132 3568 13184
rect 9404 13200 9456 13252
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 15660 13472 15712 13524
rect 17776 13472 17828 13524
rect 19800 13515 19852 13524
rect 16580 13404 16632 13456
rect 19800 13481 19809 13515
rect 19809 13481 19843 13515
rect 19843 13481 19852 13515
rect 19800 13472 19852 13481
rect 19708 13404 19760 13456
rect 20352 13404 20404 13456
rect 12624 13336 12676 13345
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 10140 13132 10192 13184
rect 10508 13132 10560 13184
rect 10968 13132 11020 13184
rect 16396 13336 16448 13388
rect 18052 13336 18104 13388
rect 19800 13336 19852 13388
rect 20812 13336 20864 13388
rect 14648 13268 14700 13320
rect 14832 13268 14884 13320
rect 15292 13268 15344 13320
rect 14740 13243 14792 13252
rect 14740 13209 14749 13243
rect 14749 13209 14783 13243
rect 14783 13209 14792 13243
rect 14740 13200 14792 13209
rect 15384 13200 15436 13252
rect 15660 13200 15712 13252
rect 15844 13200 15896 13252
rect 16396 13200 16448 13252
rect 17408 13268 17460 13320
rect 18696 13268 18748 13320
rect 18788 13268 18840 13320
rect 19340 13311 19392 13320
rect 19340 13277 19349 13311
rect 19349 13277 19383 13311
rect 19383 13277 19392 13311
rect 20444 13311 20496 13320
rect 19340 13268 19392 13277
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 20444 13268 20496 13277
rect 17132 13200 17184 13252
rect 17316 13200 17368 13252
rect 18144 13200 18196 13252
rect 19708 13200 19760 13252
rect 20720 13268 20772 13320
rect 18696 13132 18748 13184
rect 19524 13132 19576 13184
rect 19892 13132 19944 13184
rect 21272 13200 21324 13252
rect 20904 13132 20956 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1492 12928 1544 12980
rect 2596 12928 2648 12980
rect 4160 12971 4212 12980
rect 4160 12937 4169 12971
rect 4169 12937 4203 12971
rect 4203 12937 4212 12971
rect 4160 12928 4212 12937
rect 4804 12928 4856 12980
rect 4712 12860 4764 12912
rect 3148 12792 3200 12844
rect 3700 12792 3752 12844
rect 4068 12792 4120 12844
rect 5540 12792 5592 12844
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 2136 12724 2188 12776
rect 3792 12724 3844 12776
rect 5264 12724 5316 12776
rect 2044 12656 2096 12708
rect 8484 12928 8536 12980
rect 10048 12928 10100 12980
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 11704 12928 11756 12980
rect 9588 12860 9640 12912
rect 12072 12928 12124 12980
rect 12624 12928 12676 12980
rect 14464 12928 14516 12980
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 7380 12724 7432 12776
rect 8392 12724 8444 12776
rect 9680 12724 9732 12776
rect 3056 12588 3108 12640
rect 7840 12656 7892 12708
rect 8300 12656 8352 12708
rect 8576 12656 8628 12708
rect 9220 12656 9272 12708
rect 7564 12588 7616 12640
rect 10324 12792 10376 12844
rect 12164 12860 12216 12912
rect 9956 12588 10008 12640
rect 11888 12724 11940 12776
rect 12900 12860 12952 12912
rect 13268 12860 13320 12912
rect 14648 12860 14700 12912
rect 17040 12928 17092 12980
rect 17684 12971 17736 12980
rect 17684 12937 17693 12971
rect 17693 12937 17727 12971
rect 17727 12937 17736 12971
rect 17684 12928 17736 12937
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 14004 12792 14056 12844
rect 14740 12792 14792 12844
rect 17592 12860 17644 12912
rect 19524 12928 19576 12980
rect 19892 12928 19944 12980
rect 20076 12860 20128 12912
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 16304 12835 16356 12844
rect 16304 12801 16313 12835
rect 16313 12801 16347 12835
rect 16347 12801 16356 12835
rect 16304 12792 16356 12801
rect 17316 12792 17368 12844
rect 18512 12792 18564 12844
rect 12532 12724 12584 12776
rect 13820 12724 13872 12776
rect 14464 12724 14516 12776
rect 18880 12724 18932 12776
rect 19156 12792 19208 12844
rect 19340 12792 19392 12844
rect 20444 12860 20496 12912
rect 19524 12724 19576 12776
rect 20444 12724 20496 12776
rect 14280 12656 14332 12708
rect 17316 12656 17368 12708
rect 17776 12656 17828 12708
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 10968 12588 11020 12640
rect 11244 12588 11296 12640
rect 11980 12588 12032 12640
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12900 12631 12952 12640
rect 12440 12588 12492 12597
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 13636 12588 13688 12640
rect 15384 12588 15436 12640
rect 16764 12588 16816 12640
rect 18144 12588 18196 12640
rect 18696 12588 18748 12640
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 19248 12656 19300 12708
rect 21088 12656 21140 12708
rect 18880 12588 18932 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 3608 12427 3660 12436
rect 3608 12393 3617 12427
rect 3617 12393 3651 12427
rect 3651 12393 3660 12427
rect 3608 12384 3660 12393
rect 2228 12316 2280 12368
rect 2964 12316 3016 12368
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 8208 12427 8260 12436
rect 5080 12384 5132 12393
rect 8208 12393 8217 12427
rect 8217 12393 8251 12427
rect 8251 12393 8260 12427
rect 8208 12384 8260 12393
rect 8484 12316 8536 12368
rect 1584 12248 1636 12300
rect 2504 12248 2556 12300
rect 3148 12248 3200 12300
rect 4068 12248 4120 12300
rect 5264 12248 5316 12300
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 6368 12248 6420 12300
rect 8944 12291 8996 12300
rect 4988 12180 5040 12232
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 9128 12248 9180 12300
rect 5632 12180 5684 12189
rect 2044 12044 2096 12096
rect 3884 12112 3936 12164
rect 8576 12180 8628 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9588 12180 9640 12232
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 11152 12248 11204 12300
rect 12992 12316 13044 12368
rect 13636 12384 13688 12436
rect 17316 12384 17368 12436
rect 17868 12384 17920 12436
rect 19156 12384 19208 12436
rect 20812 12384 20864 12436
rect 14372 12316 14424 12368
rect 15292 12316 15344 12368
rect 15568 12316 15620 12368
rect 12164 12248 12216 12300
rect 12624 12248 12676 12300
rect 15200 12248 15252 12300
rect 14372 12223 14424 12232
rect 10416 12180 10468 12189
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 16304 12316 16356 12368
rect 16396 12291 16448 12300
rect 16396 12257 16430 12291
rect 16430 12257 16448 12291
rect 16396 12248 16448 12257
rect 16580 12316 16632 12368
rect 17132 12316 17184 12368
rect 17684 12316 17736 12368
rect 19248 12248 19300 12300
rect 19340 12248 19392 12300
rect 19892 12291 19944 12300
rect 19892 12257 19901 12291
rect 19901 12257 19935 12291
rect 19935 12257 19944 12291
rect 19892 12248 19944 12257
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 3424 12044 3476 12096
rect 9312 12112 9364 12164
rect 10048 12112 10100 12164
rect 13084 12112 13136 12164
rect 13360 12112 13412 12164
rect 19248 12112 19300 12164
rect 20996 12180 21048 12232
rect 10600 12044 10652 12096
rect 13452 12087 13504 12096
rect 13452 12053 13461 12087
rect 13461 12053 13495 12087
rect 13495 12053 13504 12087
rect 13452 12044 13504 12053
rect 15476 12087 15528 12096
rect 15476 12053 15485 12087
rect 15485 12053 15519 12087
rect 15519 12053 15528 12087
rect 15476 12044 15528 12053
rect 16396 12044 16448 12096
rect 17960 12044 18012 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2320 11840 2372 11892
rect 3516 11840 3568 11892
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2504 11636 2556 11688
rect 3608 11568 3660 11620
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 1952 11500 2004 11552
rect 2228 11500 2280 11552
rect 4620 11772 4672 11824
rect 5264 11815 5316 11824
rect 5264 11781 5273 11815
rect 5273 11781 5307 11815
rect 5307 11781 5316 11815
rect 5264 11772 5316 11781
rect 7656 11840 7708 11892
rect 7380 11772 7432 11824
rect 8484 11840 8536 11892
rect 8576 11840 8628 11892
rect 10508 11840 10560 11892
rect 10600 11840 10652 11892
rect 11704 11840 11756 11892
rect 5632 11704 5684 11756
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 9496 11772 9548 11824
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 10324 11772 10376 11824
rect 10968 11772 11020 11824
rect 11980 11772 12032 11824
rect 14188 11772 14240 11824
rect 12164 11704 12216 11756
rect 15476 11840 15528 11892
rect 16304 11840 16356 11892
rect 16764 11840 16816 11892
rect 19800 11840 19852 11892
rect 21456 11840 21508 11892
rect 16028 11704 16080 11756
rect 16212 11704 16264 11756
rect 16488 11747 16540 11756
rect 16488 11713 16497 11747
rect 16497 11713 16531 11747
rect 16531 11713 16540 11747
rect 16488 11704 16540 11713
rect 20444 11772 20496 11824
rect 17592 11747 17644 11756
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 18512 11704 18564 11756
rect 19248 11704 19300 11756
rect 21548 11772 21600 11824
rect 4252 11636 4304 11688
rect 4528 11636 4580 11688
rect 4804 11636 4856 11688
rect 10324 11636 10376 11688
rect 10692 11636 10744 11688
rect 10876 11636 10928 11688
rect 10968 11636 11020 11688
rect 11336 11636 11388 11688
rect 8208 11568 8260 11620
rect 8668 11568 8720 11620
rect 9036 11568 9088 11620
rect 11796 11568 11848 11620
rect 4528 11500 4580 11552
rect 5264 11500 5316 11552
rect 6828 11500 6880 11552
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 7288 11543 7340 11552
rect 7288 11509 7297 11543
rect 7297 11509 7331 11543
rect 7331 11509 7340 11543
rect 7288 11500 7340 11509
rect 9772 11500 9824 11552
rect 10784 11500 10836 11552
rect 10876 11500 10928 11552
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 11612 11500 11664 11552
rect 12348 11636 12400 11688
rect 12716 11679 12768 11688
rect 12716 11645 12750 11679
rect 12750 11645 12768 11679
rect 12716 11636 12768 11645
rect 13452 11636 13504 11688
rect 14556 11679 14608 11688
rect 14556 11645 14590 11679
rect 14590 11645 14608 11679
rect 16304 11679 16356 11688
rect 14556 11636 14608 11645
rect 16304 11645 16313 11679
rect 16313 11645 16347 11679
rect 16347 11645 16356 11679
rect 16304 11636 16356 11645
rect 16396 11679 16448 11688
rect 16396 11645 16405 11679
rect 16405 11645 16439 11679
rect 16439 11645 16448 11679
rect 16396 11636 16448 11645
rect 18052 11636 18104 11688
rect 18696 11636 18748 11688
rect 19708 11636 19760 11688
rect 12164 11568 12216 11620
rect 16672 11568 16724 11620
rect 15752 11500 15804 11552
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 18604 11568 18656 11620
rect 21088 11679 21140 11688
rect 21088 11645 21097 11679
rect 21097 11645 21131 11679
rect 21131 11645 21140 11679
rect 21088 11636 21140 11645
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 18696 11500 18748 11552
rect 19708 11500 19760 11552
rect 20444 11543 20496 11552
rect 20444 11509 20453 11543
rect 20453 11509 20487 11543
rect 20487 11509 20496 11543
rect 20444 11500 20496 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 5172 11296 5224 11348
rect 5724 11296 5776 11348
rect 7196 11296 7248 11348
rect 7380 11296 7432 11348
rect 11520 11296 11572 11348
rect 5080 11228 5132 11280
rect 8208 11228 8260 11280
rect 9588 11228 9640 11280
rect 10048 11228 10100 11280
rect 12164 11296 12216 11348
rect 12440 11296 12492 11348
rect 12808 11296 12860 11348
rect 18420 11296 18472 11348
rect 19708 11339 19760 11348
rect 11980 11228 12032 11280
rect 17776 11228 17828 11280
rect 17960 11228 18012 11280
rect 19708 11305 19717 11339
rect 19717 11305 19751 11339
rect 19751 11305 19760 11339
rect 19708 11296 19760 11305
rect 20628 11296 20680 11348
rect 21180 11271 21232 11280
rect 21180 11237 21189 11271
rect 21189 11237 21223 11271
rect 21223 11237 21232 11271
rect 21180 11228 21232 11237
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 2688 11160 2740 11212
rect 3056 11160 3108 11212
rect 5632 11160 5684 11212
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 6828 11160 6880 11212
rect 2228 11092 2280 11144
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 2780 11024 2832 11076
rect 4068 11024 4120 11076
rect 4620 11092 4672 11144
rect 5816 11092 5868 11144
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 7564 11092 7616 11144
rect 7012 11024 7064 11076
rect 7840 11067 7892 11076
rect 7840 11033 7849 11067
rect 7849 11033 7883 11067
rect 7883 11033 7892 11067
rect 7840 11024 7892 11033
rect 9680 11160 9732 11212
rect 10324 11203 10376 11212
rect 10324 11169 10333 11203
rect 10333 11169 10367 11203
rect 10367 11169 10376 11203
rect 10324 11160 10376 11169
rect 9588 11092 9640 11144
rect 10232 11092 10284 11144
rect 10508 11092 10560 11144
rect 12532 11160 12584 11212
rect 12808 11160 12860 11212
rect 14004 11160 14056 11212
rect 14188 11160 14240 11212
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 17132 11160 17184 11212
rect 19156 11160 19208 11212
rect 19340 11160 19392 11212
rect 19708 11160 19760 11212
rect 20720 11160 20772 11212
rect 12440 11092 12492 11144
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 15844 11135 15896 11144
rect 12716 11092 12768 11101
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 11796 11024 11848 11076
rect 4896 10956 4948 11008
rect 6276 10956 6328 11008
rect 7472 10956 7524 11008
rect 8576 10999 8628 11008
rect 8576 10965 8585 10999
rect 8585 10965 8619 10999
rect 8619 10965 8628 10999
rect 8576 10956 8628 10965
rect 10048 10956 10100 11008
rect 12164 10999 12216 11008
rect 12164 10965 12173 10999
rect 12173 10965 12207 10999
rect 12207 10965 12216 10999
rect 12164 10956 12216 10965
rect 14464 11024 14516 11076
rect 16672 11024 16724 11076
rect 13912 10956 13964 11008
rect 14188 10956 14240 11008
rect 16488 10956 16540 11008
rect 19248 11092 19300 11144
rect 20628 11092 20680 11144
rect 18788 10956 18840 11008
rect 19248 10999 19300 11008
rect 19248 10965 19257 10999
rect 19257 10965 19291 10999
rect 19291 10965 19300 10999
rect 19248 10956 19300 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 1768 10752 1820 10804
rect 4068 10752 4120 10804
rect 5632 10752 5684 10804
rect 6184 10752 6236 10804
rect 9220 10752 9272 10804
rect 9680 10795 9732 10804
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 11796 10752 11848 10804
rect 16488 10752 16540 10804
rect 16948 10752 17000 10804
rect 17684 10752 17736 10804
rect 2228 10616 2280 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 7472 10616 7524 10668
rect 9220 10616 9272 10668
rect 11612 10684 11664 10736
rect 12164 10684 12216 10736
rect 10140 10616 10192 10668
rect 12624 10616 12676 10668
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 14372 10616 14424 10668
rect 15384 10616 15436 10668
rect 15844 10616 15896 10668
rect 17592 10684 17644 10736
rect 2964 10548 3016 10600
rect 3516 10548 3568 10600
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 4896 10548 4948 10600
rect 4712 10480 4764 10532
rect 5540 10480 5592 10532
rect 6736 10480 6788 10532
rect 6920 10480 6972 10532
rect 7840 10548 7892 10600
rect 11244 10548 11296 10600
rect 11336 10591 11388 10600
rect 11336 10557 11345 10591
rect 11345 10557 11379 10591
rect 11379 10557 11388 10591
rect 11336 10548 11388 10557
rect 14464 10548 14516 10600
rect 15936 10548 15988 10600
rect 17500 10548 17552 10600
rect 9128 10480 9180 10532
rect 9220 10480 9272 10532
rect 9404 10480 9456 10532
rect 13176 10480 13228 10532
rect 2228 10412 2280 10464
rect 3884 10412 3936 10464
rect 5356 10412 5408 10464
rect 7012 10412 7064 10464
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 8392 10412 8444 10464
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 10232 10412 10284 10464
rect 11704 10412 11756 10464
rect 12716 10412 12768 10464
rect 13820 10412 13872 10464
rect 17224 10523 17276 10532
rect 15660 10455 15712 10464
rect 15660 10421 15669 10455
rect 15669 10421 15703 10455
rect 15703 10421 15712 10455
rect 15660 10412 15712 10421
rect 15936 10412 15988 10464
rect 17224 10489 17233 10523
rect 17233 10489 17267 10523
rect 17267 10489 17276 10523
rect 17224 10480 17276 10489
rect 17868 10480 17920 10532
rect 21364 10752 21416 10804
rect 18788 10616 18840 10668
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 19432 10480 19484 10532
rect 20076 10548 20128 10600
rect 20996 10591 21048 10600
rect 20996 10557 21005 10591
rect 21005 10557 21039 10591
rect 21039 10557 21048 10591
rect 20996 10548 21048 10557
rect 20812 10480 20864 10532
rect 17684 10412 17736 10464
rect 17776 10412 17828 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 3884 10208 3936 10260
rect 5540 10208 5592 10260
rect 6368 10208 6420 10260
rect 7104 10208 7156 10260
rect 8208 10251 8260 10260
rect 7380 10140 7432 10192
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 8576 10251 8628 10260
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 10232 10251 10284 10260
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 11152 10208 11204 10260
rect 4160 10072 4212 10124
rect 2596 9936 2648 9988
rect 3608 10004 3660 10056
rect 6368 10072 6420 10124
rect 8944 10140 8996 10192
rect 9128 10140 9180 10192
rect 11244 10140 11296 10192
rect 11796 10140 11848 10192
rect 12900 10208 12952 10260
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 9772 10072 9824 10124
rect 12164 10072 12216 10124
rect 14188 10140 14240 10192
rect 13544 10072 13596 10124
rect 15752 10140 15804 10192
rect 15384 10072 15436 10124
rect 9588 9936 9640 9988
rect 11704 9936 11756 9988
rect 12992 10004 13044 10056
rect 14372 10004 14424 10056
rect 16948 10004 17000 10056
rect 17132 10004 17184 10056
rect 17224 10004 17276 10056
rect 6000 9868 6052 9920
rect 6552 9868 6604 9920
rect 7748 9868 7800 9920
rect 11796 9868 11848 9920
rect 12624 9868 12676 9920
rect 17960 9936 18012 9988
rect 16764 9868 16816 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 18420 10208 18472 10260
rect 19248 10208 19300 10260
rect 20076 10208 20128 10260
rect 19340 10140 19392 10192
rect 21272 10140 21324 10192
rect 18788 10072 18840 10124
rect 20444 9868 20496 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 2320 9664 2372 9716
rect 2964 9664 3016 9716
rect 5356 9664 5408 9716
rect 6736 9664 6788 9716
rect 7564 9664 7616 9716
rect 3056 9460 3108 9512
rect 4068 9460 4120 9512
rect 3332 9392 3384 9444
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 7196 9596 7248 9648
rect 7288 9596 7340 9648
rect 8116 9664 8168 9716
rect 9956 9664 10008 9716
rect 8944 9639 8996 9648
rect 6920 9528 6972 9580
rect 8944 9605 8953 9639
rect 8953 9605 8987 9639
rect 8987 9605 8996 9639
rect 8944 9596 8996 9605
rect 5448 9460 5500 9512
rect 7012 9460 7064 9512
rect 7564 9460 7616 9512
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 3240 9324 3292 9376
rect 4804 9324 4856 9376
rect 5080 9324 5132 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 7472 9392 7524 9444
rect 8392 9392 8444 9444
rect 9312 9528 9364 9580
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 10692 9664 10744 9716
rect 12716 9664 12768 9716
rect 10968 9596 11020 9648
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 9956 9460 10008 9512
rect 10692 9528 10744 9580
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 13820 9596 13872 9648
rect 14464 9596 14516 9648
rect 14648 9596 14700 9648
rect 11888 9460 11940 9512
rect 12624 9460 12676 9512
rect 13176 9460 13228 9512
rect 13820 9460 13872 9512
rect 14004 9528 14056 9580
rect 14556 9460 14608 9512
rect 15752 9664 15804 9716
rect 16212 9528 16264 9580
rect 16396 9528 16448 9580
rect 16764 9528 16816 9580
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 16948 9460 17000 9512
rect 17408 9460 17460 9512
rect 18788 9664 18840 9716
rect 19984 9664 20036 9716
rect 20628 9664 20680 9716
rect 19248 9596 19300 9648
rect 19340 9596 19392 9648
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 19156 9460 19208 9512
rect 19708 9460 19760 9512
rect 20444 9460 20496 9512
rect 7380 9324 7432 9376
rect 8668 9324 8720 9376
rect 9772 9324 9824 9376
rect 10140 9324 10192 9376
rect 18788 9392 18840 9444
rect 18880 9392 18932 9444
rect 21180 9392 21232 9444
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 14740 9324 14792 9376
rect 15200 9324 15252 9376
rect 16028 9324 16080 9376
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 16488 9367 16540 9376
rect 16488 9333 16497 9367
rect 16497 9333 16531 9367
rect 16531 9333 16540 9367
rect 16488 9324 16540 9333
rect 16672 9324 16724 9376
rect 18512 9324 18564 9376
rect 19984 9324 20036 9376
rect 20720 9324 20772 9376
rect 21732 9324 21784 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 3332 9120 3384 9172
rect 3976 9120 4028 9172
rect 6644 9120 6696 9172
rect 8944 9163 8996 9172
rect 4988 9052 5040 9104
rect 6828 9052 6880 9104
rect 7012 9052 7064 9104
rect 8024 9052 8076 9104
rect 1952 8984 2004 9036
rect 5264 8984 5316 9036
rect 5356 8984 5408 9036
rect 7380 8984 7432 9036
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 3240 8916 3292 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 6552 8959 6604 8968
rect 5632 8916 5684 8925
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 6828 8916 6880 8968
rect 8944 8984 8996 9036
rect 9588 9052 9640 9104
rect 10232 9120 10284 9172
rect 11888 9120 11940 9172
rect 12900 9120 12952 9172
rect 13084 9120 13136 9172
rect 15200 9120 15252 9172
rect 16488 9120 16540 9172
rect 18144 9120 18196 9172
rect 19248 9120 19300 9172
rect 19432 9120 19484 9172
rect 21640 9120 21692 9172
rect 9680 8984 9732 9036
rect 4252 8780 4304 8832
rect 8300 8780 8352 8832
rect 8668 8848 8720 8900
rect 9404 8916 9456 8968
rect 9772 8848 9824 8900
rect 10508 8780 10560 8832
rect 11060 9052 11112 9104
rect 11520 9052 11572 9104
rect 12440 9052 12492 9104
rect 13636 9052 13688 9104
rect 10968 8984 11020 9036
rect 13084 8984 13136 9036
rect 12164 8916 12216 8968
rect 13360 8916 13412 8968
rect 11244 8891 11296 8900
rect 11244 8857 11253 8891
rect 11253 8857 11287 8891
rect 11287 8857 11296 8891
rect 11244 8848 11296 8857
rect 13728 8891 13780 8900
rect 13728 8857 13737 8891
rect 13737 8857 13771 8891
rect 13771 8857 13780 8891
rect 15292 8984 15344 9036
rect 16672 9027 16724 9036
rect 16672 8993 16681 9027
rect 16681 8993 16715 9027
rect 16715 8993 16724 9027
rect 16672 8984 16724 8993
rect 17500 8984 17552 9036
rect 18144 8984 18196 9036
rect 15200 8916 15252 8968
rect 16212 8916 16264 8968
rect 16580 8916 16632 8968
rect 13728 8848 13780 8857
rect 13820 8780 13872 8832
rect 15108 8780 15160 8832
rect 16120 8848 16172 8900
rect 16396 8848 16448 8900
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 17408 8959 17460 8968
rect 16856 8916 16908 8925
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 18512 9052 18564 9104
rect 21272 9052 21324 9104
rect 19340 8984 19392 9036
rect 19800 8984 19852 9036
rect 16948 8848 17000 8900
rect 18788 8891 18840 8900
rect 18788 8857 18797 8891
rect 18797 8857 18831 8891
rect 18831 8857 18840 8891
rect 18788 8848 18840 8857
rect 19800 8848 19852 8900
rect 15384 8780 15436 8832
rect 16212 8780 16264 8832
rect 17316 8780 17368 8832
rect 18144 8780 18196 8832
rect 18972 8780 19024 8832
rect 19524 8780 19576 8832
rect 20076 8780 20128 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 4804 8576 4856 8628
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 1952 8372 2004 8424
rect 3056 8372 3108 8424
rect 3332 8372 3384 8424
rect 5632 8440 5684 8492
rect 7196 8576 7248 8628
rect 8300 8576 8352 8628
rect 2688 8304 2740 8356
rect 3884 8347 3936 8356
rect 3884 8313 3918 8347
rect 3918 8313 3936 8347
rect 3884 8304 3936 8313
rect 4068 8236 4120 8288
rect 5540 8304 5592 8356
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 7104 8415 7156 8424
rect 7104 8381 7138 8415
rect 7138 8381 7156 8415
rect 7104 8372 7156 8381
rect 7472 8372 7524 8424
rect 9404 8576 9456 8628
rect 9588 8576 9640 8628
rect 12256 8576 12308 8628
rect 14096 8576 14148 8628
rect 16672 8576 16724 8628
rect 20628 8576 20680 8628
rect 18144 8508 18196 8560
rect 19432 8508 19484 8560
rect 11336 8440 11388 8492
rect 14004 8440 14056 8492
rect 15016 8440 15068 8492
rect 15108 8440 15160 8492
rect 16764 8440 16816 8492
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 17040 8440 17092 8492
rect 9496 8372 9548 8424
rect 10232 8372 10284 8424
rect 14096 8372 14148 8424
rect 8484 8304 8536 8356
rect 8944 8304 8996 8356
rect 10600 8304 10652 8356
rect 11704 8304 11756 8356
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 14372 8304 14424 8356
rect 14648 8304 14700 8356
rect 11152 8236 11204 8288
rect 11244 8236 11296 8288
rect 13912 8236 13964 8288
rect 14096 8279 14148 8288
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 14096 8236 14148 8245
rect 15292 8372 15344 8424
rect 15660 8415 15712 8424
rect 15660 8381 15669 8415
rect 15669 8381 15703 8415
rect 15703 8381 15712 8415
rect 15660 8372 15712 8381
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 19064 8440 19116 8492
rect 20996 8508 21048 8560
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 15108 8304 15160 8356
rect 16764 8347 16816 8356
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 17684 8304 17736 8356
rect 18788 8304 18840 8356
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 17592 8236 17644 8288
rect 17776 8236 17828 8288
rect 18328 8236 18380 8288
rect 19340 8236 19392 8288
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 20352 8236 20404 8288
rect 21456 8236 21508 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 2412 8032 2464 8084
rect 5540 8032 5592 8084
rect 5632 8032 5684 8084
rect 1676 7964 1728 8016
rect 2596 8007 2648 8016
rect 2596 7973 2605 8007
rect 2605 7973 2639 8007
rect 2639 7973 2648 8007
rect 2596 7964 2648 7973
rect 6000 7964 6052 8016
rect 6368 7964 6420 8016
rect 7380 7964 7432 8016
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 8668 8032 8720 8084
rect 13176 8032 13228 8084
rect 14096 8032 14148 8084
rect 15660 8032 15712 8084
rect 16212 8032 16264 8084
rect 16672 8032 16724 8084
rect 17040 8032 17092 8084
rect 17408 8075 17460 8084
rect 17408 8041 17417 8075
rect 17417 8041 17451 8075
rect 17451 8041 17460 8075
rect 17408 8032 17460 8041
rect 18328 8032 18380 8084
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 5816 7896 5868 7948
rect 6920 7896 6972 7948
rect 8208 7896 8260 7948
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 3884 7828 3936 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 8024 7828 8076 7880
rect 9588 7828 9640 7880
rect 9772 7964 9824 8016
rect 14740 7964 14792 8016
rect 13728 7896 13780 7948
rect 14372 7939 14424 7948
rect 14372 7905 14381 7939
rect 14381 7905 14415 7939
rect 14415 7905 14424 7939
rect 14372 7896 14424 7905
rect 14648 7896 14700 7948
rect 15752 7964 15804 8016
rect 18880 7964 18932 8016
rect 19984 7964 20036 8016
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15384 7896 15436 7948
rect 19156 7896 19208 7948
rect 9772 7828 9824 7880
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 10876 7828 10928 7880
rect 11796 7828 11848 7880
rect 3976 7760 4028 7812
rect 7196 7760 7248 7812
rect 6184 7692 6236 7744
rect 7564 7692 7616 7744
rect 17500 7871 17552 7880
rect 17500 7837 17509 7871
rect 17509 7837 17543 7871
rect 17543 7837 17552 7871
rect 17500 7828 17552 7837
rect 17684 7828 17736 7880
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 10876 7692 10928 7744
rect 11244 7692 11296 7744
rect 12164 7692 12216 7744
rect 12716 7692 12768 7744
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14556 7735 14608 7744
rect 14096 7692 14148 7701
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 16856 7692 16908 7744
rect 17592 7692 17644 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 20628 7692 20680 7744
rect 21548 7692 21600 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 2504 7488 2556 7540
rect 4068 7488 4120 7540
rect 2688 7420 2740 7472
rect 3516 7420 3568 7472
rect 3700 7420 3752 7472
rect 5816 7488 5868 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 8024 7488 8076 7540
rect 8576 7488 8628 7540
rect 9128 7488 9180 7540
rect 2596 7352 2648 7404
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 3056 7284 3108 7336
rect 3424 7284 3476 7336
rect 10692 7420 10744 7472
rect 12256 7488 12308 7540
rect 13452 7420 13504 7472
rect 16856 7420 16908 7472
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 7748 7352 7800 7404
rect 8944 7352 8996 7404
rect 3148 7216 3200 7268
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 3700 7148 3752 7200
rect 4160 7148 4212 7200
rect 6644 7148 6696 7200
rect 6920 7216 6972 7268
rect 9128 7284 9180 7336
rect 9496 7352 9548 7404
rect 14464 7352 14516 7404
rect 9588 7284 9640 7336
rect 9680 7284 9732 7336
rect 10508 7284 10560 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 12716 7284 12768 7336
rect 15200 7284 15252 7336
rect 15568 7284 15620 7336
rect 16304 7352 16356 7404
rect 16488 7395 16540 7404
rect 16488 7361 16497 7395
rect 16497 7361 16531 7395
rect 16531 7361 16540 7395
rect 17592 7395 17644 7404
rect 16488 7352 16540 7361
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 18880 7488 18932 7540
rect 20260 7488 20312 7540
rect 16212 7284 16264 7336
rect 17316 7327 17368 7336
rect 7564 7216 7616 7268
rect 7472 7148 7524 7200
rect 8300 7148 8352 7200
rect 8668 7191 8720 7200
rect 8668 7157 8677 7191
rect 8677 7157 8711 7191
rect 8711 7157 8720 7191
rect 8668 7148 8720 7157
rect 8852 7216 8904 7268
rect 10416 7216 10468 7268
rect 10600 7216 10652 7268
rect 14004 7216 14056 7268
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 18512 7284 18564 7336
rect 19800 7352 19852 7404
rect 20260 7352 20312 7404
rect 9404 7148 9456 7200
rect 10048 7148 10100 7200
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 11796 7148 11848 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 12624 7148 12676 7200
rect 14464 7148 14516 7200
rect 14740 7148 14792 7200
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 19892 7216 19944 7268
rect 18052 7148 18104 7200
rect 19064 7148 19116 7200
rect 21824 7284 21876 7336
rect 21916 7216 21968 7268
rect 21088 7148 21140 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 3240 6944 3292 6996
rect 3884 6944 3936 6996
rect 4160 6944 4212 6996
rect 5264 6944 5316 6996
rect 5724 6944 5776 6996
rect 6184 6987 6236 6996
rect 6184 6953 6193 6987
rect 6193 6953 6227 6987
rect 6227 6953 6236 6987
rect 6184 6944 6236 6953
rect 7564 6944 7616 6996
rect 8668 6944 8720 6996
rect 8944 6944 8996 6996
rect 9128 6944 9180 6996
rect 10416 6944 10468 6996
rect 4344 6876 4396 6928
rect 6092 6919 6144 6928
rect 6092 6885 6101 6919
rect 6101 6885 6135 6919
rect 6135 6885 6144 6919
rect 6092 6876 6144 6885
rect 6552 6876 6604 6928
rect 6644 6876 6696 6928
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 2780 6808 2832 6860
rect 3240 6808 3292 6860
rect 4068 6740 4120 6792
rect 6000 6808 6052 6860
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6644 6740 6696 6792
rect 6828 6740 6880 6792
rect 1860 6604 1912 6656
rect 3516 6604 3568 6656
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 6092 6672 6144 6724
rect 7288 6672 7340 6724
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 9128 6783 9180 6792
rect 8944 6740 8996 6749
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9588 6740 9640 6792
rect 9496 6672 9548 6724
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 11796 6808 11848 6860
rect 12532 6808 12584 6860
rect 13728 6944 13780 6996
rect 15844 6944 15896 6996
rect 15936 6944 15988 6996
rect 18604 6944 18656 6996
rect 10048 6740 10100 6792
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 15752 6876 15804 6928
rect 13912 6740 13964 6792
rect 15384 6740 15436 6792
rect 16120 6876 16172 6928
rect 16488 6919 16540 6928
rect 16488 6885 16497 6919
rect 16497 6885 16531 6919
rect 16531 6885 16540 6919
rect 16488 6876 16540 6885
rect 16672 6876 16724 6928
rect 18880 6876 18932 6928
rect 17408 6808 17460 6860
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 18788 6851 18840 6860
rect 18788 6817 18822 6851
rect 18822 6817 18840 6851
rect 18788 6808 18840 6817
rect 16304 6740 16356 6792
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 20720 6740 20772 6792
rect 11888 6672 11940 6724
rect 11704 6604 11756 6656
rect 17224 6672 17276 6724
rect 19892 6715 19944 6724
rect 19892 6681 19901 6715
rect 19901 6681 19935 6715
rect 19935 6681 19944 6715
rect 19892 6672 19944 6681
rect 15384 6604 15436 6656
rect 15660 6604 15712 6656
rect 17776 6604 17828 6656
rect 18052 6604 18104 6656
rect 18696 6604 18748 6656
rect 20904 6604 20956 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 3056 6443 3108 6452
rect 2780 6400 2832 6409
rect 3056 6409 3065 6443
rect 3065 6409 3099 6443
rect 3099 6409 3108 6443
rect 3056 6400 3108 6409
rect 4252 6400 4304 6452
rect 5816 6400 5868 6452
rect 6552 6400 6604 6452
rect 8208 6400 8260 6452
rect 8300 6400 8352 6452
rect 9680 6400 9732 6452
rect 10416 6400 10468 6452
rect 15476 6400 15528 6452
rect 16488 6400 16540 6452
rect 16580 6400 16632 6452
rect 17684 6400 17736 6452
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 1952 6196 2004 6248
rect 3332 6196 3384 6248
rect 4712 6196 4764 6248
rect 4804 6196 4856 6248
rect 5816 6264 5868 6316
rect 6276 6264 6328 6316
rect 6828 6264 6880 6316
rect 9496 6332 9548 6384
rect 10692 6332 10744 6384
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 15200 6332 15252 6384
rect 17592 6332 17644 6384
rect 20168 6400 20220 6452
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 16120 6264 16172 6316
rect 2320 6128 2372 6180
rect 3884 6128 3936 6180
rect 4252 6128 4304 6180
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 3976 6060 4028 6112
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 6644 6060 6696 6112
rect 7196 6060 7248 6112
rect 7748 6060 7800 6112
rect 10048 6196 10100 6248
rect 11244 6196 11296 6248
rect 12440 6196 12492 6248
rect 12716 6196 12768 6248
rect 14740 6196 14792 6248
rect 15568 6196 15620 6248
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 16580 6307 16632 6316
rect 16580 6273 16589 6307
rect 16589 6273 16623 6307
rect 16623 6273 16632 6307
rect 16580 6264 16632 6273
rect 18788 6264 18840 6316
rect 19340 6264 19392 6316
rect 20996 6332 21048 6384
rect 19892 6264 19944 6316
rect 20260 6264 20312 6316
rect 17224 6196 17276 6248
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 19616 6196 19668 6248
rect 20536 6239 20588 6248
rect 20536 6205 20545 6239
rect 20545 6205 20579 6239
rect 20579 6205 20588 6239
rect 20536 6196 20588 6205
rect 21180 6196 21232 6248
rect 8208 6171 8260 6180
rect 8208 6137 8242 6171
rect 8242 6137 8260 6171
rect 8208 6128 8260 6137
rect 8300 6128 8352 6180
rect 8392 6060 8444 6112
rect 8944 6128 8996 6180
rect 9588 6060 9640 6112
rect 9680 6060 9732 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 10784 6060 10836 6112
rect 11244 6060 11296 6112
rect 11796 6060 11848 6112
rect 12164 6060 12216 6112
rect 15568 6060 15620 6112
rect 16028 6060 16080 6112
rect 18604 6128 18656 6180
rect 18788 6128 18840 6180
rect 18236 6060 18288 6112
rect 18696 6060 18748 6112
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2320 5856 2372 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 4068 5899 4120 5908
rect 4068 5865 4077 5899
rect 4077 5865 4111 5899
rect 4111 5865 4120 5899
rect 4068 5856 4120 5865
rect 5540 5856 5592 5908
rect 6092 5856 6144 5908
rect 6368 5856 6420 5908
rect 6736 5856 6788 5908
rect 7104 5856 7156 5908
rect 10048 5856 10100 5908
rect 10416 5856 10468 5908
rect 11152 5856 11204 5908
rect 5724 5788 5776 5840
rect 8300 5788 8352 5840
rect 1952 5720 2004 5772
rect 2596 5720 2648 5772
rect 6000 5720 6052 5772
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 8668 5720 8720 5772
rect 9312 5720 9364 5772
rect 4252 5652 4304 5704
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6828 5584 6880 5636
rect 8300 5652 8352 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 8392 5584 8444 5636
rect 9496 5720 9548 5772
rect 11612 5788 11664 5840
rect 13820 5788 13872 5840
rect 14280 5788 14332 5840
rect 15660 5831 15712 5840
rect 15660 5797 15694 5831
rect 15694 5797 15712 5831
rect 15660 5788 15712 5797
rect 16396 5856 16448 5908
rect 18236 5856 18288 5908
rect 17500 5788 17552 5840
rect 18880 5788 18932 5840
rect 19340 5856 19392 5908
rect 19708 5856 19760 5908
rect 19616 5788 19668 5840
rect 11796 5720 11848 5772
rect 12440 5720 12492 5772
rect 13084 5763 13136 5772
rect 13084 5729 13093 5763
rect 13093 5729 13127 5763
rect 13127 5729 13136 5763
rect 13084 5720 13136 5729
rect 13176 5695 13228 5704
rect 12072 5584 12124 5636
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 6092 5559 6144 5568
rect 6092 5525 6101 5559
rect 6101 5525 6135 5559
rect 6135 5525 6144 5559
rect 6092 5516 6144 5525
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 7748 5516 7800 5568
rect 7932 5516 7984 5568
rect 9588 5516 9640 5568
rect 10324 5516 10376 5568
rect 11796 5516 11848 5568
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 14004 5720 14056 5772
rect 14648 5720 14700 5772
rect 14924 5720 14976 5772
rect 15476 5720 15528 5772
rect 18512 5763 18564 5772
rect 18512 5729 18521 5763
rect 18521 5729 18555 5763
rect 18555 5729 18564 5763
rect 18512 5720 18564 5729
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 17500 5695 17552 5704
rect 14648 5584 14700 5636
rect 12440 5516 12492 5568
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 17868 5652 17920 5704
rect 21088 5720 21140 5772
rect 21180 5652 21232 5704
rect 21364 5584 21416 5636
rect 15660 5516 15712 5568
rect 15752 5516 15804 5568
rect 16396 5516 16448 5568
rect 16488 5516 16540 5568
rect 20996 5516 21048 5568
rect 21824 5516 21876 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 3424 5312 3476 5364
rect 7472 5312 7524 5364
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 8300 5312 8352 5364
rect 9036 5312 9088 5364
rect 9312 5312 9364 5364
rect 2320 5176 2372 5228
rect 3240 5108 3292 5160
rect 4160 5108 4212 5160
rect 5816 5108 5868 5160
rect 6092 5151 6144 5160
rect 6092 5117 6101 5151
rect 6101 5117 6135 5151
rect 6135 5117 6144 5151
rect 6092 5108 6144 5117
rect 6644 5108 6696 5160
rect 8300 5176 8352 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 9588 5176 9640 5228
rect 10324 5176 10376 5228
rect 11796 5244 11848 5296
rect 15936 5312 15988 5364
rect 16304 5312 16356 5364
rect 17224 5312 17276 5364
rect 17500 5312 17552 5364
rect 19432 5312 19484 5364
rect 20168 5355 20220 5364
rect 20168 5321 20177 5355
rect 20177 5321 20211 5355
rect 20211 5321 20220 5355
rect 20168 5312 20220 5321
rect 13084 5244 13136 5296
rect 14832 5244 14884 5296
rect 15476 5244 15528 5296
rect 20444 5244 20496 5296
rect 12072 5176 12124 5228
rect 13544 5176 13596 5228
rect 13636 5176 13688 5228
rect 15200 5176 15252 5228
rect 2136 5040 2188 5092
rect 3148 5040 3200 5092
rect 3608 5040 3660 5092
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 2596 4972 2648 5024
rect 4252 4972 4304 5024
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 9496 5108 9548 5160
rect 10140 5108 10192 5160
rect 11060 5108 11112 5160
rect 11796 5151 11848 5160
rect 11796 5117 11805 5151
rect 11805 5117 11839 5151
rect 11839 5117 11848 5151
rect 11796 5108 11848 5117
rect 7104 5083 7156 5092
rect 7104 5049 7138 5083
rect 7138 5049 7156 5083
rect 7104 5040 7156 5049
rect 7196 5040 7248 5092
rect 7472 4972 7524 5024
rect 7748 5040 7800 5092
rect 9312 5040 9364 5092
rect 13360 5040 13412 5092
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 9128 4972 9180 5024
rect 10416 4972 10468 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 11336 4972 11388 5024
rect 12624 4972 12676 5024
rect 13084 4972 13136 5024
rect 14740 5108 14792 5160
rect 15292 5040 15344 5092
rect 19708 5219 19760 5228
rect 15660 5151 15712 5160
rect 15660 5117 15669 5151
rect 15669 5117 15703 5151
rect 15703 5117 15712 5151
rect 15660 5108 15712 5117
rect 16488 5108 16540 5160
rect 16672 5108 16724 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 19708 5185 19717 5219
rect 19717 5185 19751 5219
rect 19751 5185 19760 5219
rect 19708 5176 19760 5185
rect 20996 5219 21048 5228
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 19340 5108 19392 5160
rect 20168 5108 20220 5160
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 16028 5040 16080 5092
rect 17960 5040 18012 5092
rect 13820 4972 13872 5024
rect 14188 4972 14240 5024
rect 15476 4972 15528 5024
rect 16488 4972 16540 5024
rect 18420 4972 18472 5024
rect 19616 5015 19668 5024
rect 19616 4981 19625 5015
rect 19625 4981 19659 5015
rect 19659 4981 19668 5015
rect 19616 4972 19668 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 5172 4768 5224 4820
rect 7288 4768 7340 4820
rect 9036 4768 9088 4820
rect 9956 4768 10008 4820
rect 10692 4768 10744 4820
rect 13452 4768 13504 4820
rect 15568 4768 15620 4820
rect 15660 4768 15712 4820
rect 1768 4496 1820 4548
rect 9128 4700 9180 4752
rect 10048 4743 10100 4752
rect 10048 4709 10057 4743
rect 10057 4709 10091 4743
rect 10091 4709 10100 4743
rect 10048 4700 10100 4709
rect 10968 4700 11020 4752
rect 5632 4632 5684 4684
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 11060 4675 11112 4684
rect 11060 4641 11069 4675
rect 11069 4641 11103 4675
rect 11103 4641 11112 4675
rect 11060 4632 11112 4641
rect 11336 4632 11388 4684
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 4252 4564 4304 4616
rect 5172 4564 5224 4616
rect 5356 4564 5408 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 7748 4607 7800 4616
rect 2964 4496 3016 4548
rect 4068 4428 4120 4480
rect 7104 4496 7156 4548
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 8484 4564 8536 4616
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 8852 4607 8904 4616
rect 8852 4573 8861 4607
rect 8861 4573 8895 4607
rect 8895 4573 8904 4607
rect 8852 4564 8904 4573
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 11152 4564 11204 4616
rect 9588 4496 9640 4548
rect 9956 4496 10008 4548
rect 12532 4564 12584 4616
rect 13912 4632 13964 4684
rect 15752 4632 15804 4684
rect 17868 4768 17920 4820
rect 19616 4768 19668 4820
rect 16304 4700 16356 4752
rect 18420 4700 18472 4752
rect 15200 4564 15252 4616
rect 19340 4632 19392 4684
rect 19800 4675 19852 4684
rect 19800 4641 19809 4675
rect 19809 4641 19843 4675
rect 19843 4641 19852 4675
rect 19800 4632 19852 4641
rect 21272 4632 21324 4684
rect 20996 4564 21048 4616
rect 14096 4496 14148 4548
rect 15568 4496 15620 4548
rect 17224 4539 17276 4548
rect 17224 4505 17233 4539
rect 17233 4505 17267 4539
rect 17267 4505 17276 4539
rect 17224 4496 17276 4505
rect 18880 4539 18932 4548
rect 18880 4505 18889 4539
rect 18889 4505 18923 4539
rect 18923 4505 18932 4539
rect 18880 4496 18932 4505
rect 7196 4471 7248 4480
rect 7196 4437 7205 4471
rect 7205 4437 7239 4471
rect 7239 4437 7248 4471
rect 7196 4428 7248 4437
rect 7656 4428 7708 4480
rect 8300 4428 8352 4480
rect 13544 4428 13596 4480
rect 13636 4428 13688 4480
rect 14188 4428 14240 4480
rect 14832 4428 14884 4480
rect 19340 4428 19392 4480
rect 22744 4428 22796 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2412 4267 2464 4276
rect 2412 4233 2421 4267
rect 2421 4233 2455 4267
rect 2455 4233 2464 4267
rect 2412 4224 2464 4233
rect 2688 4156 2740 4208
rect 3792 4088 3844 4140
rect 4160 4088 4212 4140
rect 2872 4020 2924 4072
rect 3240 4020 3292 4072
rect 4988 4063 5040 4072
rect 4988 4029 4997 4063
rect 4997 4029 5031 4063
rect 5031 4029 5040 4063
rect 4988 4020 5040 4029
rect 7748 4224 7800 4276
rect 8852 4224 8904 4276
rect 8944 4224 8996 4276
rect 9588 4224 9640 4276
rect 13452 4224 13504 4276
rect 6736 4156 6788 4208
rect 7196 4088 7248 4140
rect 9036 4156 9088 4208
rect 9312 4156 9364 4208
rect 4160 3952 4212 4004
rect 5448 3952 5500 4004
rect 8852 4088 8904 4140
rect 9864 4088 9916 4140
rect 10508 4156 10560 4208
rect 13728 4224 13780 4276
rect 14188 4224 14240 4276
rect 14648 4224 14700 4276
rect 15108 4224 15160 4276
rect 11152 4131 11204 4140
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 11888 4088 11940 4140
rect 13636 4156 13688 4208
rect 14096 4088 14148 4140
rect 14740 4156 14792 4208
rect 15844 4224 15896 4276
rect 19892 4224 19944 4276
rect 15568 4156 15620 4208
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 16396 4156 16448 4208
rect 17868 4156 17920 4208
rect 20260 4156 20312 4208
rect 16948 4088 17000 4140
rect 17132 4088 17184 4140
rect 17224 4088 17276 4140
rect 17592 4088 17644 4140
rect 18880 4088 18932 4140
rect 20168 4088 20220 4140
rect 20812 4088 20864 4140
rect 3608 3884 3660 3936
rect 5632 3884 5684 3936
rect 6736 3884 6788 3936
rect 7380 3952 7432 4004
rect 7472 3952 7524 4004
rect 9312 3952 9364 4004
rect 9772 4020 9824 4072
rect 10876 4020 10928 4072
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 13176 4020 13228 4072
rect 11888 3952 11940 4004
rect 17316 4020 17368 4072
rect 18052 4020 18104 4072
rect 14924 3995 14976 4004
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 10876 3927 10928 3936
rect 10876 3893 10885 3927
rect 10885 3893 10919 3927
rect 10919 3893 10928 3927
rect 10876 3884 10928 3893
rect 11244 3884 11296 3936
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 14924 3961 14933 3995
rect 14933 3961 14967 3995
rect 14967 3961 14976 3995
rect 14924 3952 14976 3961
rect 15016 3995 15068 4004
rect 15016 3961 15025 3995
rect 15025 3961 15059 3995
rect 15059 3961 15068 3995
rect 15016 3952 15068 3961
rect 15200 3952 15252 4004
rect 20996 3952 21048 4004
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 18236 3884 18288 3936
rect 18604 3884 18656 3936
rect 19800 3884 19852 3936
rect 19984 3884 20036 3936
rect 20812 3927 20864 3936
rect 20812 3893 20821 3927
rect 20821 3893 20855 3927
rect 20855 3893 20864 3927
rect 20812 3884 20864 3893
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 5724 3680 5776 3732
rect 3240 3544 3292 3596
rect 3608 3544 3660 3596
rect 4988 3544 5040 3596
rect 5540 3544 5592 3596
rect 6092 3680 6144 3732
rect 6828 3680 6880 3732
rect 6184 3612 6236 3664
rect 10508 3612 10560 3664
rect 10876 3680 10928 3732
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 13176 3680 13228 3732
rect 13268 3680 13320 3732
rect 13728 3680 13780 3732
rect 14280 3680 14332 3732
rect 15292 3723 15344 3732
rect 12716 3612 12768 3664
rect 15292 3689 15301 3723
rect 15301 3689 15335 3723
rect 15335 3689 15344 3723
rect 15292 3680 15344 3689
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 16580 3680 16632 3732
rect 17040 3723 17092 3732
rect 7288 3544 7340 3596
rect 9864 3544 9916 3596
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 2964 3476 3016 3528
rect 3976 3476 4028 3528
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 5632 3476 5684 3528
rect 7472 3476 7524 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 12624 3544 12676 3596
rect 13636 3544 13688 3596
rect 16764 3612 16816 3664
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 16672 3544 16724 3596
rect 17500 3612 17552 3664
rect 18696 3680 18748 3732
rect 21180 3655 21232 3664
rect 21180 3621 21189 3655
rect 21189 3621 21223 3655
rect 21223 3621 21232 3655
rect 21180 3612 21232 3621
rect 17684 3544 17736 3596
rect 18880 3544 18932 3596
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 12532 3476 12584 3528
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 13820 3476 13872 3528
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 16028 3476 16080 3528
rect 17500 3476 17552 3528
rect 20352 3544 20404 3596
rect 21088 3544 21140 3596
rect 20168 3519 20220 3528
rect 1952 3451 2004 3460
rect 1952 3417 1961 3451
rect 1961 3417 1995 3451
rect 1995 3417 2004 3451
rect 1952 3408 2004 3417
rect 9312 3451 9364 3460
rect 3056 3340 3108 3392
rect 5724 3340 5776 3392
rect 7288 3340 7340 3392
rect 7748 3340 7800 3392
rect 9312 3417 9321 3451
rect 9321 3417 9355 3451
rect 9355 3417 9364 3451
rect 9312 3408 9364 3417
rect 15200 3408 15252 3460
rect 16212 3408 16264 3460
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 8300 3340 8352 3392
rect 11152 3383 11204 3392
rect 11152 3349 11161 3383
rect 11161 3349 11195 3383
rect 11195 3349 11204 3383
rect 11152 3340 11204 3349
rect 11704 3340 11756 3392
rect 13176 3340 13228 3392
rect 13544 3340 13596 3392
rect 17224 3340 17276 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3056 3136 3108 3188
rect 5264 3136 5316 3188
rect 6920 3136 6972 3188
rect 7196 3179 7248 3188
rect 7196 3145 7205 3179
rect 7205 3145 7239 3179
rect 7239 3145 7248 3179
rect 7196 3136 7248 3145
rect 7932 3136 7984 3188
rect 3700 3000 3752 3052
rect 7288 3068 7340 3120
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 4988 2932 5040 2984
rect 8576 3000 8628 3052
rect 9772 3136 9824 3188
rect 9864 3136 9916 3188
rect 12072 3136 12124 3188
rect 14096 3136 14148 3188
rect 15752 3136 15804 3188
rect 17132 3136 17184 3188
rect 18696 3136 18748 3188
rect 20812 3136 20864 3188
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 16304 3111 16356 3120
rect 16304 3077 16313 3111
rect 16313 3077 16347 3111
rect 16347 3077 16356 3111
rect 16304 3068 16356 3077
rect 1952 2864 2004 2916
rect 3240 2796 3292 2848
rect 3516 2796 3568 2848
rect 4252 2907 4304 2916
rect 4252 2873 4286 2907
rect 4286 2873 4304 2907
rect 4252 2864 4304 2873
rect 5264 2796 5316 2848
rect 5540 2864 5592 2916
rect 8208 2864 8260 2916
rect 6000 2839 6052 2848
rect 6000 2805 6009 2839
rect 6009 2805 6043 2839
rect 6043 2805 6052 2839
rect 6000 2796 6052 2805
rect 6276 2796 6328 2848
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 9588 2796 9640 2848
rect 10048 2796 10100 2848
rect 11612 2864 11664 2916
rect 13268 2864 13320 2916
rect 15568 3000 15620 3052
rect 16028 3000 16080 3052
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 16304 2932 16356 2984
rect 18328 3068 18380 3120
rect 20628 3068 20680 3120
rect 16488 3000 16540 3052
rect 17132 3000 17184 3052
rect 18420 3000 18472 3052
rect 18512 3000 18564 3052
rect 19524 3000 19576 3052
rect 20260 3000 20312 3052
rect 21548 3000 21600 3052
rect 11152 2796 11204 2848
rect 14188 2839 14240 2848
rect 14188 2805 14197 2839
rect 14197 2805 14231 2839
rect 14231 2805 14240 2839
rect 14188 2796 14240 2805
rect 15200 2796 15252 2848
rect 18328 2932 18380 2984
rect 20076 2932 20128 2984
rect 19524 2864 19576 2916
rect 19708 2864 19760 2916
rect 21088 2864 21140 2916
rect 19432 2796 19484 2848
rect 19800 2796 19852 2848
rect 20628 2796 20680 2848
rect 20996 2796 21048 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 5540 2592 5592 2644
rect 6000 2592 6052 2644
rect 6276 2635 6328 2644
rect 6276 2601 6285 2635
rect 6285 2601 6319 2635
rect 6319 2601 6328 2635
rect 6276 2592 6328 2601
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 8208 2592 8260 2644
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 11244 2592 11296 2644
rect 12992 2635 13044 2644
rect 3332 2524 3384 2576
rect 2412 2456 2464 2508
rect 5356 2456 5408 2508
rect 5724 2524 5776 2576
rect 10784 2567 10836 2576
rect 10784 2533 10793 2567
rect 10793 2533 10827 2567
rect 10827 2533 10836 2567
rect 10784 2524 10836 2533
rect 11612 2524 11664 2576
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 14740 2592 14792 2644
rect 16304 2592 16356 2644
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 8208 2456 8260 2508
rect 9864 2499 9916 2508
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5908 2388 5960 2440
rect 7104 2388 7156 2440
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 9036 2388 9088 2440
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 12440 2456 12492 2508
rect 14372 2524 14424 2576
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 18788 2635 18840 2644
rect 18788 2601 18797 2635
rect 18797 2601 18831 2635
rect 18831 2601 18840 2635
rect 18788 2592 18840 2601
rect 20076 2592 20128 2644
rect 17408 2524 17460 2576
rect 17868 2524 17920 2576
rect 9956 2388 10008 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12900 2388 12952 2440
rect 14004 2456 14056 2508
rect 14648 2499 14700 2508
rect 14648 2465 14657 2499
rect 14657 2465 14691 2499
rect 14691 2465 14700 2499
rect 14648 2456 14700 2465
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 12624 2363 12676 2372
rect 6184 2252 6236 2304
rect 6828 2252 6880 2304
rect 9680 2252 9732 2304
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 11060 2252 11112 2304
rect 12624 2329 12633 2363
rect 12633 2329 12667 2363
rect 12667 2329 12676 2363
rect 12624 2320 12676 2329
rect 17132 2456 17184 2508
rect 18972 2456 19024 2508
rect 19248 2456 19300 2508
rect 16764 2388 16816 2440
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 18512 2388 18564 2440
rect 15016 2252 15068 2304
rect 22284 2252 22336 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 1492 2048 1544 2100
rect 8208 2048 8260 2100
rect 9680 2048 9732 2100
rect 13912 2048 13964 2100
rect 12164 1980 12216 2032
rect 12900 1980 12952 2032
rect 5356 1912 5408 1964
rect 12992 1912 13044 1964
rect 8392 1844 8444 1896
rect 17132 1844 17184 1896
rect 204 1776 256 1828
rect 8484 1776 8536 1828
rect 11152 1776 11204 1828
rect 5264 1708 5316 1760
rect 9772 1708 9824 1760
rect 16764 1708 16816 1760
rect 1032 1368 1084 1420
rect 8392 1368 8444 1420
rect 3148 1300 3200 1352
rect 5172 1300 5224 1352
rect 10048 1232 10100 1284
rect 16396 1232 16448 1284
rect 13084 552 13136 604
rect 14096 552 14148 604
rect 19340 552 19392 604
rect 19984 552 20036 604
<< metal2 >>
rect 202 22520 258 23000
rect 662 22520 718 23000
rect 1122 22520 1178 23000
rect 1582 22520 1638 23000
rect 1858 22672 1914 22681
rect 1858 22607 1914 22616
rect 216 16726 244 22520
rect 676 19310 704 22520
rect 664 19304 716 19310
rect 664 19246 716 19252
rect 1136 18698 1164 22520
rect 1596 18766 1624 22520
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1780 18902 1808 20334
rect 1872 20058 1900 22607
rect 2042 22520 2098 23000
rect 2594 22520 2650 23000
rect 3054 22520 3110 23000
rect 3514 22520 3570 23000
rect 3974 22520 4030 23000
rect 4434 22520 4490 23000
rect 4986 22520 5042 23000
rect 5446 22520 5502 23000
rect 5906 22520 5962 23000
rect 6366 22520 6422 23000
rect 6826 22520 6882 23000
rect 7378 22520 7434 23000
rect 7838 22520 7894 23000
rect 8298 22520 8354 23000
rect 8758 22520 8814 23000
rect 9218 22520 9274 23000
rect 9770 22520 9826 23000
rect 10230 22520 10286 23000
rect 10690 22520 10746 23000
rect 11150 22520 11206 23000
rect 11702 22520 11758 23000
rect 12162 22522 12218 23000
rect 12162 22520 12480 22522
rect 12622 22520 12678 23000
rect 13082 22520 13138 23000
rect 13542 22520 13598 23000
rect 14094 22520 14150 23000
rect 14554 22520 14610 23000
rect 15014 22520 15070 23000
rect 15474 22520 15530 23000
rect 15934 22520 15990 23000
rect 16486 22520 16542 23000
rect 16946 22520 17002 23000
rect 17406 22520 17462 23000
rect 17866 22520 17922 23000
rect 18326 22520 18382 23000
rect 18878 22520 18934 23000
rect 19338 22520 19394 23000
rect 19798 22520 19854 23000
rect 20258 22520 20314 23000
rect 20442 22672 20498 22681
rect 20442 22607 20498 22616
rect 1950 21176 2006 21185
rect 1950 21111 2006 21120
rect 1964 20602 1992 21111
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 1860 20052 1912 20058
rect 1860 19994 1912 20000
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1872 18970 1900 19751
rect 1950 19272 2006 19281
rect 1950 19207 2006 19216
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1124 18692 1176 18698
rect 1124 18634 1176 18640
rect 1490 18320 1546 18329
rect 1490 18255 1546 18264
rect 1504 17338 1532 18255
rect 1582 17912 1638 17921
rect 1582 17847 1584 17856
rect 1636 17847 1638 17856
rect 1584 17818 1636 17824
rect 1582 17368 1638 17377
rect 1492 17332 1544 17338
rect 1582 17303 1638 17312
rect 1492 17274 1544 17280
rect 1490 16960 1546 16969
rect 1490 16895 1546 16904
rect 204 16720 256 16726
rect 204 16662 256 16668
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 15638 1440 16594
rect 1504 16182 1532 16895
rect 1596 16794 1624 17303
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1688 16561 1716 18770
rect 1964 18426 1992 19207
rect 2056 19009 2084 22520
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2332 19825 2360 19858
rect 2318 19816 2374 19825
rect 2318 19751 2374 19760
rect 2608 19310 2636 22520
rect 2870 22128 2926 22137
rect 2870 22063 2926 22072
rect 2778 20768 2834 20777
rect 2778 20703 2834 20712
rect 2792 20602 2820 20703
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 2792 19922 2820 20266
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2884 19718 2912 22063
rect 2962 21720 3018 21729
rect 2962 21655 3018 21664
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2596 19304 2648 19310
rect 2976 19258 3004 21655
rect 3068 20346 3096 22520
rect 3332 20392 3384 20398
rect 3068 20318 3188 20346
rect 3332 20334 3384 20340
rect 3054 20224 3110 20233
rect 3054 20159 3110 20168
rect 3068 20058 3096 20159
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 2596 19246 2648 19252
rect 2884 19242 3004 19258
rect 2872 19236 3004 19242
rect 2924 19230 3004 19236
rect 2872 19178 2924 19184
rect 3160 19174 3188 20318
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 2042 19000 2098 19009
rect 2042 18935 2098 18944
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1780 17814 1808 18158
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1780 17134 1808 17546
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1674 16552 1730 16561
rect 1674 16487 1730 16496
rect 1952 16448 2004 16454
rect 1674 16416 1730 16425
rect 1952 16390 2004 16396
rect 1674 16351 1730 16360
rect 1492 16176 1544 16182
rect 1492 16118 1544 16124
rect 1688 15706 1716 16351
rect 1964 16153 1992 16390
rect 1950 16144 2006 16153
rect 1950 16079 2006 16088
rect 1858 16008 1914 16017
rect 1858 15943 1914 15952
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1400 15632 1452 15638
rect 1400 15574 1452 15580
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 11218 1440 13262
rect 1504 12986 1532 15506
rect 1872 15162 1900 15943
rect 1950 15464 2006 15473
rect 1950 15399 2006 15408
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1582 14512 1638 14521
rect 1780 14482 1808 14826
rect 1964 14618 1992 15399
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2056 14498 2084 18770
rect 2608 18290 2636 19110
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2792 18426 2820 18799
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2596 18284 2648 18290
rect 2596 18226 2648 18232
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2148 15502 2176 17682
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 1582 14447 1638 14456
rect 1768 14476 1820 14482
rect 1596 14074 1624 14447
rect 1768 14418 1820 14424
rect 1872 14470 2084 14498
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1596 12306 1624 12718
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1780 10810 1808 11494
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 570 3768 626 3777
rect 570 3703 626 3712
rect 204 1828 256 1834
rect 204 1770 256 1776
rect 216 480 244 1770
rect 584 480 612 3703
rect 1688 3505 1716 7958
rect 1872 6662 1900 14470
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2056 13394 2084 14214
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2148 12782 2176 13670
rect 2240 12889 2268 17614
rect 2332 16522 2360 18158
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2516 16697 2544 16730
rect 2884 16726 2912 18090
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2976 16794 3004 16934
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2872 16720 2924 16726
rect 2502 16688 2558 16697
rect 2872 16662 2924 16668
rect 2502 16623 2558 16632
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2516 15366 2544 15846
rect 2608 15745 2636 16526
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2594 15736 2650 15745
rect 2594 15671 2650 15680
rect 2792 15638 2820 15914
rect 2884 15706 2912 16390
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2884 15570 2912 15642
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2976 15366 3004 16050
rect 3068 16046 3096 17274
rect 3160 17066 3188 19110
rect 3238 19000 3294 19009
rect 3238 18935 3240 18944
rect 3292 18935 3294 18944
rect 3240 18906 3292 18912
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3252 17882 3280 18022
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2226 12880 2282 12889
rect 2226 12815 2282 12824
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 2056 12102 2084 12650
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11762 2084 12038
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2240 11558 2268 12310
rect 2332 11898 2360 13670
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 1964 11354 1992 11494
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2240 11150 2268 11494
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10674 2268 11086
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2240 10266 2268 10406
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2424 9738 2452 14418
rect 3068 14278 3096 15982
rect 3160 15706 3188 16526
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3252 15162 3280 16662
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3344 14822 3372 20334
rect 3528 19666 3556 22520
rect 3700 20596 3752 20602
rect 3700 20538 3752 20544
rect 3712 19854 3740 20538
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3804 20058 3832 20334
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3804 19854 3832 19994
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3436 19638 3556 19666
rect 3436 17882 3464 19638
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 18698 3556 19314
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18970 3648 19110
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3528 17678 3556 18634
rect 3712 18290 3740 18702
rect 3700 18284 3752 18290
rect 3620 18244 3700 18272
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3528 15978 3556 17614
rect 3620 17134 3648 18244
rect 3700 18226 3752 18232
rect 3804 18204 3832 19790
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3896 18834 3924 19110
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3884 18216 3936 18222
rect 3804 18176 3884 18204
rect 3884 18158 3936 18164
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3712 17184 3740 17546
rect 3896 17338 3924 18158
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3792 17196 3844 17202
rect 3712 17156 3792 17184
rect 3792 17138 3844 17144
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3620 16590 3648 17070
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3422 15872 3478 15881
rect 3422 15807 3478 15816
rect 3436 15706 3464 15807
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3528 15502 3556 15914
rect 3882 15872 3938 15881
rect 3882 15807 3938 15816
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3436 14464 3464 15098
rect 3514 15056 3570 15065
rect 3804 15026 3832 15438
rect 3514 14991 3570 15000
rect 3792 15020 3844 15026
rect 3528 14618 3556 14991
rect 3792 14962 3844 14968
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3252 14436 3464 14464
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 2778 14104 2834 14113
rect 2778 14039 2834 14048
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2516 12306 2544 13398
rect 2608 13394 2636 13874
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2608 12986 2636 13330
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2516 11694 2544 12242
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2700 10962 2728 11154
rect 2792 11082 2820 14039
rect 3068 13938 3096 14214
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 12374 3004 13806
rect 3068 13462 3096 13874
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3160 12850 3188 13738
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 3068 11218 3096 12582
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2700 10934 2912 10962
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2332 9722 2452 9738
rect 2320 9716 2452 9722
rect 2372 9710 2452 9716
rect 2320 9658 2372 9664
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1964 8430 1992 8978
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2424 8090 2452 9318
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2516 7546 2544 9318
rect 2608 8022 2636 9930
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2700 7886 2728 8298
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2700 7562 2728 7822
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2608 7534 2728 7562
rect 2608 7410 2636 7534
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2700 7206 2728 7414
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1964 6254 1992 6802
rect 2792 6458 2820 6802
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1964 5778 1992 6190
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 2332 5914 2360 6122
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 2332 5234 2360 5850
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2136 5092 2188 5098
rect 2136 5034 2188 5040
rect 2148 4826 2176 5034
rect 2608 5030 2636 5714
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1780 3097 1808 4490
rect 2424 4282 2452 4966
rect 2608 4842 2636 4966
rect 2608 4814 2728 4842
rect 2700 4622 2728 4814
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2700 4214 2728 4558
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2884 4078 2912 10934
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2976 9722 3004 10542
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2976 4554 3004 9658
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3068 8430 3096 9454
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6458 3096 7278
rect 3160 7274 3188 12242
rect 3252 9625 3280 14436
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3238 9616 3294 9625
rect 3238 9551 3294 9560
rect 3344 9450 3372 14282
rect 3620 13870 3648 14758
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3700 13796 3752 13802
rect 3700 13738 3752 13744
rect 3606 13560 3662 13569
rect 3606 13495 3662 13504
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12617 3556 13126
rect 3514 12608 3570 12617
rect 3514 12543 3570 12552
rect 3620 12442 3648 13495
rect 3712 13258 3740 13738
rect 3896 13326 3924 15807
rect 3988 15162 4016 22520
rect 4448 20890 4476 22520
rect 4448 20862 4936 20890
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 19378 4108 19654
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4540 18884 4568 19178
rect 4816 19174 4844 19246
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4620 18896 4672 18902
rect 4540 18856 4620 18884
rect 4620 18838 4672 18844
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4080 16833 4108 18770
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4160 18148 4212 18154
rect 4160 18090 4212 18096
rect 4172 17678 4200 18090
rect 4356 17882 4384 18566
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4908 18465 4936 20862
rect 5000 18630 5028 22520
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19990 5304 20198
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5276 19378 5304 19926
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 4894 18456 4950 18465
rect 4804 18420 4856 18426
rect 4894 18391 4950 18400
rect 4804 18362 4856 18368
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4172 17338 4200 17614
rect 4448 17610 4476 18090
rect 4816 17814 4844 18362
rect 5184 18222 5212 19246
rect 5262 19000 5318 19009
rect 5262 18935 5318 18944
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 4804 17808 4856 17814
rect 4804 17750 4856 17756
rect 4436 17604 4488 17610
rect 4436 17546 4488 17552
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 5184 17202 5212 18158
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5276 17066 5304 18935
rect 5356 18760 5408 18766
rect 5460 18737 5488 22520
rect 5814 19816 5870 19825
rect 5814 19751 5870 19760
rect 5828 19718 5856 19751
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5356 18702 5408 18708
rect 5446 18728 5502 18737
rect 5368 18358 5396 18702
rect 5446 18663 5502 18672
rect 5552 18426 5580 18770
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5356 17672 5408 17678
rect 5408 17632 5488 17660
rect 5356 17614 5408 17620
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4066 16824 4122 16833
rect 4908 16794 4936 16934
rect 4066 16759 4122 16768
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5184 16726 5212 17002
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4080 15706 4108 16594
rect 4172 16250 4200 16594
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4816 16250 4844 16526
rect 5000 16454 5028 16526
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15706 4844 15846
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11665 3464 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3422 11656 3478 11665
rect 3422 11591 3478 11600
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 8974 3280 9318
rect 3344 9178 3372 9386
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8634 3280 8910
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3240 6996 3292 7002
rect 3344 6984 3372 8366
rect 3436 7342 3464 11086
rect 3528 10606 3556 11834
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3620 11150 3648 11562
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3620 10674 3648 11086
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 7478 3556 10542
rect 3620 10062 3648 10610
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3712 7478 3740 12786
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3516 7472 3568 7478
rect 3700 7472 3752 7478
rect 3568 7432 3648 7460
rect 3516 7414 3568 7420
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3292 6956 3372 6984
rect 3240 6938 3292 6944
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3252 5914 3280 6802
rect 3344 6254 3372 6956
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3436 6202 3464 7278
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6322 3556 6598
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3240 5160 3292 5166
rect 3344 5148 3372 6190
rect 3436 6174 3556 6202
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5370 3464 6054
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3292 5120 3372 5148
rect 3240 5102 3292 5108
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2872 4072 2924 4078
rect 2792 4020 2872 4026
rect 2792 4014 2924 4020
rect 2792 3998 2912 4014
rect 2594 3904 2650 3913
rect 2594 3839 2650 3848
rect 2608 3534 2636 3839
rect 2596 3528 2648 3534
rect 1950 3496 2006 3505
rect 2596 3470 2648 3476
rect 1950 3431 1952 3440
rect 2004 3431 2006 3440
rect 1952 3402 2004 3408
rect 1766 3088 1822 3097
rect 1766 3023 1822 3032
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1492 2100 1544 2106
rect 1492 2042 1544 2048
rect 1032 1420 1084 1426
rect 1032 1362 1084 1368
rect 1044 480 1072 1362
rect 1504 480 1532 2042
rect 1964 480 1992 2858
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 2424 480 2452 2450
rect 2792 2145 2820 3998
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2976 3194 3004 3470
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3068 3194 3096 3334
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2870 2816 2926 2825
rect 2870 2751 2926 2760
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 2884 480 2912 2751
rect 3160 2553 3188 5034
rect 3252 4078 3280 5102
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3238 3632 3294 3641
rect 3238 3567 3240 3576
rect 3292 3567 3294 3576
rect 3240 3538 3292 3544
rect 3424 2984 3476 2990
rect 3422 2952 3424 2961
rect 3476 2952 3478 2961
rect 3422 2887 3478 2896
rect 3528 2854 3556 6174
rect 3620 5098 3648 7432
rect 3700 7414 3752 7420
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3620 3602 3648 3878
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3712 3058 3740 7142
rect 3804 4146 3832 12718
rect 3882 12200 3938 12209
rect 3882 12135 3884 12144
rect 3936 12135 3938 12144
rect 3884 12106 3936 12112
rect 3882 10704 3938 10713
rect 3882 10639 3938 10648
rect 3896 10470 3924 10639
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3896 10169 3924 10202
rect 3882 10160 3938 10169
rect 3882 10095 3938 10104
rect 3988 9178 4016 14486
rect 4080 12850 4108 14758
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4264 14074 4292 14554
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12986 4200 13330
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4080 11354 4108 12242
rect 4264 11694 4292 13806
rect 4356 13530 4384 14758
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4816 13802 4844 14214
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4066 11112 4122 11121
rect 4066 11047 4068 11056
rect 4120 11047 4122 11056
rect 4068 11018 4120 11024
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4080 9761 4108 10746
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4172 10130 4200 10542
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4066 9752 4122 9761
rect 4066 9687 4122 9696
rect 4068 9512 4120 9518
rect 4172 9500 4200 10066
rect 4120 9472 4200 9500
rect 4068 9454 4120 9460
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4252 8832 4304 8838
rect 4250 8800 4252 8809
rect 4304 8800 4306 8809
rect 4250 8735 4306 8744
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3896 7886 3924 8298
rect 4068 8288 4120 8294
rect 4066 8256 4068 8265
rect 4120 8256 4122 8265
rect 4356 8242 4384 13262
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4816 12986 4844 13262
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12912 4764 12918
rect 4764 12860 4844 12866
rect 4712 12854 4844 12860
rect 4724 12838 4844 12854
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4540 11558 4568 11630
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4632 11150 4660 11766
rect 4816 11694 4844 12838
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4724 10282 4752 10474
rect 4816 10452 4844 11630
rect 4908 11014 4936 15506
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5000 13326 5028 13806
rect 5092 13530 5120 14758
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10606 4936 10950
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4816 10424 4936 10452
rect 4724 10254 4844 10282
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4816 9382 4844 10254
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4066 8191 4122 8200
rect 4264 8214 4384 8242
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4066 7848 4122 7857
rect 3896 7410 3924 7822
rect 3976 7812 4028 7818
rect 4066 7783 4122 7792
rect 3976 7754 4028 7760
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3896 7002 3924 7346
rect 3988 7313 4016 7754
rect 4080 7546 4108 7783
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3974 7304 4030 7313
rect 3974 7239 4030 7248
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 7002 4200 7142
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4264 6882 4292 8214
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4816 7410 4844 8570
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 3988 6854 4292 6882
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 3988 6361 4016 6854
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3974 6352 4030 6361
rect 3974 6287 4030 6296
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3792 4140 3844 4146
rect 3896 4128 3924 6122
rect 3988 6118 4016 6287
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 4080 5914 4108 6734
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4264 6186 4292 6394
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 5160 4212 5166
rect 3974 5128 4030 5137
rect 4160 5102 4212 5108
rect 3974 5063 4030 5072
rect 3988 4457 4016 5063
rect 4066 4992 4122 5001
rect 4066 4927 4122 4936
rect 4080 4486 4108 4927
rect 4068 4480 4120 4486
rect 3974 4448 4030 4457
rect 4068 4422 4120 4428
rect 3974 4383 4030 4392
rect 4172 4146 4200 5102
rect 4264 5030 4292 5646
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4264 4622 4292 4966
rect 4356 4826 4384 6870
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4816 6440 4844 7346
rect 4724 6412 4844 6440
rect 4724 6254 4752 6412
rect 4908 6361 4936 10424
rect 5000 9110 5028 12174
rect 5092 11286 5120 12378
rect 5184 11354 5212 14758
rect 5276 12782 5304 14894
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5276 11830 5304 12242
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 5092 7721 5120 9318
rect 5276 9160 5304 11494
rect 5368 10470 5396 16526
rect 5460 15502 5488 17632
rect 5552 17338 5580 18022
rect 5644 17814 5672 18226
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5724 17808 5776 17814
rect 5724 17750 5776 17756
rect 5736 17338 5764 17750
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5828 17105 5856 19110
rect 5814 17096 5870 17105
rect 5814 17031 5870 17040
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5552 15745 5580 16594
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5538 15736 5594 15745
rect 5538 15671 5594 15680
rect 5552 15570 5580 15671
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 14822 5488 15438
rect 5736 15026 5764 15982
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5460 13870 5488 14214
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5552 12850 5580 14486
rect 5644 14074 5672 14962
rect 5736 14618 5764 14962
rect 5828 14890 5856 17031
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5736 13530 5764 14214
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5828 13462 5856 14214
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5722 12880 5778 12889
rect 5540 12844 5592 12850
rect 5722 12815 5778 12824
rect 5540 12786 5592 12792
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 9722 5396 10406
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5460 9518 5488 12242
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5644 11937 5672 12174
rect 5630 11928 5686 11937
rect 5630 11863 5686 11872
rect 5644 11762 5672 11863
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11218 5672 11698
rect 5736 11354 5764 12815
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5644 10810 5672 11154
rect 5828 11150 5856 11698
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10266 5580 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5722 9616 5778 9625
rect 5722 9551 5778 9560
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5184 9132 5304 9160
rect 5184 8537 5212 9132
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5276 8634 5304 8978
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5170 8528 5226 8537
rect 5170 8463 5226 8472
rect 5368 8344 5396 8978
rect 5276 8316 5396 8344
rect 5078 7712 5134 7721
rect 5078 7647 5134 7656
rect 5276 7002 5304 8316
rect 5354 7984 5410 7993
rect 5354 7919 5356 7928
rect 5408 7919 5410 7928
rect 5356 7890 5408 7896
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 4894 6352 4950 6361
rect 4894 6287 4950 6296
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4160 4140 4212 4146
rect 3896 4100 4016 4128
rect 3792 4082 3844 4088
rect 3804 4026 3832 4082
rect 3804 3998 3924 4026
rect 3790 3088 3846 3097
rect 3700 3052 3752 3058
rect 3790 3023 3846 3032
rect 3700 2994 3752 3000
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3146 2544 3202 2553
rect 3146 2479 3202 2488
rect 3252 1601 3280 2790
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 3238 1592 3294 1601
rect 3238 1527 3294 1536
rect 3148 1352 3200 1358
rect 3148 1294 3200 1300
rect 3160 649 3188 1294
rect 3146 640 3202 649
rect 3146 575 3202 584
rect 3344 480 3372 2518
rect 3804 480 3832 3023
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1490 0 1546 480
rect 1950 0 2006 480
rect 2410 0 2466 480
rect 2870 0 2926 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 3896 241 3924 3998
rect 3988 3534 4016 4100
rect 4160 4082 4212 4088
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4066 1184 4122 1193
rect 4172 1170 4200 3946
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4122 1142 4200 1170
rect 4066 1119 4122 1128
rect 4264 480 4292 2858
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1442 4844 6190
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5184 4826 5212 5510
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5000 3602 5028 4014
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5000 2990 5028 3538
rect 5184 3346 5212 4558
rect 5276 3890 5304 6938
rect 5368 4622 5396 7890
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5460 4010 5488 9454
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 8498 5672 8910
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5552 8090 5580 8298
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8090 5672 8230
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5736 7002 5764 9551
rect 5920 8809 5948 22520
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6012 18970 6040 20198
rect 6288 19514 6316 20198
rect 6380 20074 6408 22520
rect 6380 20046 6500 20074
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6380 19378 6408 19926
rect 6472 19446 6500 20046
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6460 19440 6512 19446
rect 6460 19382 6512 19388
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6380 18766 6408 19314
rect 6656 19310 6684 19858
rect 6840 19530 6868 22520
rect 7392 20482 7420 22520
rect 7300 20454 7420 20482
rect 7196 20324 7248 20330
rect 7196 20266 7248 20272
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6748 19502 6868 19530
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6368 18760 6420 18766
rect 6748 18714 6776 19502
rect 6828 19440 6880 19446
rect 6828 19382 6880 19388
rect 6840 18986 6868 19382
rect 6932 19242 6960 20198
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6840 18970 7052 18986
rect 6840 18964 7064 18970
rect 6840 18958 7012 18964
rect 7012 18906 7064 18912
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6368 18702 6420 18708
rect 6656 18686 6776 18714
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5998 16144 6054 16153
rect 5998 16079 6054 16088
rect 6012 15910 6040 16079
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 6012 13326 6040 14826
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5906 8800 5962 8809
rect 5906 8735 5962 8744
rect 6012 8650 6040 9862
rect 5920 8622 6040 8650
rect 5814 8256 5870 8265
rect 5814 8191 5870 8200
rect 5828 7954 5856 8191
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5914 5580 6054
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5736 5846 5764 6598
rect 5828 6458 5856 7482
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 5840 5776 5846
rect 5828 5817 5856 6258
rect 5920 6118 5948 8622
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 6012 6866 6040 7958
rect 6104 6934 6132 18566
rect 6656 17377 6684 18686
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6642 17368 6698 17377
rect 6642 17303 6698 17312
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6656 16794 6684 17002
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 16046 6224 16390
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6288 15162 6316 15846
rect 6380 15450 6408 16050
rect 6380 15434 6500 15450
rect 6380 15428 6512 15434
rect 6380 15422 6460 15428
rect 6460 15370 6512 15376
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13530 6224 14350
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6288 11937 6316 14962
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 13802 6408 14758
rect 6472 14074 6500 14894
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6380 12306 6408 13738
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6274 11928 6330 11937
rect 6274 11863 6330 11872
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 10810 6224 11154
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 8673 6224 9318
rect 6182 8664 6238 8673
rect 6182 8599 6238 8608
rect 6288 8004 6316 10950
rect 6380 10266 6408 11086
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9586 6408 10066
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6368 8016 6420 8022
rect 6288 7976 6368 8004
rect 6368 7958 6420 7964
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7546 6224 7686
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6196 6769 6224 6938
rect 6276 6792 6328 6798
rect 6182 6760 6238 6769
rect 6092 6724 6144 6730
rect 6276 6734 6328 6740
rect 6182 6695 6238 6704
rect 6092 6666 6144 6672
rect 6000 6248 6052 6254
rect 5998 6216 6000 6225
rect 6052 6216 6054 6225
rect 5998 6151 6054 6160
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5724 5782 5776 5788
rect 5814 5808 5870 5817
rect 5814 5743 5870 5752
rect 5828 5710 5856 5743
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5828 5166 5856 5646
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5276 3862 5488 3890
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5092 3318 5212 3346
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4724 1414 4844 1442
rect 4724 480 4752 1414
rect 5092 480 5120 3318
rect 5276 3194 5304 3470
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5460 2938 5488 3862
rect 5552 3602 5580 4558
rect 5644 3942 5672 4626
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5644 3534 5672 3878
rect 5736 3738 5764 4966
rect 5920 4729 5948 6054
rect 6104 5914 6132 6666
rect 6288 6322 6316 6734
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5914 6408 6054
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5906 4720 5962 4729
rect 5906 4655 5962 4664
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5724 3392 5776 3398
rect 5630 3360 5686 3369
rect 6012 3380 6040 5714
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6104 5166 6132 5510
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5724 3334 5776 3340
rect 5828 3352 6040 3380
rect 5630 3295 5686 3304
rect 5184 2910 5488 2938
rect 5540 2916 5592 2922
rect 5184 1358 5212 2910
rect 5540 2858 5592 2864
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5276 2446 5304 2790
rect 5552 2650 5580 2858
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5276 1766 5304 2382
rect 5368 1970 5396 2450
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 5264 1760 5316 1766
rect 5264 1702 5316 1708
rect 5644 1442 5672 3295
rect 5736 2582 5764 3334
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5828 2292 5856 3352
rect 6104 3210 6132 3674
rect 6184 3664 6236 3670
rect 6182 3632 6184 3641
rect 6236 3632 6238 3641
rect 6182 3567 6238 3576
rect 5920 3182 6132 3210
rect 5920 2446 5948 3182
rect 6288 2854 6316 2885
rect 6000 2848 6052 2854
rect 6276 2848 6328 2854
rect 6000 2790 6052 2796
rect 6274 2816 6276 2825
rect 6328 2816 6330 2825
rect 6012 2650 6040 2790
rect 6274 2751 6330 2760
rect 6288 2650 6316 2751
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6196 2310 6224 2450
rect 6184 2304 6236 2310
rect 5828 2264 6040 2292
rect 5552 1414 5672 1442
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5552 480 5580 1414
rect 6012 480 6040 2264
rect 6184 2246 6236 2252
rect 6472 480 6500 13398
rect 6564 9926 6592 14282
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6656 9178 6684 15098
rect 6748 12073 6776 18566
rect 6840 18426 6868 18770
rect 7208 18630 7236 20266
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 17134 6868 17478
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6828 16244 6880 16250
rect 6932 16232 6960 17002
rect 6880 16204 6960 16232
rect 6828 16186 6880 16192
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6840 15094 6868 15914
rect 6932 15570 6960 16050
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14618 6868 14758
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6932 14482 6960 15098
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7024 14362 7052 18022
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7116 16289 7144 16526
rect 7102 16280 7158 16289
rect 7102 16215 7158 16224
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7116 14600 7144 15098
rect 7208 14793 7236 18566
rect 7194 14784 7250 14793
rect 7194 14719 7250 14728
rect 7116 14572 7236 14600
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 6932 14334 7052 14362
rect 6828 13456 6880 13462
rect 6932 13433 6960 14334
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6828 13398 6880 13404
rect 6918 13424 6974 13433
rect 6840 13297 6868 13398
rect 6918 13359 6974 13368
rect 6826 13288 6882 13297
rect 6826 13223 6882 13232
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 6748 10538 6776 11999
rect 6918 11656 6974 11665
rect 6918 11591 6974 11600
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11218 6868 11494
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6932 11098 6960 11591
rect 6840 11070 6960 11098
rect 7024 11082 7052 13806
rect 7116 13530 7144 14418
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7208 11801 7236 14572
rect 7300 14249 7328 20454
rect 7380 20392 7432 20398
rect 7852 20346 7880 22520
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 7380 20334 7432 20340
rect 7392 20058 7420 20334
rect 7484 20318 7880 20346
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7392 17882 7420 18702
rect 7484 18154 7512 20318
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8220 20058 8248 20402
rect 8312 20346 8340 22520
rect 8312 20318 8432 20346
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7668 19281 7696 19790
rect 7654 19272 7710 19281
rect 7564 19236 7616 19242
rect 8220 19258 8248 19994
rect 8312 19514 8340 20198
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8128 19242 8248 19258
rect 7654 19207 7710 19216
rect 8116 19236 8248 19242
rect 7564 19178 7616 19184
rect 7576 18766 7604 19178
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7576 18290 7604 18702
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 17513 7512 17614
rect 7470 17504 7526 17513
rect 7470 17439 7526 17448
rect 7378 17232 7434 17241
rect 7378 17167 7380 17176
rect 7432 17167 7434 17176
rect 7380 17138 7432 17144
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16794 7420 16934
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7392 16425 7420 16458
rect 7378 16416 7434 16425
rect 7378 16351 7434 16360
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7286 14240 7342 14249
rect 7286 14175 7342 14184
rect 7392 13326 7420 14962
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7392 12209 7420 12718
rect 7378 12200 7434 12209
rect 7378 12135 7434 12144
rect 7380 11824 7432 11830
rect 7194 11792 7250 11801
rect 7380 11766 7432 11772
rect 7194 11727 7250 11736
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7208 11354 7236 11494
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7012 11076 7064 11082
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6552 8968 6604 8974
rect 6550 8936 6552 8945
rect 6604 8936 6606 8945
rect 6550 8871 6606 8880
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 6934 6684 7142
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6564 6458 6592 6870
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6656 6338 6684 6734
rect 6564 6310 6684 6338
rect 6564 3210 6592 6310
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5166 6684 6054
rect 6748 5914 6776 9658
rect 6840 9110 6868 11070
rect 7012 11018 7064 11024
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 9586 6960 10474
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7024 9518 7052 10406
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7012 9512 7064 9518
rect 6918 9480 6974 9489
rect 7012 9454 7064 9460
rect 6918 9415 6974 9424
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 7886 6868 8910
rect 6932 7954 6960 9415
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6932 7732 6960 7890
rect 6840 7704 6960 7732
rect 6840 6798 6868 7704
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6840 5642 6868 6258
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6748 3942 6776 4150
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6734 3224 6790 3233
rect 6564 3182 6734 3210
rect 6734 3159 6790 3168
rect 6748 2122 6776 3159
rect 6840 2310 6868 3674
rect 6932 3194 6960 7210
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6828 2304 6880 2310
rect 7024 2292 7052 9046
rect 7116 8430 7144 10202
rect 7208 9654 7236 10406
rect 7300 9654 7328 11494
rect 7392 11354 7420 11766
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7484 11014 7512 17439
rect 7668 17202 7696 19207
rect 8168 19230 8248 19236
rect 8116 19178 8168 19184
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18426 7788 19110
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7944 18222 7972 18702
rect 8220 18630 8248 18770
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18222 8340 18566
rect 8404 18426 8432 20318
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8680 18698 8708 19110
rect 8772 18698 8800 22520
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8864 18902 8892 20198
rect 9232 20074 9260 22520
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 8956 20046 9260 20074
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7760 17785 7788 17818
rect 7746 17776 7802 17785
rect 7746 17711 7802 17720
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7576 16046 7604 17138
rect 7668 16658 7696 17138
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7668 16250 7696 16594
rect 7930 16552 7986 16561
rect 7930 16487 7986 16496
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15706 7604 15982
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7668 15094 7696 16186
rect 7944 15978 7972 16487
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8208 15360 8260 15366
rect 8022 15328 8078 15337
rect 8208 15302 8260 15308
rect 8022 15263 8078 15272
rect 7838 15192 7894 15201
rect 7838 15127 7840 15136
rect 7892 15127 7894 15136
rect 7840 15098 7892 15104
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7576 13530 7604 15030
rect 7668 13802 7696 15030
rect 8036 14958 8064 15263
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7564 13524 7616 13530
rect 8220 13512 8248 15302
rect 8312 14958 8340 17478
rect 8404 16250 8432 18022
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8496 15858 8524 18090
rect 8666 17912 8722 17921
rect 8956 17864 8984 20046
rect 9324 19990 9352 20402
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 8666 17847 8722 17856
rect 8680 17746 8708 17847
rect 8772 17836 8984 17864
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16726 8616 17070
rect 8576 16720 8628 16726
rect 8668 16720 8720 16726
rect 8576 16662 8628 16668
rect 8666 16688 8668 16697
rect 8720 16688 8722 16697
rect 8588 16182 8616 16662
rect 8666 16623 8722 16632
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8404 15830 8524 15858
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8404 15065 8432 15830
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8390 15056 8446 15065
rect 8496 15026 8524 15642
rect 8390 14991 8446 15000
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8404 14074 8432 14894
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8496 14521 8524 14758
rect 8574 14648 8630 14657
rect 8574 14583 8630 14592
rect 8482 14512 8538 14521
rect 8482 14447 8538 14456
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8300 13524 8352 13530
rect 8220 13484 8300 13512
rect 7564 13466 7616 13472
rect 8300 13466 8352 13472
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 11150 7604 12582
rect 7668 11898 7696 13398
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 7852 12714 7880 13262
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8220 12442 8248 13262
rect 8404 12782 8432 13738
rect 8496 12986 8524 14350
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7746 12336 7802 12345
rect 7746 12271 7802 12280
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7654 11792 7710 11801
rect 7654 11727 7710 11736
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7392 10198 7420 10610
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7484 9874 7512 10610
rect 7392 9846 7512 9874
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7392 9466 7420 9846
rect 7470 9752 7526 9761
rect 7576 9722 7604 11086
rect 7470 9687 7526 9696
rect 7564 9716 7616 9722
rect 7208 9438 7420 9466
rect 7484 9450 7512 9687
rect 7564 9658 7616 9664
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7472 9444 7524 9450
rect 7208 8634 7236 9438
rect 7472 9386 7524 9392
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 9042 7420 9318
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7484 8922 7512 9386
rect 7300 8894 7512 8922
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7194 8528 7250 8537
rect 7194 8463 7250 8472
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7208 7936 7236 8463
rect 7116 7908 7236 7936
rect 7116 5914 7144 7908
rect 7194 7848 7250 7857
rect 7194 7783 7196 7792
rect 7248 7783 7250 7792
rect 7196 7754 7248 7760
rect 7208 6254 7236 7754
rect 7300 6730 7328 8894
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7208 5574 7236 6054
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7194 5264 7250 5273
rect 7194 5199 7250 5208
rect 7208 5098 7236 5199
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7116 4554 7144 5034
rect 7300 4826 7328 5510
rect 7392 5409 7420 7958
rect 7484 7206 7512 8366
rect 7576 7750 7604 9454
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7378 5400 7434 5409
rect 7484 5370 7512 7142
rect 7576 7002 7604 7210
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7668 6848 7696 11727
rect 7760 9926 7788 12271
rect 7838 12200 7894 12209
rect 7838 12135 7894 12144
rect 7852 11762 7880 12135
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 8220 11626 8248 12378
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7852 10606 7880 11018
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8220 10266 8248 11222
rect 8312 10826 8340 12650
rect 8496 12374 8524 12922
rect 8588 12714 8616 14583
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8496 11898 8524 12310
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11898 8616 12174
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8680 11626 8708 15846
rect 8772 15337 8800 17836
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8758 15328 8814 15337
rect 8758 15263 8814 15272
rect 8772 15026 8800 15263
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8864 14618 8892 17682
rect 8942 16416 8998 16425
rect 8942 16351 8998 16360
rect 8956 16250 8984 16351
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 9048 15638 9076 19858
rect 9324 19378 9352 19926
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9220 19304 9272 19310
rect 9218 19272 9220 19281
rect 9272 19272 9274 19281
rect 9218 19207 9274 19216
rect 9324 18766 9352 19314
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9140 18426 9168 18566
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 15632 9088 15638
rect 9036 15574 9088 15580
rect 8944 15496 8996 15502
rect 9140 15484 9168 17614
rect 9232 17270 9260 17682
rect 9324 17610 9352 18702
rect 9416 17921 9444 20266
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9586 19272 9642 19281
rect 9402 17912 9458 17921
rect 9402 17847 9458 17856
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9232 16833 9260 17206
rect 9218 16824 9274 16833
rect 9218 16759 9274 16768
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 8996 15456 9168 15484
rect 8944 15438 8996 15444
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8772 14521 8800 14554
rect 8758 14512 8814 14521
rect 8758 14447 8814 14456
rect 8956 14414 8984 15438
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8944 14408 8996 14414
rect 8758 14376 8814 14385
rect 8944 14350 8996 14356
rect 8758 14311 8814 14320
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8312 10798 8524 10826
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7748 9920 7800 9926
rect 8404 9897 8432 10406
rect 7748 9862 7800 9868
rect 8390 9888 8446 9897
rect 7760 8265 7788 9862
rect 8390 9823 8446 9832
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8128 9364 8156 9658
rect 8390 9616 8446 9625
rect 8390 9551 8446 9560
rect 8404 9450 8432 9551
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8128 9336 8248 9364
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8036 8809 8064 9046
rect 8022 8800 8078 8809
rect 8022 8735 8078 8744
rect 7746 8256 7802 8265
rect 7746 8191 7802 8200
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 8220 7954 8248 9336
rect 8298 9344 8354 9353
rect 8298 9279 8354 9288
rect 8312 8838 8340 9279
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8404 8650 8432 9143
rect 8496 9058 8524 10798
rect 8588 10266 8616 10950
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8772 9432 8800 14311
rect 8852 14272 8904 14278
rect 8944 14272 8996 14278
rect 8852 14214 8904 14220
rect 8942 14240 8944 14249
rect 8996 14240 8998 14249
rect 8864 13530 8892 14214
rect 8942 14175 8998 14184
rect 8956 13734 8984 14175
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8763 9404 8800 9432
rect 8668 9376 8720 9382
rect 8666 9344 8668 9353
rect 8720 9344 8722 9353
rect 8666 9279 8722 9288
rect 8763 9194 8791 9404
rect 8763 9166 8800 9194
rect 8496 9030 8616 9058
rect 8300 8628 8352 8634
rect 8404 8622 8524 8650
rect 8300 8570 8352 8576
rect 8312 8090 8340 8570
rect 8496 8362 8524 8622
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8300 8084 8352 8090
rect 8352 8044 8432 8072
rect 8300 8026 8352 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7852 7721 7880 7822
rect 7838 7712 7894 7721
rect 7838 7647 7894 7656
rect 8036 7546 8064 7822
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7760 7313 7788 7346
rect 7746 7304 7802 7313
rect 7746 7239 7802 7248
rect 7576 6820 7696 6848
rect 7378 5335 7434 5344
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7470 5264 7526 5273
rect 7470 5199 7526 5208
rect 7484 5030 7512 5199
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 2446 7144 4490
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 4146 7236 4422
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7484 4010 7512 4966
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7286 3904 7342 3913
rect 7208 3194 7236 3878
rect 7286 3839 7342 3848
rect 7300 3602 7328 3839
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7300 3126 7328 3334
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7392 2650 7420 3946
rect 7484 3534 7512 3946
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7024 2264 7420 2292
rect 6828 2246 6880 2252
rect 6748 2094 6960 2122
rect 6932 480 6960 2094
rect 7392 480 7420 2264
rect 7576 1884 7604 6820
rect 7760 6118 7788 7239
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8312 6458 8340 7142
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8220 6338 8248 6394
rect 8220 6310 8340 6338
rect 8312 6186 8340 6310
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5778 7788 6054
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7930 5808 7986 5817
rect 7748 5772 7800 5778
rect 7930 5743 7986 5752
rect 7748 5714 7800 5720
rect 7944 5574 7972 5743
rect 7748 5568 7800 5574
rect 7746 5536 7748 5545
rect 7932 5568 7984 5574
rect 7800 5536 7802 5545
rect 7932 5510 7984 5516
rect 7746 5471 7802 5480
rect 8220 5370 8248 6122
rect 8404 6118 8432 8044
rect 8496 7954 8524 8298
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8588 7698 8616 9030
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8680 8090 8708 8842
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8496 7670 8616 7698
rect 8496 7449 8524 7670
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8482 7440 8538 7449
rect 8482 7375 8538 7384
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5840 8352 5846
rect 8298 5808 8300 5817
rect 8352 5808 8354 5817
rect 8298 5743 8354 5752
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8312 5370 8340 5646
rect 8404 5642 8432 6054
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8404 5273 8432 5578
rect 8390 5264 8446 5273
rect 8300 5228 8352 5234
rect 8390 5199 8446 5208
rect 8300 5170 8352 5176
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4622 7788 5034
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8312 4865 8340 5170
rect 8588 5001 8616 7482
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 7002 8708 7142
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8772 6780 8800 9166
rect 8864 7449 8892 13330
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8956 10198 8984 12242
rect 9048 11744 9076 15302
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 13870 9168 14758
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9232 13530 9260 16526
rect 9324 16454 9352 17546
rect 9416 17338 9444 17682
rect 9508 17678 9536 19246
rect 9586 19207 9642 19216
rect 9600 18850 9628 19207
rect 9600 18834 9720 18850
rect 9588 18828 9720 18834
rect 9640 18822 9720 18828
rect 9588 18770 9640 18776
rect 9496 17672 9548 17678
rect 9692 17649 9720 18822
rect 9496 17614 9548 17620
rect 9678 17640 9734 17649
rect 9678 17575 9734 17584
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 16114 9352 16390
rect 9586 16280 9642 16289
rect 9586 16215 9642 16224
rect 9600 16114 9628 16215
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9496 16040 9548 16046
rect 9494 16008 9496 16017
rect 9548 16008 9550 16017
rect 9494 15943 9550 15952
rect 9600 15144 9628 16050
rect 9692 15570 9720 16934
rect 9784 16017 9812 22520
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9876 20058 9904 20742
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9968 19514 9996 20470
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9876 16182 9904 18634
rect 10152 18601 10180 18702
rect 10138 18592 10194 18601
rect 10138 18527 10194 18536
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9770 16008 9826 16017
rect 9770 15943 9826 15952
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9508 15116 9720 15144
rect 9508 15065 9536 15116
rect 9494 15056 9550 15065
rect 9692 15026 9720 15116
rect 9494 14991 9550 15000
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9310 14920 9366 14929
rect 9310 14855 9366 14864
rect 9324 13802 9352 14855
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9508 14346 9536 14758
rect 9600 14618 9628 14962
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9416 13394 9444 13942
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9140 12209 9168 12242
rect 9232 12238 9260 12650
rect 9220 12232 9272 12238
rect 9126 12200 9182 12209
rect 9220 12174 9272 12180
rect 9126 12135 9182 12144
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9048 11716 9168 11744
rect 9140 11665 9168 11716
rect 9126 11656 9182 11665
rect 9036 11620 9088 11626
rect 9126 11591 9182 11600
rect 9036 11562 9088 11568
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8956 9178 8984 9590
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8956 8362 8984 8978
rect 9048 8537 9076 11562
rect 9218 10840 9274 10849
rect 9218 10775 9220 10784
rect 9272 10775 9274 10784
rect 9220 10746 9272 10752
rect 9220 10668 9272 10674
rect 9140 10628 9220 10656
rect 9140 10538 9168 10628
rect 9220 10610 9272 10616
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 9034 8528 9090 8537
rect 9034 8463 9090 8472
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8850 7440 8906 7449
rect 8956 7410 8984 8298
rect 9034 7712 9090 7721
rect 9034 7647 9090 7656
rect 8850 7375 8906 7384
rect 8944 7404 8996 7410
rect 8864 7274 8892 7375
rect 8944 7346 8996 7352
rect 8942 7304 8998 7313
rect 8852 7268 8904 7274
rect 8942 7239 8998 7248
rect 8852 7210 8904 7216
rect 8956 7002 8984 7239
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8944 6792 8996 6798
rect 8772 6752 8944 6780
rect 8944 6734 8996 6740
rect 8666 6352 8722 6361
rect 8666 6287 8722 6296
rect 8680 6089 8708 6287
rect 8956 6186 8984 6734
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8666 6080 8722 6089
rect 9048 6066 9076 7647
rect 9140 7546 9168 10134
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 7002 9168 7278
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8666 6015 8722 6024
rect 8772 6038 9076 6066
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8390 4992 8446 5001
rect 8390 4927 8446 4936
rect 8574 4992 8630 5001
rect 8574 4927 8630 4936
rect 8298 4856 8354 4865
rect 8298 4791 8354 4800
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7668 3058 7696 4422
rect 7760 4282 7788 4558
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7760 3398 7788 4218
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3058 7788 3334
rect 7944 3194 7972 3470
rect 8312 3398 8340 4422
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8404 3210 8432 4927
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8484 4616 8536 4622
rect 8588 4593 8616 4626
rect 8680 4622 8708 5714
rect 8668 4616 8720 4622
rect 8484 4558 8536 4564
rect 8574 4584 8630 4593
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8312 3182 8432 3210
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8220 2650 8248 2858
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8220 2106 8248 2450
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 7576 1856 7880 1884
rect 7852 480 7880 1856
rect 8312 480 8340 3182
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8404 1902 8432 2382
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 8404 1426 8432 1838
rect 8496 1834 8524 4558
rect 8668 4558 8720 4564
rect 8574 4519 8630 4528
rect 8588 3641 8616 4519
rect 8574 3632 8630 3641
rect 8574 3567 8630 3576
rect 8576 3052 8628 3058
rect 8772 3040 8800 6038
rect 9140 5710 9168 6734
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8850 5536 8906 5545
rect 8850 5471 8906 5480
rect 9126 5536 9182 5545
rect 9126 5471 9182 5480
rect 8864 4622 8892 5471
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8864 4282 8892 4558
rect 8956 4282 8984 4966
rect 9048 4826 9076 5306
rect 9140 5234 9168 5471
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9140 4758 9168 4966
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8628 3012 8800 3040
rect 8576 2994 8628 3000
rect 8864 2088 8892 4082
rect 9048 2446 9076 4150
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8772 2060 8892 2088
rect 8484 1828 8536 1834
rect 8484 1770 8536 1776
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8772 480 8800 2060
rect 9232 480 9260 10474
rect 9324 9586 9352 12106
rect 9416 10538 9444 13194
rect 9600 12918 9628 13874
rect 9692 13530 9720 14418
rect 9784 13802 9812 15846
rect 9968 13938 9996 16730
rect 10060 15162 10088 16934
rect 10152 15473 10180 18362
rect 10138 15464 10194 15473
rect 10138 15399 10194 15408
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9968 13394 9996 13466
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10060 12986 10088 14486
rect 10152 14482 10180 15030
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9588 12912 9640 12918
rect 10152 12866 10180 13126
rect 9588 12854 9640 12860
rect 9600 12238 9628 12854
rect 10060 12838 10180 12866
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9494 11928 9550 11937
rect 9494 11863 9550 11872
rect 9508 11830 9536 11863
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9692 11529 9720 12718
rect 9956 12640 10008 12646
rect 9876 12600 9956 12628
rect 9772 11552 9824 11558
rect 9678 11520 9734 11529
rect 9772 11494 9824 11500
rect 9678 11455 9734 11464
rect 9588 11280 9640 11286
rect 9586 11248 9588 11257
rect 9640 11248 9642 11257
rect 9586 11183 9642 11192
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9600 10470 9628 11086
rect 9692 10810 9720 11154
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9588 10464 9640 10470
rect 9402 10432 9458 10441
rect 9588 10406 9640 10412
rect 9402 10367 9458 10376
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9416 9058 9444 10367
rect 9600 9994 9628 10406
rect 9784 10130 9812 11494
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9324 9030 9444 9058
rect 9324 5778 9352 9030
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8634 9444 8910
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9402 8528 9458 8537
rect 9402 8463 9458 8472
rect 9416 7206 9444 8463
rect 9508 8430 9536 9522
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9600 8634 9628 9046
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 7410 9536 8366
rect 9600 7886 9628 8570
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9692 7585 9720 8978
rect 9784 8906 9812 9318
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9770 8392 9826 8401
rect 9770 8327 9826 8336
rect 9784 8265 9812 8327
rect 9770 8256 9826 8265
rect 9770 8191 9826 8200
rect 9784 8022 9812 8191
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9678 7576 9734 7585
rect 9678 7511 9734 7520
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9324 5098 9352 5306
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9416 5001 9444 7142
rect 9508 6730 9536 7346
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9680 7336 9732 7342
rect 9784 7313 9812 7822
rect 9680 7278 9732 7284
rect 9770 7304 9826 7313
rect 9600 6798 9628 7278
rect 9692 6905 9720 7278
rect 9770 7239 9826 7248
rect 9678 6896 9734 6905
rect 9678 6831 9734 6840
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9508 6390 9536 6666
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9692 6202 9720 6394
rect 9600 6174 9720 6202
rect 9600 6118 9628 6174
rect 9588 6112 9640 6118
rect 9494 6080 9550 6089
rect 9588 6054 9640 6060
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9494 6015 9550 6024
rect 9508 5778 9536 6015
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9508 5166 9536 5714
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5234 9628 5510
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9402 4992 9458 5001
rect 9402 4927 9458 4936
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9600 4282 9628 4490
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9324 4010 9352 4150
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9324 3466 9352 3946
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9600 480 9628 2790
rect 9692 2394 9720 6054
rect 9784 4078 9812 7239
rect 9876 4146 9904 12600
rect 9956 12582 10008 12588
rect 10060 12170 10088 12838
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9954 11928 10010 11937
rect 9954 11863 10010 11872
rect 9968 9722 9996 11863
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10046 11384 10102 11393
rect 10046 11319 10102 11328
rect 10060 11286 10088 11319
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10060 9602 10088 10950
rect 10152 10674 10180 11698
rect 10244 11150 10272 22520
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10704 20482 10732 22520
rect 11060 20528 11112 20534
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10428 19310 10456 20402
rect 10612 19990 10640 20470
rect 10704 20454 10824 20482
rect 11060 20470 11112 20476
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10704 18698 10732 20334
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10508 18080 10560 18086
rect 10692 18080 10744 18086
rect 10508 18022 10560 18028
rect 10612 18028 10692 18034
rect 10612 18022 10744 18028
rect 10322 17232 10378 17241
rect 10322 17167 10378 17176
rect 10336 15609 10364 17167
rect 10428 16794 10456 18022
rect 10520 17814 10548 18022
rect 10612 18006 10732 18022
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10612 17660 10640 18006
rect 10520 17632 10640 17660
rect 10692 17672 10744 17678
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10428 15745 10456 15914
rect 10414 15736 10470 15745
rect 10414 15671 10470 15680
rect 10322 15600 10378 15609
rect 10322 15535 10378 15544
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10428 14958 10456 15506
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10336 13462 10364 13942
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12850 10364 13262
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10428 12238 10456 14894
rect 10520 13190 10548 17632
rect 10692 17614 10744 17620
rect 10704 17338 10732 17614
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10704 15706 10732 16390
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10598 15600 10654 15609
rect 10796 15586 10824 20454
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10980 19990 11008 20402
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 11072 19514 11100 20470
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11164 19394 11192 22520
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11716 20346 11744 22520
rect 12176 22494 12480 22520
rect 11716 20318 11836 20346
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11348 20058 11376 20198
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11428 19440 11480 19446
rect 11164 19366 11376 19394
rect 11428 19382 11480 19388
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10598 15535 10654 15544
rect 10704 15558 10824 15586
rect 10612 13530 10640 15535
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10612 12102 10640 12582
rect 10600 12096 10652 12102
rect 10414 12064 10470 12073
rect 10600 12038 10652 12044
rect 10414 11999 10470 12008
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10336 11694 10364 11766
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10232 11144 10284 11150
rect 10336 11121 10364 11154
rect 10232 11086 10284 11092
rect 10322 11112 10378 11121
rect 10322 11047 10378 11056
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10266 10272 10406
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10060 9574 10364 9602
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9968 4826 9996 9454
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10230 9344 10286 9353
rect 10046 8392 10102 8401
rect 10046 8327 10102 8336
rect 10060 7721 10088 8327
rect 10046 7712 10102 7721
rect 10046 7647 10102 7656
rect 10046 7576 10102 7585
rect 10046 7511 10102 7520
rect 10060 7206 10088 7511
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10152 6866 10180 9318
rect 10230 9279 10286 9288
rect 10244 9178 10272 9279
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6254 10088 6734
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5914 10088 6054
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10244 5817 10272 8366
rect 10230 5808 10286 5817
rect 10230 5743 10286 5752
rect 10336 5658 10364 9574
rect 10428 7274 10456 11999
rect 10704 11937 10732 15558
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10796 14958 10824 15438
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10796 13938 10824 14418
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10690 11928 10746 11937
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10600 11892 10652 11898
rect 10690 11863 10746 11872
rect 10600 11834 10652 11840
rect 10520 11801 10548 11834
rect 10506 11792 10562 11801
rect 10506 11727 10562 11736
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10520 8838 10548 11086
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8129 10548 8774
rect 10612 8673 10640 11834
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 9722 10732 11630
rect 10796 11558 10824 13466
rect 10888 11694 10916 18770
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10980 18306 11008 18702
rect 11072 18426 11100 18770
rect 11164 18766 11192 19178
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11256 18873 11284 19110
rect 11242 18864 11298 18873
rect 11242 18799 11298 18808
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 11164 18358 11192 18702
rect 11348 18612 11376 19366
rect 11440 19009 11468 19382
rect 11610 19136 11666 19145
rect 11610 19071 11666 19080
rect 11624 19009 11652 19071
rect 11426 19000 11482 19009
rect 11426 18935 11482 18944
rect 11610 19000 11666 19009
rect 11610 18935 11666 18944
rect 11716 18630 11744 20198
rect 11808 19666 11836 20318
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11808 19638 11928 19666
rect 11796 19168 11848 19174
rect 11794 19136 11796 19145
rect 11848 19136 11850 19145
rect 11794 19071 11850 19080
rect 11256 18584 11376 18612
rect 11704 18624 11756 18630
rect 11152 18352 11204 18358
rect 10980 18290 11100 18306
rect 11152 18294 11204 18300
rect 10980 18284 11112 18290
rect 10980 18278 11060 18284
rect 11060 18226 11112 18232
rect 10966 18048 11022 18057
rect 10966 17983 11022 17992
rect 10980 17513 11008 17983
rect 11072 17746 11100 18226
rect 11164 17882 11192 18294
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11058 17640 11114 17649
rect 11058 17575 11114 17584
rect 11072 17542 11100 17575
rect 11060 17536 11112 17542
rect 10966 17504 11022 17513
rect 11060 17478 11112 17484
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 10966 17439 11022 17448
rect 11164 17377 11192 17478
rect 11150 17368 11206 17377
rect 11060 17332 11112 17338
rect 11150 17303 11206 17312
rect 11060 17274 11112 17280
rect 11072 17134 11100 17274
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10980 14550 11008 16526
rect 11072 15201 11100 17070
rect 11152 16992 11204 16998
rect 11150 16960 11152 16969
rect 11204 16960 11206 16969
rect 11150 16895 11206 16904
rect 11150 16552 11206 16561
rect 11150 16487 11206 16496
rect 11164 16250 11192 16487
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11152 16040 11204 16046
rect 11150 16008 11152 16017
rect 11204 16008 11206 16017
rect 11150 15943 11206 15952
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15609 11192 15846
rect 11150 15600 11206 15609
rect 11150 15535 11206 15544
rect 11058 15192 11114 15201
rect 11058 15127 11114 15136
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10980 13190 11008 14486
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 11830 11008 12582
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10980 11694 11008 11766
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10796 10305 10824 11494
rect 10782 10296 10838 10305
rect 10782 10231 10838 10240
rect 10782 10160 10838 10169
rect 10782 10095 10838 10104
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10598 8664 10654 8673
rect 10598 8599 10654 8608
rect 10612 8362 10640 8599
rect 10704 8537 10732 9522
rect 10690 8528 10746 8537
rect 10690 8463 10746 8472
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10506 8120 10562 8129
rect 10506 8055 10562 8064
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10506 7712 10562 7721
rect 10506 7647 10562 7656
rect 10520 7342 10548 7647
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10612 7274 10640 7822
rect 10704 7478 10732 8463
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10428 6458 10456 6938
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10244 5630 10364 5658
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10244 5114 10272 5630
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10336 5234 10364 5510
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10152 5012 10180 5102
rect 10244 5086 10364 5114
rect 10152 4984 10272 5012
rect 10244 4865 10272 4984
rect 10230 4856 10286 4865
rect 9956 4820 10008 4826
rect 10230 4791 10286 4800
rect 9956 4762 10008 4768
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9784 3194 9812 3470
rect 9876 3194 9904 3538
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9862 2544 9918 2553
rect 9862 2479 9864 2488
rect 9916 2479 9918 2488
rect 9864 2450 9916 2456
rect 9968 2446 9996 4490
rect 10060 2854 10088 4694
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10152 3777 10180 4626
rect 10244 4622 10272 4791
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10230 4448 10286 4457
rect 10230 4383 10286 4392
rect 10244 3913 10272 4383
rect 10336 4185 10364 5086
rect 10428 5030 10456 5850
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10322 4176 10378 4185
rect 10322 4111 10378 4120
rect 10230 3904 10286 3913
rect 10230 3839 10286 3848
rect 10138 3768 10194 3777
rect 10138 3703 10194 3712
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10244 2689 10272 3839
rect 10230 2680 10286 2689
rect 10230 2615 10286 2624
rect 9956 2440 10008 2446
rect 9692 2366 9812 2394
rect 9956 2382 10008 2388
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 2106 9720 2246
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9784 1766 9812 2366
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 10060 1290 10088 2246
rect 10048 1284 10100 1290
rect 10048 1226 10100 1232
rect 10336 1170 10364 4111
rect 10428 3516 10456 4966
rect 10520 4214 10548 7142
rect 10704 6798 10732 7278
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6390 10732 6734
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10796 6225 10824 10095
rect 10888 7886 10916 11494
rect 11072 10826 11100 13262
rect 11164 12986 11192 13330
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12646 11284 18584
rect 11704 18566 11756 18572
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 11348 17882 11376 18090
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11716 17202 11744 18090
rect 11900 18034 11928 19638
rect 11992 19514 12020 19790
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11992 18766 12020 19450
rect 12268 19417 12296 19654
rect 12360 19446 12388 19654
rect 12348 19440 12400 19446
rect 12254 19408 12310 19417
rect 12348 19382 12400 19388
rect 12254 19343 12310 19352
rect 12164 18896 12216 18902
rect 12164 18838 12216 18844
rect 11980 18760 12032 18766
rect 12176 18737 12204 18838
rect 12256 18760 12308 18766
rect 11980 18702 12032 18708
rect 12162 18728 12218 18737
rect 12308 18720 12388 18748
rect 12256 18702 12308 18708
rect 12162 18663 12218 18672
rect 11808 18006 11928 18034
rect 12070 18048 12126 18057
rect 11808 17202 11836 18006
rect 12070 17983 12126 17992
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11900 17241 11928 17818
rect 11886 17232 11942 17241
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11796 17196 11848 17202
rect 11886 17167 11942 17176
rect 11796 17138 11848 17144
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11348 16590 11376 16934
rect 11440 16590 11468 17138
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11336 15564 11388 15570
rect 11532 15552 11560 15982
rect 11716 15609 11744 16458
rect 11388 15524 11560 15552
rect 11702 15600 11758 15609
rect 11702 15535 11758 15544
rect 11336 15506 11388 15512
rect 11702 15464 11758 15473
rect 11702 15399 11758 15408
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11532 14618 11560 15030
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11716 14464 11744 15399
rect 11808 14657 11836 17138
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16182 11928 16934
rect 12084 16674 12112 17983
rect 12162 17504 12218 17513
rect 12162 17439 12218 17448
rect 12176 17270 12204 17439
rect 12254 17368 12310 17377
rect 12254 17303 12256 17312
rect 12308 17303 12310 17312
rect 12256 17274 12308 17280
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12360 17134 12388 18720
rect 12452 18057 12480 22494
rect 12636 19394 12664 22520
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12636 19366 12848 19394
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 19145 12572 19246
rect 12820 19174 12848 19366
rect 12808 19168 12860 19174
rect 12530 19136 12586 19145
rect 12808 19110 12860 19116
rect 12530 19071 12586 19080
rect 12438 18048 12494 18057
rect 12438 17983 12494 17992
rect 12544 17678 12572 19071
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12714 18592 12770 18601
rect 12714 18527 12770 18536
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12636 17882 12664 18090
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12728 17762 12756 18527
rect 12820 18426 12848 18770
rect 13004 18426 13032 20198
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12806 17912 12862 17921
rect 12806 17847 12862 17856
rect 12636 17734 12756 17762
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 11992 16646 12112 16674
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11794 14648 11850 14657
rect 11794 14583 11850 14592
rect 11716 14436 11836 14464
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11426 13832 11482 13841
rect 11426 13767 11428 13776
rect 11480 13767 11482 13776
rect 11428 13738 11480 13744
rect 11426 13696 11482 13705
rect 11426 13631 11482 13640
rect 11440 13462 11468 13631
rect 11428 13456 11480 13462
rect 11520 13456 11572 13462
rect 11428 13398 11480 13404
rect 11518 13424 11520 13433
rect 11572 13424 11574 13433
rect 11440 13326 11468 13398
rect 11518 13359 11574 13368
rect 11716 13326 11744 14282
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11242 12336 11298 12345
rect 11152 12300 11204 12306
rect 11242 12271 11298 12280
rect 11152 12242 11204 12248
rect 10980 10798 11100 10826
rect 10980 10169 11008 10798
rect 11164 10266 11192 12242
rect 11256 10606 11284 12271
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11898 11744 12922
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11808 11744 11836 14436
rect 11886 14240 11942 14249
rect 11886 14175 11942 14184
rect 11900 12782 11928 14175
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11992 12646 12020 16646
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12084 13530 12112 16526
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12268 15570 12296 16458
rect 12360 16046 12388 17070
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12268 15434 12296 15506
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12268 15162 12296 15370
rect 12452 15162 12480 16662
rect 12636 15706 12664 17734
rect 12820 17066 12848 17847
rect 12898 17640 12954 17649
rect 12898 17575 12954 17584
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12728 16096 12756 16186
rect 12728 16068 12848 16096
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12622 15600 12678 15609
rect 12622 15535 12678 15544
rect 12636 15502 12664 15535
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12728 15366 12756 15914
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 14385 12204 14418
rect 12452 14414 12480 14962
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12256 14408 12308 14414
rect 12162 14376 12218 14385
rect 12256 14350 12308 14356
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12162 14311 12218 14320
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11980 12640 12032 12646
rect 11886 12608 11942 12617
rect 11980 12582 12032 12588
rect 11886 12543 11942 12552
rect 11716 11716 11836 11744
rect 11336 11688 11388 11694
rect 11334 11656 11336 11665
rect 11388 11656 11390 11665
rect 11334 11591 11390 11600
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11532 11354 11560 11494
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11624 11257 11652 11494
rect 11610 11248 11666 11257
rect 11610 11183 11666 11192
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11612 10736 11664 10742
rect 11334 10704 11390 10713
rect 11612 10678 11664 10684
rect 11334 10639 11390 10648
rect 11348 10606 11376 10639
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11624 10441 11652 10678
rect 11716 10470 11744 11716
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11808 11082 11836 11562
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11704 10464 11756 10470
rect 11610 10432 11666 10441
rect 11704 10406 11756 10412
rect 11610 10367 11666 10376
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11808 10198 11836 10746
rect 11244 10192 11296 10198
rect 10966 10160 11022 10169
rect 10966 10095 11022 10104
rect 11150 10160 11206 10169
rect 11244 10134 11296 10140
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11150 10095 11206 10104
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10980 9353 11008 9590
rect 10966 9344 11022 9353
rect 10966 9279 11022 9288
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10782 6216 10838 6225
rect 10782 6151 10838 6160
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10598 5400 10654 5409
rect 10598 5335 10654 5344
rect 10612 4865 10640 5335
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10598 4856 10654 4865
rect 10704 4826 10732 4966
rect 10598 4791 10654 4800
rect 10692 4820 10744 4826
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3670 10548 3878
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10428 3488 10548 3516
rect 10060 1142 10364 1170
rect 10060 480 10088 1142
rect 10520 480 10548 3488
rect 10612 2122 10640 4791
rect 10692 4762 10744 4768
rect 10796 2582 10824 6054
rect 10888 4078 10916 7686
rect 10980 4758 11008 8978
rect 11072 5166 11100 9046
rect 11164 8294 11192 10095
rect 11256 8906 11284 10134
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 9110 11560 9522
rect 11716 9489 11744 9930
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 11808 9217 11836 9862
rect 11900 9518 11928 12543
rect 11992 11937 12020 12582
rect 11978 11928 12034 11937
rect 11978 11863 12034 11872
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11992 11286 12020 11766
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11978 11112 12034 11121
rect 11978 11047 12034 11056
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11886 9344 11942 9353
rect 11886 9279 11942 9288
rect 11794 9208 11850 9217
rect 11900 9178 11928 9279
rect 11794 9143 11850 9152
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11348 8401 11376 8434
rect 11334 8392 11390 8401
rect 11334 8327 11390 8336
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7868 11284 8230
rect 11164 7840 11284 7868
rect 11164 5914 11192 7840
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 6254 11284 7686
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11716 6746 11744 8298
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11808 7206 11836 7822
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11808 6866 11836 7142
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11716 6718 11836 6746
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11612 6316 11664 6322
rect 11716 6304 11744 6598
rect 11664 6276 11744 6304
rect 11612 6258 11664 6264
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11256 4842 11284 6054
rect 11624 5846 11652 6258
rect 11808 6236 11836 6718
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11716 6208 11836 6236
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11334 5264 11390 5273
rect 11334 5199 11390 5208
rect 11348 5030 11376 5199
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11256 4814 11376 4842
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11348 4690 11376 4814
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3738 10916 3878
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10874 2680 10930 2689
rect 10874 2615 10876 2624
rect 10928 2615 10930 2624
rect 10876 2586 10928 2592
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 11072 2310 11100 4626
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4146 11192 4558
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 3398 11192 4082
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 2854 11192 3334
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11256 2650 11284 3878
rect 11716 3398 11744 6208
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5778 11836 6054
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5302 11836 5510
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11808 4146 11836 5102
rect 11900 4146 11928 6666
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11900 3738 11928 3946
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11992 2938 12020 11047
rect 12084 5953 12112 12922
rect 12176 12918 12204 14311
rect 12268 13530 12296 14350
rect 12544 14006 12572 14758
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12636 13938 12664 14894
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12728 14006 12756 14554
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12360 12322 12388 13806
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12986 12664 13330
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12268 12294 12388 12322
rect 12176 11762 12204 12242
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12176 11354 12204 11562
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10849 12204 10950
rect 12162 10840 12218 10849
rect 12162 10775 12218 10784
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12176 10130 12204 10678
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12176 8974 12204 10066
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 7750 12204 8910
rect 12268 8634 12296 12294
rect 12346 12064 12402 12073
rect 12346 11999 12402 12008
rect 12360 11694 12388 11999
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12346 11520 12402 11529
rect 12346 11455 12402 11464
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12162 7440 12218 7449
rect 12162 7375 12218 7384
rect 12176 7041 12204 7375
rect 12268 7177 12296 7482
rect 12254 7168 12310 7177
rect 12254 7103 12310 7112
rect 12162 7032 12218 7041
rect 12162 6967 12218 6976
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12070 5944 12126 5953
rect 12070 5879 12126 5888
rect 12070 5672 12126 5681
rect 12070 5607 12072 5616
rect 12124 5607 12126 5616
rect 12072 5578 12124 5584
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12084 3534 12112 5170
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12084 3194 12112 3470
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11716 2910 12020 2938
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11624 2582 11652 2858
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 11150 2408 11206 2417
rect 11150 2343 11206 2352
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 10612 2094 11008 2122
rect 10980 480 11008 2094
rect 11164 1834 11192 2343
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11152 1828 11204 1834
rect 11152 1770 11204 1776
rect 11716 1442 11744 2910
rect 11886 2816 11942 2825
rect 11886 2751 11942 2760
rect 11440 1414 11744 1442
rect 11440 480 11468 1414
rect 11900 480 11928 2751
rect 12084 2446 12112 3130
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12176 2038 12204 6054
rect 12254 3632 12310 3641
rect 12254 3567 12310 3576
rect 12268 2961 12296 3567
rect 12254 2952 12310 2961
rect 12254 2887 12310 2896
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 12360 480 12388 11455
rect 12452 11354 12480 12582
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12544 11218 12572 12718
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12452 9654 12480 11086
rect 12636 10674 12664 12242
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11150 12756 11630
rect 12820 11354 12848 16068
rect 12912 12918 12940 17575
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 13802 13032 16390
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12900 12912 12952 12918
rect 12898 12880 12900 12889
rect 12952 12880 12954 12889
rect 12898 12815 12954 12824
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12820 10674 12848 11154
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12530 10296 12586 10305
rect 12530 10231 12586 10240
rect 12544 9761 12572 10231
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12636 9518 12664 9862
rect 12728 9722 12756 10406
rect 12912 10266 12940 12582
rect 13004 12374 13032 12786
rect 12992 12368 13044 12374
rect 12992 12310 13044 12316
rect 13004 11506 13032 12310
rect 13096 12170 13124 22520
rect 13556 20806 13584 22520
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13372 19718 13400 20402
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13372 19145 13400 19654
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13452 19168 13504 19174
rect 13358 19136 13414 19145
rect 13452 19110 13504 19116
rect 13358 19071 13414 19080
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17882 13400 18022
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13188 12764 13216 17750
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 15978 13400 16390
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13280 14006 13308 15506
rect 13372 15162 13400 15914
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13372 14113 13400 14418
rect 13358 14104 13414 14113
rect 13358 14039 13414 14048
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13268 13864 13320 13870
rect 13360 13864 13412 13870
rect 13268 13806 13320 13812
rect 13358 13832 13360 13841
rect 13412 13832 13414 13841
rect 13280 12918 13308 13806
rect 13358 13767 13414 13776
rect 13372 13326 13400 13767
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13188 12736 13308 12764
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13004 11478 13124 11506
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12440 9104 12492 9110
rect 12492 9064 12572 9092
rect 12440 9046 12492 9052
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6254 12480 7142
rect 12544 6866 12572 9064
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 7342 12756 7686
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12530 5944 12586 5953
rect 12530 5879 12586 5888
rect 12544 5794 12572 5879
rect 12452 5778 12572 5794
rect 12440 5772 12572 5778
rect 12492 5766 12572 5772
rect 12440 5714 12492 5720
rect 12636 5681 12664 7142
rect 12728 6254 12756 7278
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12622 5672 12678 5681
rect 12622 5607 12678 5616
rect 12440 5568 12492 5574
rect 12728 5556 12756 6190
rect 12440 5510 12492 5516
rect 12544 5528 12756 5556
rect 12452 2514 12480 5510
rect 12544 4622 12572 5528
rect 12624 5024 12676 5030
rect 12820 4978 12848 8298
rect 12624 4966 12676 4972
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12544 3534 12572 4558
rect 12636 3913 12664 4966
rect 12728 4950 12848 4978
rect 12728 4049 12756 4950
rect 12806 4720 12862 4729
rect 12806 4655 12862 4664
rect 12820 4185 12848 4655
rect 12806 4176 12862 4185
rect 12806 4111 12862 4120
rect 12714 4040 12770 4049
rect 12714 3975 12770 3984
rect 12716 3936 12768 3942
rect 12622 3904 12678 3913
rect 12716 3878 12768 3884
rect 12622 3839 12678 3848
rect 12728 3670 12756 3878
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12636 2378 12664 3538
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12820 2990 12848 3470
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12912 2836 12940 9114
rect 12820 2808 12940 2836
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12820 480 12848 2808
rect 13004 2650 13032 9998
rect 13096 9586 13124 11478
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13188 9518 13216 10474
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13096 9042 13124 9114
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13082 6352 13138 6361
rect 13082 6287 13138 6296
rect 13096 5778 13124 6287
rect 13188 5794 13216 8026
rect 13280 7857 13308 12736
rect 13464 12617 13492 19110
rect 13832 18902 13860 19450
rect 13924 18970 13952 20266
rect 14004 19712 14056 19718
rect 14002 19680 14004 19689
rect 14056 19680 14058 19689
rect 14002 19615 14058 19624
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13820 18896 13872 18902
rect 14004 18896 14056 18902
rect 13820 18838 13872 18844
rect 13910 18864 13966 18873
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13556 17134 13584 18702
rect 13832 18290 13860 18838
rect 14004 18838 14056 18844
rect 13910 18799 13966 18808
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13832 17882 13860 18090
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13648 15473 13676 17682
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 17241 13860 17614
rect 13818 17232 13874 17241
rect 13818 17167 13874 17176
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16454 13860 17070
rect 13924 16998 13952 18799
rect 14016 18737 14044 18838
rect 14002 18728 14058 18737
rect 14002 18663 14058 18672
rect 14108 18630 14136 22520
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14200 18290 14228 19926
rect 14292 19242 14320 20470
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14476 19417 14504 19722
rect 14462 19408 14518 19417
rect 14462 19343 14518 19352
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14384 18970 14412 19110
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14016 17649 14044 18226
rect 14292 18170 14320 18566
rect 14200 18142 14320 18170
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14002 17640 14058 17649
rect 14002 17575 14058 17584
rect 14002 17096 14058 17105
rect 14002 17031 14058 17040
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 14016 16726 14044 17031
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13924 16250 13952 16594
rect 14108 16250 14136 17682
rect 14200 16833 14228 18142
rect 14186 16824 14242 16833
rect 14186 16759 14242 16768
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14200 16130 14228 16390
rect 14108 16102 14228 16130
rect 13634 15464 13690 15473
rect 13634 15399 13690 15408
rect 13648 14634 13676 15399
rect 14108 15162 14136 16102
rect 14292 15638 14320 16730
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 14384 15434 14412 18770
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14476 15337 14504 19343
rect 14568 18426 14596 22520
rect 15028 20602 15056 22520
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14568 16114 14596 16730
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14660 15609 14688 20334
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14752 19310 14780 19994
rect 14740 19304 14792 19310
rect 15212 19281 15240 20334
rect 15488 20058 15516 22520
rect 15948 20602 15976 22520
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15396 19310 15424 19858
rect 15384 19304 15436 19310
rect 14740 19246 14792 19252
rect 15198 19272 15254 19281
rect 15384 19246 15436 19252
rect 15198 19207 15254 19216
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14844 18193 14872 18362
rect 14830 18184 14886 18193
rect 14830 18119 14886 18128
rect 15198 18048 15254 18057
rect 14817 17980 15113 18000
rect 15198 17983 15254 17992
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16522 14780 17002
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14752 16114 14780 16458
rect 15212 16454 15240 17983
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14646 15600 14702 15609
rect 14646 15535 14702 15544
rect 15212 15366 15240 15982
rect 15200 15360 15252 15366
rect 14462 15328 14518 15337
rect 15200 15302 15252 15308
rect 14462 15263 14518 15272
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13556 14606 13676 14634
rect 13450 12608 13506 12617
rect 13450 12543 13506 12552
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13372 9081 13400 12106
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 11694 13492 12038
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13556 10130 13584 14606
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13648 13462 13676 14486
rect 13740 14074 13768 14894
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14346 13952 14758
rect 14292 14550 14320 15098
rect 15304 15042 15332 18838
rect 15396 15162 15424 18906
rect 15580 18698 15608 19858
rect 16304 19372 16356 19378
rect 16304 19314 16356 19320
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 17338 15884 17614
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15488 16046 15516 17274
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15580 16402 15608 16730
rect 15672 16590 15700 17138
rect 16040 16794 16068 19178
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15856 16674 15884 16730
rect 15764 16646 15884 16674
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15660 16448 15712 16454
rect 15580 16396 15660 16402
rect 15580 16390 15712 16396
rect 15580 16374 15700 16390
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 14648 15020 14700 15026
rect 15304 15014 15424 15042
rect 14648 14962 14700 14968
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14292 14385 14320 14486
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14278 14376 14334 14385
rect 13912 14340 13964 14346
rect 14278 14311 14334 14320
rect 13912 14282 13964 14288
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13832 12782 13860 14214
rect 13924 13161 13952 14282
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13910 13152 13966 13161
rect 13910 13087 13966 13096
rect 14016 12850 14044 14214
rect 14278 14104 14334 14113
rect 14278 14039 14334 14048
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13910 12608 13966 12617
rect 13648 12442 13676 12582
rect 14200 12594 14228 13738
rect 14292 12714 14320 14039
rect 14384 13705 14412 14418
rect 14370 13696 14426 13705
rect 14370 13631 14426 13640
rect 14384 13025 14412 13631
rect 14370 13016 14426 13025
rect 14476 12986 14504 14758
rect 14568 14278 14596 14758
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14556 14000 14608 14006
rect 14660 13988 14688 14962
rect 15292 14952 15344 14958
rect 15106 14920 15162 14929
rect 15292 14894 15344 14900
rect 15106 14855 15108 14864
rect 15160 14855 15162 14864
rect 15108 14826 15160 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14608 13960 14688 13988
rect 14556 13942 14608 13948
rect 14370 12951 14426 12960
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14464 12776 14516 12782
rect 14370 12744 14426 12753
rect 14280 12708 14332 12714
rect 14464 12718 14516 12724
rect 14370 12679 14426 12688
rect 14280 12650 14332 12656
rect 14200 12566 14320 12594
rect 13910 12543 13966 12552
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13818 11248 13874 11257
rect 13818 11183 13874 11192
rect 13832 10470 13860 11183
rect 13924 11014 13952 12543
rect 14094 12200 14150 12209
rect 14094 12135 14150 12144
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13820 10464 13872 10470
rect 13634 10432 13690 10441
rect 13820 10406 13872 10412
rect 13634 10367 13690 10376
rect 13648 10266 13676 10367
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13832 10146 13860 10406
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13648 10118 13860 10146
rect 13358 9072 13414 9081
rect 13358 9007 13414 9016
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13266 7848 13322 7857
rect 13266 7783 13322 7792
rect 13084 5772 13136 5778
rect 13188 5766 13308 5794
rect 13084 5714 13136 5720
rect 13096 5302 13124 5714
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4078 13124 4966
rect 13188 4078 13216 5646
rect 13280 4321 13308 5766
rect 13372 5098 13400 8910
rect 13452 7472 13504 7478
rect 13556 7460 13584 10066
rect 13648 9110 13676 10118
rect 13924 10010 13952 10950
rect 13832 9982 13952 10010
rect 13832 9738 13860 9982
rect 13740 9710 13860 9738
rect 13740 9364 13768 9710
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13832 9518 13860 9590
rect 14016 9586 14044 11154
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13820 9376 13872 9382
rect 13740 9336 13820 9364
rect 13820 9318 13872 9324
rect 13636 9104 13688 9110
rect 13832 9081 13860 9318
rect 13636 9046 13688 9052
rect 13818 9072 13874 9081
rect 13818 9007 13874 9016
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13740 7954 13768 8842
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13504 7432 13584 7460
rect 13452 7414 13504 7420
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13740 6225 13768 6938
rect 13726 6216 13782 6225
rect 13726 6151 13782 6160
rect 13832 5846 13860 8774
rect 14016 8498 14044 9522
rect 14108 8634 14136 12135
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14200 11665 14228 11766
rect 14186 11656 14242 11665
rect 14186 11591 14242 11600
rect 14200 11218 14228 11591
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10198 14228 10950
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14186 10024 14242 10033
rect 14186 9959 14242 9968
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14108 8430 14136 8570
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 13924 6798 13952 8230
rect 14108 8090 14136 8230
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7290 14136 7686
rect 14016 7274 14136 7290
rect 14004 7268 14136 7274
rect 14056 7262 14136 7268
rect 14004 7210 14056 7216
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 5840 13872 5846
rect 13818 5808 13820 5817
rect 13872 5808 13874 5817
rect 14016 5778 14044 7210
rect 13818 5743 13874 5752
rect 14004 5772 14056 5778
rect 14056 5732 14136 5760
rect 14004 5714 14056 5720
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 13266 4312 13322 4321
rect 13266 4247 13322 4256
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13082 3904 13138 3913
rect 13082 3839 13138 3848
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12912 2038 12940 2382
rect 12900 2032 12952 2038
rect 12900 1974 12952 1980
rect 13004 1970 13032 2586
rect 12992 1964 13044 1970
rect 12992 1906 13044 1912
rect 13096 610 13124 3839
rect 13188 3738 13216 4014
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 2802 13216 3334
rect 13280 2922 13308 3674
rect 13372 3210 13400 5034
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13464 4282 13492 4762
rect 13556 4729 13584 5170
rect 13542 4720 13598 4729
rect 13542 4655 13598 4664
rect 13648 4486 13676 5170
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13556 3398 13584 4422
rect 13648 4214 13676 4422
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13648 3602 13676 4150
rect 13740 3738 13768 4218
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13832 3534 13860 4966
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13372 3182 13768 3210
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13188 2774 13308 2802
rect 13084 604 13136 610
rect 13084 546 13136 552
rect 13280 480 13308 2774
rect 13740 480 13768 3182
rect 13924 2106 13952 4626
rect 14108 4554 14136 5732
rect 14200 5681 14228 9959
rect 14292 9625 14320 12566
rect 14384 12374 14412 12679
rect 14476 12481 14504 12718
rect 14462 12472 14518 12481
rect 14462 12407 14518 12416
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14384 10674 14412 12174
rect 14568 11694 14596 13942
rect 14752 13870 14780 14758
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14844 13870 14872 14486
rect 15304 14328 15332 14894
rect 15396 14396 15424 15014
rect 15488 14958 15516 15302
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14550 15516 14894
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15396 14368 15516 14396
rect 15304 14300 15424 14328
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 14740 13864 14792 13870
rect 14832 13864 14884 13870
rect 14740 13806 14792 13812
rect 14830 13832 14832 13841
rect 14884 13832 14886 13841
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13326 14688 13738
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14752 13258 14780 13806
rect 14830 13767 14886 13776
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14462 11112 14518 11121
rect 14462 11047 14464 11056
rect 14516 11047 14518 11056
rect 14464 11018 14516 11024
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 10062 14412 10610
rect 14476 10606 14504 11018
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14568 10452 14596 11154
rect 14476 10424 14596 10452
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14370 9752 14426 9761
rect 14370 9687 14426 9696
rect 14278 9616 14334 9625
rect 14278 9551 14334 9560
rect 14292 5846 14320 9551
rect 14384 8362 14412 9687
rect 14476 9654 14504 10424
rect 14660 9654 14688 12854
rect 14752 12850 14780 13194
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14844 12628 14872 13262
rect 14752 12600 14872 12628
rect 14464 9648 14516 9654
rect 14648 9648 14700 9654
rect 14464 9590 14516 9596
rect 14554 9616 14610 9625
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 14186 5672 14242 5681
rect 14186 5607 14242 5616
rect 14200 5030 14228 5607
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14188 4480 14240 4486
rect 14108 4428 14188 4434
rect 14108 4422 14240 4428
rect 14108 4406 14228 4422
rect 14108 4146 14136 4406
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3194 14136 3878
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14200 2854 14228 4218
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14292 3641 14320 3674
rect 14278 3632 14334 3641
rect 14278 3567 14334 3576
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14002 2680 14058 2689
rect 14002 2615 14004 2624
rect 14056 2615 14058 2624
rect 14004 2586 14056 2592
rect 14002 2544 14058 2553
rect 14002 2479 14004 2488
rect 14056 2479 14058 2488
rect 14004 2450 14056 2456
rect 14200 2446 14228 2790
rect 14384 2582 14412 7890
rect 14476 7410 14504 9590
rect 14752 9625 14780 12600
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15212 12306 15240 14010
rect 15396 13977 15424 14300
rect 15382 13968 15438 13977
rect 15382 13903 15438 13912
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12986 15332 13262
rect 15396 13258 15424 13903
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14922 10024 14978 10033
rect 14922 9959 14978 9968
rect 14648 9590 14700 9596
rect 14738 9616 14794 9625
rect 14554 9551 14610 9560
rect 14738 9551 14794 9560
rect 14568 9518 14596 9551
rect 14556 9512 14608 9518
rect 14936 9466 14964 9959
rect 14556 9454 14608 9460
rect 14660 9438 14964 9466
rect 14660 9364 14688 9438
rect 14568 9353 14688 9364
rect 14554 9344 14688 9353
rect 14610 9336 14688 9344
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14554 9279 14610 9288
rect 14568 7834 14596 9279
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14752 8344 14780 9318
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15212 9178 15240 9318
rect 15304 9217 15332 12310
rect 15396 11132 15424 12582
rect 15488 12186 15516 14368
rect 15580 12374 15608 16374
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15672 13530 15700 14486
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15488 12158 15608 12186
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15488 11898 15516 12038
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15396 11104 15516 11132
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15396 10130 15424 10610
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15290 9208 15346 9217
rect 15200 9172 15252 9178
rect 15290 9143 15346 9152
rect 15200 9114 15252 9120
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15014 8528 15070 8537
rect 15120 8498 15148 8774
rect 15014 8463 15016 8472
rect 15068 8463 15070 8472
rect 15108 8492 15160 8498
rect 15016 8434 15068 8440
rect 15108 8434 15160 8440
rect 15108 8356 15160 8362
rect 14752 8316 15108 8344
rect 14660 7954 14688 8298
rect 14752 8022 14780 8316
rect 15108 8298 15160 8304
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14568 7806 14688 7834
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 3126 14504 7142
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14372 2576 14424 2582
rect 14372 2518 14424 2524
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 13912 2100 13964 2106
rect 13912 2042 13964 2048
rect 14096 604 14148 610
rect 14096 546 14148 552
rect 14108 480 14136 546
rect 14568 480 14596 7686
rect 14660 5778 14688 7806
rect 15212 7342 15240 8910
rect 15304 8430 15332 8978
rect 15396 8838 15424 10066
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15382 8528 15438 8537
rect 15382 8463 15438 8472
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15396 8072 15424 8463
rect 15304 8044 15424 8072
rect 15304 7954 15332 8044
rect 15488 7993 15516 11104
rect 15474 7984 15530 7993
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15384 7948 15436 7954
rect 15474 7919 15530 7928
rect 15384 7890 15436 7896
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 6254 14780 7142
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15396 6798 15424 7890
rect 15580 7342 15608 12158
rect 15672 10554 15700 13194
rect 15764 12730 15792 16646
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16040 16425 16068 16458
rect 16026 16416 16082 16425
rect 16026 16351 16082 16360
rect 15844 15496 15896 15502
rect 15896 15456 16068 15484
rect 15844 15438 15896 15444
rect 15844 14544 15896 14550
rect 15896 14504 15976 14532
rect 15844 14486 15896 14492
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14074 15884 14350
rect 15948 14346 15976 14504
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15856 13258 15884 14010
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15948 12850 15976 13806
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15764 12702 15976 12730
rect 15948 11642 15976 12702
rect 16040 11762 16068 15456
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15948 11614 16068 11642
rect 15752 11552 15804 11558
rect 15936 11552 15988 11558
rect 15804 11512 15884 11540
rect 15752 11494 15804 11500
rect 15856 11150 15884 11512
rect 15936 11494 15988 11500
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10674 15884 11086
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15948 10606 15976 11494
rect 15936 10600 15988 10606
rect 15672 10526 15884 10554
rect 15936 10542 15988 10548
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 8430 15700 10406
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15764 9722 15792 10134
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15764 8537 15792 9658
rect 15750 8528 15806 8537
rect 15750 8463 15806 8472
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15750 8256 15806 8265
rect 15750 8191 15806 8200
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15568 7336 15620 7342
rect 15566 7304 15568 7313
rect 15620 7304 15622 7313
rect 15566 7239 15622 7248
rect 15384 6792 15436 6798
rect 15672 6769 15700 8026
rect 15764 8022 15792 8191
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15856 7426 15884 10526
rect 15936 10464 15988 10470
rect 15934 10432 15936 10441
rect 15988 10432 15990 10441
rect 15934 10367 15990 10376
rect 15948 8401 15976 10367
rect 16040 9382 16068 11614
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16132 8906 16160 19246
rect 16316 17762 16344 19314
rect 16224 17734 16344 17762
rect 16224 15745 16252 17734
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16316 16794 16344 17614
rect 16408 17377 16436 20334
rect 16500 19174 16528 22520
rect 16960 20602 16988 22520
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17420 20058 17448 22520
rect 17880 20058 17908 22520
rect 17958 21176 18014 21185
rect 17958 21111 18014 21120
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16592 19310 16620 19858
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16684 18601 16712 19246
rect 16670 18592 16726 18601
rect 16670 18527 16726 18536
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17814 16620 18022
rect 16580 17808 16632 17814
rect 16580 17750 16632 17756
rect 16684 17762 16712 18226
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17882 16804 18022
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16684 17734 16804 17762
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16394 17368 16450 17377
rect 16592 17338 16620 17614
rect 16394 17303 16450 17312
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16408 16114 16436 17138
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16592 16794 16620 16934
rect 16776 16810 16804 17734
rect 16948 17128 17000 17134
rect 16946 17096 16948 17105
rect 17000 17096 17002 17105
rect 16946 17031 17002 17040
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16684 16782 16804 16810
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15994 16436 16050
rect 16316 15966 16436 15994
rect 16210 15736 16266 15745
rect 16210 15671 16266 15680
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16224 12617 16252 15574
rect 16316 15570 16344 15966
rect 16500 15910 16528 16390
rect 16592 16046 16620 16594
rect 16684 16182 16712 16782
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16394 15736 16450 15745
rect 16394 15671 16450 15680
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 14414 16344 14758
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16316 13841 16344 13942
rect 16302 13832 16358 13841
rect 16302 13767 16358 13776
rect 16316 12850 16344 13767
rect 16408 13394 16436 15671
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 14822 16528 15302
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16486 14376 16542 14385
rect 16486 14311 16542 14320
rect 16500 13734 16528 14311
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16210 12608 16266 12617
rect 16210 12543 16266 12552
rect 16316 12374 16344 12786
rect 16408 12753 16436 13194
rect 16394 12744 16450 12753
rect 16394 12679 16450 12688
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16408 12102 16436 12242
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16302 11928 16358 11937
rect 16500 11914 16528 13670
rect 16592 13462 16620 14418
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16684 12481 16712 15846
rect 16776 15706 16804 16594
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16960 15450 16988 16118
rect 16776 15422 16988 15450
rect 16776 14362 16804 15422
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16776 14334 16896 14362
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14074 16804 14214
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16868 13682 16896 14334
rect 16960 13734 16988 14826
rect 17052 14657 17080 19926
rect 17972 19786 18000 21111
rect 18340 20890 18368 22520
rect 18156 20862 18368 20890
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 18156 19174 18184 20862
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18248 18970 18276 19246
rect 18892 19174 18920 22520
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18696 18896 18748 18902
rect 17682 18864 17738 18873
rect 18696 18838 18748 18844
rect 17682 18799 17738 18808
rect 17696 18408 17724 18799
rect 18144 18624 18196 18630
rect 18050 18592 18106 18601
rect 18144 18566 18196 18572
rect 18050 18527 18106 18536
rect 17696 18380 17908 18408
rect 17880 18329 17908 18380
rect 17866 18320 17922 18329
rect 17776 18284 17828 18290
rect 17866 18255 17922 18264
rect 17776 18226 17828 18232
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17144 16998 17172 17614
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17132 15904 17184 15910
rect 17130 15872 17132 15881
rect 17184 15872 17186 15881
rect 17130 15807 17186 15816
rect 17130 14920 17186 14929
rect 17130 14855 17186 14864
rect 17038 14648 17094 14657
rect 17038 14583 17094 14592
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17052 14249 17080 14350
rect 17038 14240 17094 14249
rect 17038 14175 17094 14184
rect 16776 13654 16896 13682
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16776 12753 16804 13654
rect 17144 13410 17172 14855
rect 16960 13382 17172 13410
rect 16762 12744 16818 12753
rect 16762 12679 16818 12688
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16670 12472 16726 12481
rect 16670 12407 16726 12416
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16302 11863 16304 11872
rect 16356 11863 16358 11872
rect 16408 11886 16528 11914
rect 16304 11834 16356 11840
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16224 9586 16252 11698
rect 16316 11694 16344 11834
rect 16408 11694 16436 11886
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16394 11384 16450 11393
rect 16394 11319 16450 11328
rect 16302 10840 16358 10849
rect 16302 10775 16358 10784
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 8974 16252 9318
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16316 8786 16344 10775
rect 16408 10690 16436 11319
rect 16500 11014 16528 11698
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10810 16528 10950
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16408 10662 16528 10690
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16408 8906 16436 9522
rect 16500 9489 16528 10662
rect 16486 9480 16542 9489
rect 16486 9415 16542 9424
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16500 9178 16528 9318
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16592 8974 16620 12310
rect 16776 11898 16804 12582
rect 16854 12200 16910 12209
rect 16854 12135 16910 12144
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16762 11792 16818 11801
rect 16762 11727 16818 11736
rect 16670 11656 16726 11665
rect 16670 11591 16672 11600
rect 16724 11591 16726 11600
rect 16672 11562 16724 11568
rect 16776 11150 16804 11727
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16684 9382 16712 11018
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9586 16804 9862
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 15934 8392 15990 8401
rect 15934 8327 15990 8336
rect 16224 8090 16252 8774
rect 16316 8758 16620 8786
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 15856 7398 16068 7426
rect 16316 7410 16344 8230
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15948 7002 15976 7142
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15384 6734 15436 6740
rect 15658 6760 15714 6769
rect 15658 6695 15714 6704
rect 15384 6656 15436 6662
rect 15660 6656 15712 6662
rect 15384 6598 15436 6604
rect 15658 6624 15660 6633
rect 15712 6624 15714 6633
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14752 5794 14780 6190
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14648 5772 14700 5778
rect 14752 5766 14872 5794
rect 14648 5714 14700 5720
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14660 4282 14688 5578
rect 14752 5166 14780 5646
rect 14844 5302 14872 5766
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14936 5012 14964 5714
rect 15212 5234 15240 6326
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14752 4984 14964 5012
rect 14752 4808 14780 4984
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14752 4780 15056 4808
rect 14922 4584 14978 4593
rect 14922 4519 14978 4528
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14738 4312 14794 4321
rect 14648 4276 14700 4282
rect 14738 4247 14794 4256
rect 14648 4218 14700 4224
rect 14752 4214 14780 4247
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14844 3924 14872 4422
rect 14936 4321 14964 4519
rect 14922 4312 14978 4321
rect 14922 4247 14978 4256
rect 14936 4010 14964 4247
rect 15028 4010 15056 4780
rect 15212 4622 15240 5170
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15120 4146 15148 4218
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15198 4040 15254 4049
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 15016 4004 15068 4010
rect 15198 3975 15200 3984
rect 15016 3946 15068 3952
rect 15252 3975 15254 3984
rect 15200 3946 15252 3952
rect 14752 3896 14872 3924
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 14660 2514 14688 3431
rect 14752 2650 14780 3896
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15304 3738 15332 5034
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 14830 3632 14886 3641
rect 14830 3567 14886 3576
rect 14844 2990 14872 3567
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 15212 2854 15240 3402
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15028 480 15056 2246
rect 15396 1442 15424 6598
rect 15658 6559 15714 6568
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15488 5778 15516 6394
rect 15566 6352 15622 6361
rect 15566 6287 15622 6296
rect 15660 6316 15712 6322
rect 15580 6254 15608 6287
rect 15660 6258 15712 6264
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15488 5030 15516 5238
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15580 4826 15608 6054
rect 15672 5846 15700 6258
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15764 5574 15792 6870
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15672 5166 15700 5510
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15672 4826 15700 5102
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15580 4706 15608 4762
rect 15580 4678 15700 4706
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15580 4214 15608 4490
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15580 3058 15608 4150
rect 15672 3738 15700 4678
rect 15752 4684 15804 4690
rect 15856 4672 15884 6938
rect 15934 6760 15990 6769
rect 15934 6695 15990 6704
rect 15948 5930 15976 6695
rect 16040 6118 16068 7398
rect 16304 7404 16356 7410
rect 16488 7404 16540 7410
rect 16304 7346 16356 7352
rect 16408 7364 16488 7392
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16132 6322 16160 6870
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15948 5902 16160 5930
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15804 4644 15884 4672
rect 15752 4626 15804 4632
rect 15856 4282 15884 4644
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15764 3194 15792 3470
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15396 1414 15516 1442
rect 15488 480 15516 1414
rect 15948 480 15976 5306
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 16040 3534 16068 5034
rect 16132 4049 16160 5902
rect 16118 4040 16174 4049
rect 16118 3975 16174 3984
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16040 3058 16068 3470
rect 16224 3466 16252 7278
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 5370 16344 6734
rect 16408 6338 16436 7364
rect 16488 7346 16540 7352
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16500 6458 16528 6870
rect 16592 6458 16620 8758
rect 16684 8634 16712 8978
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16776 8498 16804 9522
rect 16868 8974 16896 12135
rect 16960 10810 16988 13382
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17040 12980 17092 12986
rect 17144 12968 17172 13194
rect 17236 13138 17264 17614
rect 17328 16794 17356 17682
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 16794 17448 17478
rect 17592 17264 17644 17270
rect 17592 17206 17644 17212
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 13258 17356 16594
rect 17406 15056 17462 15065
rect 17406 14991 17408 15000
rect 17460 14991 17462 15000
rect 17408 14962 17460 14968
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 13938 17448 14758
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17420 13326 17448 13874
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17236 13110 17448 13138
rect 17092 12940 17172 12968
rect 17314 13016 17370 13025
rect 17314 12951 17370 12960
rect 17040 12922 17092 12928
rect 17144 12374 17172 12940
rect 17328 12850 17356 12951
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17222 12608 17278 12617
rect 17222 12543 17278 12552
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17144 10418 17172 11154
rect 17236 10538 17264 12543
rect 17328 12442 17356 12650
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17314 12200 17370 12209
rect 17314 12135 17370 12144
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 16960 10390 17172 10418
rect 16960 10062 16988 10390
rect 17328 10282 17356 12135
rect 17052 10254 17356 10282
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16960 9518 16988 9862
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 8090 16712 8230
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16684 6338 16712 6870
rect 16776 6633 16804 8298
rect 16868 7750 16896 8434
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16762 6624 16818 6633
rect 16762 6559 16818 6568
rect 16408 6310 16528 6338
rect 16500 6304 16528 6310
rect 16580 6316 16632 6322
rect 16500 6276 16580 6304
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16408 5914 16436 6190
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16500 5574 16528 6276
rect 16684 6310 16804 6338
rect 16580 6258 16632 6264
rect 16670 6080 16726 6089
rect 16670 6015 16726 6024
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16316 4758 16344 5306
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16408 4214 16436 5510
rect 16500 5166 16528 5510
rect 16684 5166 16712 6015
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16578 4992 16634 5001
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16302 3224 16358 3233
rect 16302 3159 16358 3168
rect 16316 3126 16344 3159
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16500 3058 16528 4966
rect 16578 4927 16634 4936
rect 16592 4185 16620 4927
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16040 2446 16068 2994
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16316 2650 16344 2926
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16592 2553 16620 3674
rect 16684 3602 16712 5102
rect 16776 3670 16804 6310
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16578 2544 16634 2553
rect 16578 2479 16634 2488
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16776 1766 16804 2382
rect 16764 1760 16816 1766
rect 16764 1702 16816 1708
rect 16396 1284 16448 1290
rect 16396 1226 16448 1232
rect 16408 480 16436 1226
rect 16868 480 16896 7414
rect 16960 4146 16988 8842
rect 17052 8498 17080 10254
rect 17420 10146 17448 13110
rect 17512 12481 17540 17002
rect 17604 16590 17632 17206
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17604 12918 17632 16526
rect 17696 12986 17724 17614
rect 17788 15910 17816 18226
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17866 17368 17922 17377
rect 17866 17303 17922 17312
rect 17880 16726 17908 17303
rect 17972 17105 18000 18158
rect 17958 17096 18014 17105
rect 18064 17066 18092 18527
rect 18156 18358 18184 18566
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18326 18320 18382 18329
rect 18326 18255 18328 18264
rect 18380 18255 18382 18264
rect 18328 18226 18380 18232
rect 18708 18222 18736 18838
rect 19064 18284 19116 18290
rect 18984 18244 19064 18272
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18144 18148 18196 18154
rect 18144 18090 18196 18096
rect 17958 17031 18014 17040
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17972 16590 18000 16934
rect 18156 16794 18184 18090
rect 18418 17912 18474 17921
rect 18418 17847 18474 17856
rect 18432 17610 18460 17847
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18420 17604 18472 17610
rect 18420 17546 18472 17552
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18604 17128 18656 17134
rect 18708 17105 18736 17614
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18800 17241 18828 17274
rect 18786 17232 18842 17241
rect 18786 17167 18842 17176
rect 18604 17070 18656 17076
rect 18694 17096 18750 17105
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18616 16590 18644 17070
rect 18694 17031 18750 17040
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17972 15586 18000 16526
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18800 16153 18828 16934
rect 18786 16144 18842 16153
rect 18512 16108 18564 16114
rect 18786 16079 18842 16088
rect 18512 16050 18564 16056
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 18064 15706 18092 15846
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17972 15558 18092 15586
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17788 14958 17816 15302
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17972 15065 18000 15098
rect 17958 15056 18014 15065
rect 17958 14991 18014 15000
rect 17776 14952 17828 14958
rect 18064 14940 18092 15558
rect 17776 14894 17828 14900
rect 17972 14912 18092 14940
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 13530 17816 14214
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17498 12472 17554 12481
rect 17498 12407 17554 12416
rect 17604 11914 17632 12854
rect 17696 12374 17724 12922
rect 17866 12744 17922 12753
rect 17776 12708 17828 12714
rect 17866 12679 17922 12688
rect 17776 12650 17828 12656
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17788 12073 17816 12650
rect 17880 12442 17908 12679
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17972 12102 18000 14912
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18064 14385 18092 14418
rect 18050 14376 18106 14385
rect 18050 14311 18106 14320
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 12617 18092 13330
rect 18156 13258 18184 15914
rect 18524 15638 18552 16050
rect 18800 15706 18828 16079
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18616 14618 18644 15506
rect 18708 15473 18736 15506
rect 18694 15464 18750 15473
rect 18694 15399 18750 15408
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18616 13802 18644 14350
rect 18708 14074 18736 14826
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18602 13424 18658 13433
rect 18602 13359 18658 13368
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18524 12753 18552 12786
rect 18510 12744 18566 12753
rect 18510 12679 18566 12688
rect 18144 12640 18196 12646
rect 18050 12608 18106 12617
rect 18144 12582 18196 12588
rect 18050 12543 18106 12552
rect 17960 12096 18012 12102
rect 17774 12064 17830 12073
rect 17960 12038 18012 12044
rect 17774 11999 17830 12008
rect 17604 11886 17816 11914
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17604 11257 17632 11698
rect 17788 11286 17816 11886
rect 17972 11286 18000 12038
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17776 11280 17828 11286
rect 17590 11248 17646 11257
rect 17776 11222 17828 11228
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 17590 11183 17646 11192
rect 17604 10742 17632 11183
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17236 10118 17448 10146
rect 17236 10062 17264 10118
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17052 8090 17080 8434
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17038 6896 17094 6905
rect 17038 6831 17094 6840
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17052 3738 17080 6831
rect 17144 4321 17172 9998
rect 17236 7154 17264 9998
rect 17512 9586 17540 10542
rect 17696 10470 17724 10746
rect 17788 10470 17816 11222
rect 17958 10704 18014 10713
rect 17958 10639 18014 10648
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17696 9738 17724 10406
rect 17880 9874 17908 10474
rect 17972 9994 18000 10639
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17880 9846 18000 9874
rect 17696 9710 17908 9738
rect 17774 9616 17830 9625
rect 17500 9580 17552 9586
rect 17774 9551 17830 9560
rect 17500 9522 17552 9528
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17420 8974 17448 9454
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17406 8800 17462 8809
rect 17328 7342 17356 8774
rect 17406 8735 17462 8744
rect 17420 8090 17448 8735
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17512 7886 17540 8978
rect 17682 8664 17738 8673
rect 17682 8599 17738 8608
rect 17696 8362 17724 8599
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17788 8294 17816 9551
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17500 7880 17552 7886
rect 17406 7848 17462 7857
rect 17604 7857 17632 8230
rect 17684 7880 17736 7886
rect 17500 7822 17552 7828
rect 17590 7848 17646 7857
rect 17406 7783 17462 7792
rect 17684 7822 17736 7828
rect 17590 7783 17646 7792
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17236 7126 17356 7154
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17236 6361 17264 6666
rect 17222 6352 17278 6361
rect 17222 6287 17278 6296
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17236 5370 17264 6190
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17130 4312 17186 4321
rect 17130 4247 17186 4256
rect 17236 4146 17264 4490
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17144 3194 17172 4082
rect 17328 4078 17356 7126
rect 17420 6866 17448 7783
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7410 17632 7686
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17604 6390 17632 7346
rect 17696 6798 17724 7822
rect 17684 6792 17736 6798
rect 17880 6780 17908 9710
rect 17972 7857 18000 9846
rect 18064 8430 18092 11630
rect 18156 9178 18184 12582
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11354 18460 11494
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18524 11121 18552 11698
rect 18616 11626 18644 13359
rect 18708 13326 18736 14010
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18696 13184 18748 13190
rect 18694 13152 18696 13161
rect 18748 13152 18750 13161
rect 18694 13087 18750 13096
rect 18696 12640 18748 12646
rect 18800 12628 18828 13262
rect 18892 12782 18920 17478
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18748 12600 18828 12628
rect 18880 12640 18932 12646
rect 18696 12582 18748 12588
rect 18880 12582 18932 12588
rect 18694 11792 18750 11801
rect 18694 11727 18750 11736
rect 18708 11694 18736 11727
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18696 11552 18748 11558
rect 18694 11520 18696 11529
rect 18748 11520 18750 11529
rect 18694 11455 18750 11464
rect 18510 11112 18566 11121
rect 18510 11047 18566 11056
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18800 10674 18828 10950
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18432 10266 18460 10542
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18800 10130 18828 10610
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18800 9722 18828 10066
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18892 9602 18920 12582
rect 18708 9574 18920 9602
rect 18512 9376 18564 9382
rect 18510 9344 18512 9353
rect 18564 9344 18566 9353
rect 18510 9279 18566 9288
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18512 9104 18564 9110
rect 18510 9072 18512 9081
rect 18564 9072 18566 9081
rect 18144 9036 18196 9042
rect 18510 9007 18566 9016
rect 18144 8978 18196 8984
rect 18156 8838 18184 8978
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17958 7848 18014 7857
rect 17958 7783 18014 7792
rect 17960 7744 18012 7750
rect 18012 7692 18092 7698
rect 17960 7686 18092 7692
rect 17972 7670 18092 7686
rect 17958 7576 18014 7585
rect 17958 7511 18014 7520
rect 17972 6905 18000 7511
rect 18064 7206 18092 7670
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17958 6896 18014 6905
rect 17958 6831 18014 6840
rect 17880 6752 18000 6780
rect 17684 6734 17736 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17592 6384 17644 6390
rect 17498 6352 17554 6361
rect 17592 6326 17644 6332
rect 17498 6287 17554 6296
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17144 2666 17172 2994
rect 17052 2638 17172 2666
rect 17052 2446 17080 2638
rect 17130 2544 17186 2553
rect 17130 2479 17132 2488
rect 17184 2479 17186 2488
rect 17132 2450 17184 2456
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17144 1902 17172 2450
rect 17236 2292 17264 3334
rect 17328 3097 17356 3878
rect 17314 3088 17370 3097
rect 17314 3023 17370 3032
rect 17420 2582 17448 6190
rect 17512 5846 17540 6287
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17604 5710 17632 6326
rect 17500 5704 17552 5710
rect 17498 5672 17500 5681
rect 17592 5704 17644 5710
rect 17552 5672 17554 5681
rect 17592 5646 17644 5652
rect 17498 5607 17554 5616
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17512 3670 17540 5306
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17500 3528 17552 3534
rect 17604 3516 17632 4082
rect 17696 3602 17724 6394
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17552 3488 17632 3516
rect 17500 3470 17552 3476
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17236 2264 17356 2292
rect 17132 1896 17184 1902
rect 17132 1838 17184 1844
rect 17328 480 17356 2264
rect 17788 480 17816 6598
rect 17972 6089 18000 6752
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17958 6080 18014 6089
rect 17958 6015 18014 6024
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17880 4826 17908 5646
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17972 4457 18000 5034
rect 17958 4448 18014 4457
rect 17958 4383 18014 4392
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17880 2582 17908 4150
rect 18064 4078 18092 6598
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 18156 1306 18184 8502
rect 18326 8392 18382 8401
rect 18326 8327 18382 8336
rect 18602 8392 18658 8401
rect 18602 8327 18658 8336
rect 18340 8294 18368 8327
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18340 8090 18368 8230
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18510 7440 18566 7449
rect 18510 7375 18566 7384
rect 18524 7342 18552 7375
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18524 6866 18552 7278
rect 18616 7002 18644 8327
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18512 6860 18564 6866
rect 18564 6820 18644 6848
rect 18512 6802 18564 6808
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18616 6440 18644 6820
rect 18708 6662 18736 9574
rect 18878 9480 18934 9489
rect 18788 9444 18840 9450
rect 18878 9415 18880 9424
rect 18788 9386 18840 9392
rect 18932 9415 18934 9424
rect 18880 9386 18932 9392
rect 18800 8906 18828 9386
rect 18984 8922 19012 18244
rect 19064 18226 19116 18232
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18892 8894 19012 8922
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18800 7426 18828 8298
rect 18892 8022 18920 8894
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18892 7546 18920 7958
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18800 7398 18920 7426
rect 18892 6934 18920 7398
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18524 6412 18644 6440
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5914 18276 6054
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18524 5778 18552 6412
rect 18800 6322 18828 6802
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18512 5160 18564 5166
rect 18510 5128 18512 5137
rect 18564 5128 18566 5137
rect 18510 5063 18566 5072
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18432 4758 18460 4966
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18616 3942 18644 6122
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18248 3505 18276 3878
rect 18708 3738 18736 6054
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18800 3618 18828 6122
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18892 4554 18920 5782
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18892 4146 18920 4490
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18616 3590 18828 3618
rect 18892 3602 18920 4082
rect 18880 3596 18932 3602
rect 18234 3496 18290 3505
rect 18234 3431 18290 3440
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18418 3088 18474 3097
rect 18340 2990 18368 3062
rect 18418 3023 18420 3032
rect 18472 3023 18474 3032
rect 18512 3052 18564 3058
rect 18420 2994 18472 3000
rect 18512 2994 18564 3000
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18340 2417 18368 2926
rect 18524 2446 18552 2994
rect 18512 2440 18564 2446
rect 18326 2408 18382 2417
rect 18512 2382 18564 2388
rect 18326 2343 18382 2352
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1278 18276 1306
rect 18248 480 18276 1278
rect 18616 480 18644 3590
rect 18880 3538 18932 3544
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18708 3097 18736 3130
rect 18694 3088 18750 3097
rect 18694 3023 18750 3032
rect 18694 2816 18750 2825
rect 18694 2751 18750 2760
rect 18708 2650 18736 2751
rect 18786 2680 18842 2689
rect 18696 2644 18748 2650
rect 18786 2615 18788 2624
rect 18696 2586 18748 2592
rect 18840 2615 18842 2624
rect 18788 2586 18840 2592
rect 18984 2514 19012 8774
rect 19076 8498 19104 18022
rect 19168 17678 19196 19858
rect 19352 18970 19380 22520
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19444 18902 19472 19110
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19536 18426 19564 20334
rect 19812 20058 19840 22520
rect 19890 22128 19946 22137
rect 19890 22063 19946 22072
rect 19904 20058 19932 22063
rect 20272 20602 20300 22520
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19248 18148 19300 18154
rect 19248 18090 19300 18096
rect 19260 18057 19288 18090
rect 19246 18048 19302 18057
rect 19246 17983 19302 17992
rect 19352 17921 19380 18158
rect 19338 17912 19394 17921
rect 19338 17847 19394 17856
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19156 17264 19208 17270
rect 19154 17232 19156 17241
rect 19208 17232 19210 17241
rect 19154 17167 19210 17176
rect 19156 17128 19208 17134
rect 19154 17096 19156 17105
rect 19208 17096 19210 17105
rect 19154 17031 19210 17040
rect 19260 16658 19288 17750
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19352 16522 19380 17546
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 16017 19288 16050
rect 19340 16040 19392 16046
rect 19246 16008 19302 16017
rect 19340 15982 19392 15988
rect 19246 15943 19302 15952
rect 19260 15638 19288 15943
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 19168 15162 19196 15574
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19168 14346 19196 15098
rect 19260 14618 19288 15302
rect 19352 14618 19380 15982
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19352 13326 19380 13738
rect 19340 13320 19392 13326
rect 19246 13288 19302 13297
rect 19340 13262 19392 13268
rect 19246 13223 19302 13232
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19168 12442 19196 12786
rect 19260 12714 19288 13223
rect 19352 12850 19380 13262
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19248 12708 19300 12714
rect 19248 12650 19300 12656
rect 19444 12594 19472 16594
rect 19536 13190 19564 16662
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19522 13016 19578 13025
rect 19522 12951 19524 12960
rect 19576 12951 19578 12960
rect 19524 12922 19576 12928
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19260 12566 19472 12594
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19260 12306 19288 12566
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19260 11762 19288 12106
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19168 9518 19196 11154
rect 19260 11150 19288 11698
rect 19352 11218 19380 12242
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19260 10266 19288 10950
rect 19432 10532 19484 10538
rect 19432 10474 19484 10480
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19352 9654 19380 10134
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19260 9330 19288 9590
rect 19338 9480 19394 9489
rect 19338 9415 19394 9424
rect 19168 9302 19288 9330
rect 19168 8537 19196 9302
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19154 8528 19210 8537
rect 19064 8492 19116 8498
rect 19154 8463 19210 8472
rect 19064 8434 19116 8440
rect 19168 8072 19196 8463
rect 19076 8044 19196 8072
rect 19076 7886 19104 8044
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19076 7449 19104 7822
rect 19062 7440 19118 7449
rect 19062 7375 19118 7384
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 19076 480 19104 7142
rect 19168 2825 19196 7890
rect 19154 2816 19210 2825
rect 19154 2751 19210 2760
rect 19260 2514 19288 9114
rect 19352 9042 19380 9415
rect 19444 9178 19472 10474
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8537 19380 8978
rect 19536 8838 19564 12718
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19432 8560 19484 8566
rect 19338 8528 19394 8537
rect 19484 8520 19564 8548
rect 19432 8502 19484 8508
rect 19338 8463 19394 8472
rect 19340 8288 19392 8294
rect 19321 8236 19340 8276
rect 19321 8230 19392 8236
rect 19321 8214 19380 8230
rect 19352 8129 19380 8214
rect 19338 8120 19394 8129
rect 19338 8055 19394 8064
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19352 5914 19380 6258
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19338 5808 19394 5817
rect 19338 5743 19394 5752
rect 19352 5250 19380 5743
rect 19444 5370 19472 6054
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19352 5222 19472 5250
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19352 4690 19380 5102
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19352 610 19380 4422
rect 19444 2854 19472 5222
rect 19536 3058 19564 8520
rect 19628 6254 19656 17478
rect 19720 17338 19748 18770
rect 19812 18290 19840 19246
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19812 17218 19840 18022
rect 19904 17785 19932 18770
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19890 17776 19946 17785
rect 19890 17711 19946 17720
rect 19720 17190 19840 17218
rect 19720 16114 19748 17190
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19812 16017 19840 16934
rect 19996 16726 20024 18566
rect 20088 18086 20116 20334
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 20088 17134 20116 17750
rect 20180 17678 20208 20334
rect 20456 20058 20484 22607
rect 20718 22520 20774 23000
rect 21270 22520 21326 23000
rect 21730 22520 21786 23000
rect 22190 22520 22246 23000
rect 22650 22520 22706 23000
rect 20534 21720 20590 21729
rect 20534 21655 20590 21664
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20272 19417 20300 19858
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20258 19408 20314 19417
rect 20258 19343 20314 19352
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20272 18630 20300 19246
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 19892 16176 19944 16182
rect 19892 16118 19944 16124
rect 19798 16008 19854 16017
rect 19798 15943 19854 15952
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19720 14074 19748 15846
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19812 13530 19840 15846
rect 19904 13802 19932 16118
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19708 13456 19760 13462
rect 19706 13424 19708 13433
rect 19760 13424 19762 13433
rect 19706 13359 19762 13368
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 19720 12753 19748 13194
rect 19706 12744 19762 12753
rect 19706 12679 19762 12688
rect 19720 11694 19748 12679
rect 19812 12050 19840 13330
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19904 12986 19932 13126
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19996 12594 20024 16050
rect 20088 14521 20116 17070
rect 20180 16130 20208 17478
rect 20272 16250 20300 17818
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20180 16102 20300 16130
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 15094 20208 15438
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20272 14958 20300 16102
rect 20364 16017 20392 18566
rect 20456 17542 20484 19790
rect 20548 19174 20576 21655
rect 20626 20768 20682 20777
rect 20626 20703 20682 20712
rect 20640 20602 20668 20703
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20732 19786 20760 22520
rect 21086 20224 21142 20233
rect 21086 20159 21142 20168
rect 21100 20058 21128 20159
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20640 18290 20668 18770
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20536 17672 20588 17678
rect 20732 17649 20760 19246
rect 20824 18766 20852 19858
rect 20994 19816 21050 19825
rect 20994 19751 21050 19760
rect 21008 19514 21036 19751
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21086 19272 21142 19281
rect 21284 19242 21312 22520
rect 21086 19207 21142 19216
rect 21272 19236 21324 19242
rect 21100 18970 21128 19207
rect 21272 19178 21324 19184
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21270 18864 21326 18873
rect 21270 18799 21326 18808
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 21284 18426 21312 18799
rect 21744 18698 21772 22520
rect 22204 20534 22232 22520
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 22664 18902 22692 22520
rect 22652 18896 22704 18902
rect 22652 18838 22704 18844
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21086 18320 21142 18329
rect 21086 18255 21142 18264
rect 21100 17882 21128 18255
rect 22006 17912 22062 17921
rect 21088 17876 21140 17882
rect 22006 17847 22008 17856
rect 21088 17818 21140 17824
rect 22060 17847 22062 17856
rect 22008 17818 22060 17824
rect 21640 17808 21692 17814
rect 21640 17750 21692 17756
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20536 17614 20588 17620
rect 20718 17640 20774 17649
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20548 17202 20576 17614
rect 20718 17575 20774 17584
rect 20628 17264 20680 17270
rect 20628 17206 20680 17212
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20536 16992 20588 16998
rect 20442 16960 20498 16969
rect 20536 16934 20588 16940
rect 20442 16895 20498 16904
rect 20350 16008 20406 16017
rect 20350 15943 20406 15952
rect 20456 15706 20484 16895
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20180 14618 20208 14758
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20074 14512 20130 14521
rect 20074 14447 20130 14456
rect 20364 14414 20392 14962
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20088 12918 20116 14350
rect 20364 14006 20392 14350
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 19996 12566 20116 12594
rect 19892 12300 19944 12306
rect 19944 12260 20024 12288
rect 19892 12242 19944 12248
rect 19812 12022 19932 12050
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19720 11354 19748 11494
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19720 9625 19748 11154
rect 19706 9616 19762 9625
rect 19706 9551 19762 9560
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19720 6202 19748 9454
rect 19812 9042 19840 11834
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19812 7410 19840 8842
rect 19904 7562 19932 12022
rect 19996 9722 20024 12260
rect 20088 10606 20116 12566
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20088 10266 20116 10542
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20074 10024 20130 10033
rect 20074 9959 20130 9968
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 20088 9625 20116 9959
rect 20074 9616 20130 9625
rect 20074 9551 20130 9560
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 9217 20024 9318
rect 19982 9208 20038 9217
rect 19982 9143 20038 9152
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 20088 8378 20116 8774
rect 19996 8350 20116 8378
rect 19996 8022 20024 8350
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19984 8016 20036 8022
rect 19984 7958 20036 7964
rect 19904 7534 20024 7562
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19892 7268 19944 7274
rect 19892 7210 19944 7216
rect 19904 6730 19932 7210
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19904 6322 19932 6666
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19720 6174 19932 6202
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19616 5840 19668 5846
rect 19616 5782 19668 5788
rect 19628 5114 19656 5782
rect 19720 5234 19748 5850
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19628 5086 19748 5114
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19628 4826 19656 4966
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19720 2922 19748 5086
rect 19798 4720 19854 4729
rect 19798 4655 19800 4664
rect 19852 4655 19854 4664
rect 19800 4626 19852 4632
rect 19904 4570 19932 6174
rect 19812 4542 19932 4570
rect 19812 3942 19840 4542
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19340 604 19392 610
rect 19340 546 19392 552
rect 19536 480 19564 2858
rect 19812 2854 19840 3878
rect 19800 2848 19852 2854
rect 19904 2836 19932 4218
rect 19996 3942 20024 7534
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 20088 2990 20116 8230
rect 20180 6458 20208 13670
rect 20272 7546 20300 13806
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 20364 8514 20392 13398
rect 20456 13326 20484 13874
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20442 13016 20498 13025
rect 20442 12951 20498 12960
rect 20456 12918 20484 12951
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 11830 20484 12718
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20456 11121 20484 11494
rect 20442 11112 20498 11121
rect 20442 11047 20498 11056
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 9518 20484 9862
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20364 8486 20484 8514
rect 20350 8392 20406 8401
rect 20350 8327 20406 8336
rect 20364 8294 20392 8327
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20272 6322 20300 7346
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20166 5536 20222 5545
rect 20166 5471 20222 5480
rect 20180 5370 20208 5471
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20168 5160 20220 5166
rect 20168 5102 20220 5108
rect 20180 4146 20208 5102
rect 20272 4214 20300 6258
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20180 3534 20208 4082
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20272 3058 20300 4150
rect 20364 3602 20392 8230
rect 20456 5522 20484 8486
rect 20548 6254 20576 16934
rect 20640 16114 20668 17206
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20732 16046 20760 16730
rect 20824 16454 20852 16934
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20824 15586 20852 16390
rect 20732 15558 20852 15586
rect 20626 14512 20682 14521
rect 20732 14482 20760 15558
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20824 14958 20852 15438
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20626 14447 20682 14456
rect 20720 14476 20772 14482
rect 20640 11354 20668 14447
rect 20720 14418 20772 14424
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 20824 13394 20852 13738
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20732 11218 20760 13262
rect 20916 13190 20944 17682
rect 20994 17368 21050 17377
rect 20994 17303 21050 17312
rect 21008 15162 21036 17303
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21086 16416 21142 16425
rect 21086 16351 21142 16360
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21100 14618 21128 16351
rect 21192 15366 21220 16594
rect 21454 15464 21510 15473
rect 21454 15399 21510 15408
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21362 14104 21418 14113
rect 21362 14039 21418 14048
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20640 10305 20668 11086
rect 20824 10538 20852 12378
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20626 10296 20682 10305
rect 20626 10231 20682 10240
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20640 8634 20668 9658
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20626 8528 20682 8537
rect 20626 8463 20628 8472
rect 20680 8463 20682 8472
rect 20628 8434 20680 8440
rect 20640 7750 20668 8434
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20732 6882 20760 9318
rect 20732 6854 20852 6882
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20456 5494 20668 5522
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20534 5264 20590 5273
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19904 2808 20116 2836
rect 19800 2790 19852 2796
rect 20088 2650 20116 2808
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20364 649 20392 3538
rect 20350 640 20406 649
rect 19984 604 20036 610
rect 20350 575 20406 584
rect 19984 546 20036 552
rect 19996 480 20024 546
rect 20456 480 20484 5238
rect 20534 5199 20590 5208
rect 20548 4865 20576 5199
rect 20534 4856 20590 4865
rect 20534 4791 20590 4800
rect 20640 3126 20668 5494
rect 20732 5166 20760 6734
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20824 4146 20852 6854
rect 20916 6746 20944 12242
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21008 10606 21036 12174
rect 21100 11694 21128 12650
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 21192 11286 21220 13806
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21284 13569 21312 13670
rect 21270 13560 21326 13569
rect 21270 13495 21326 13504
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21284 10198 21312 13194
rect 21376 10810 21404 14039
rect 21468 11898 21496 15399
rect 21546 12608 21602 12617
rect 21546 12543 21602 12552
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21560 11830 21588 12543
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21008 8566 21036 9522
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 20916 6718 21036 6746
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20824 3194 20852 3878
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 1601 20668 2790
rect 20626 1592 20682 1601
rect 20626 1527 20682 1536
rect 20916 480 20944 6598
rect 21008 6390 21036 6718
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 21100 5778 21128 7142
rect 21192 6254 21220 9386
rect 21652 9178 21680 17750
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20996 5568 21048 5574
rect 21048 5528 21128 5556
rect 20996 5510 21048 5516
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21008 4622 21036 5170
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 21008 3482 21036 3946
rect 21100 3602 21128 5528
rect 21192 3670 21220 5646
rect 21284 4690 21312 9046
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 21008 3454 21128 3482
rect 21100 2922 21128 3454
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 20996 2848 21048 2854
rect 20994 2816 20996 2825
rect 21048 2816 21050 2825
rect 20994 2751 21050 2760
rect 21008 2145 21036 2751
rect 21100 2553 21128 2858
rect 21086 2544 21142 2553
rect 21086 2479 21142 2488
rect 20994 2136 21050 2145
rect 20994 2071 21050 2080
rect 21376 480 21404 5578
rect 3882 232 3938 241
rect 3882 167 3938 176
rect 4250 0 4306 480
rect 4710 0 4766 480
rect 5078 0 5134 480
rect 5538 0 5594 480
rect 5998 0 6054 480
rect 6458 0 6514 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8298 0 8354 480
rect 8758 0 8814 480
rect 9218 0 9274 480
rect 9586 0 9642 480
rect 10046 0 10102 480
rect 10506 0 10562 480
rect 10966 0 11022 480
rect 11426 0 11482 480
rect 11886 0 11942 480
rect 12346 0 12402 480
rect 12806 0 12862 480
rect 13266 0 13322 480
rect 13726 0 13782 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16394 0 16450 480
rect 16854 0 16910 480
rect 17314 0 17370 480
rect 17774 0 17830 480
rect 18234 0 18290 480
rect 18602 0 18658 480
rect 19062 0 19118 480
rect 19522 0 19578 480
rect 19982 0 20038 480
rect 20442 0 20498 480
rect 20902 0 20958 480
rect 21362 0 21418 480
rect 21468 241 21496 8230
rect 21744 8129 21772 9318
rect 21730 8120 21786 8129
rect 21730 8055 21786 8064
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21560 3058 21588 7686
rect 21548 3052 21600 3058
rect 21548 2994 21600 3000
rect 21744 1193 21772 8055
rect 21836 7342 21864 17546
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21928 7274 21956 17002
rect 22374 10160 22430 10169
rect 22374 10095 22430 10104
rect 22388 9897 22416 10095
rect 22374 9888 22430 9897
rect 22374 9823 22430 9832
rect 21916 7268 21968 7274
rect 21916 7210 21968 7216
rect 22374 6080 22430 6089
rect 22374 6015 22430 6024
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21730 1184 21786 1193
rect 21730 1119 21786 1128
rect 21836 480 21864 5510
rect 22388 4457 22416 6015
rect 22744 4480 22796 4486
rect 22374 4448 22430 4457
rect 22744 4422 22796 4428
rect 22374 4383 22430 4392
rect 22284 2304 22336 2310
rect 22284 2246 22336 2252
rect 22296 480 22324 2246
rect 22756 480 22784 4422
rect 21454 232 21510 241
rect 21454 167 21510 176
rect 21822 0 21878 480
rect 22282 0 22338 480
rect 22742 0 22798 480
<< via2 >>
rect 1858 22616 1914 22672
rect 20442 22616 20498 22672
rect 1950 21120 2006 21176
rect 1858 19760 1914 19816
rect 1950 19216 2006 19272
rect 1490 18264 1546 18320
rect 1582 17876 1638 17912
rect 1582 17856 1584 17876
rect 1584 17856 1636 17876
rect 1636 17856 1638 17876
rect 1582 17312 1638 17368
rect 1490 16904 1546 16960
rect 2318 19760 2374 19816
rect 2870 22072 2926 22128
rect 2778 20712 2834 20768
rect 2962 21664 3018 21720
rect 3054 20168 3110 20224
rect 2042 18944 2098 19000
rect 1674 16496 1730 16552
rect 1674 16360 1730 16416
rect 1950 16088 2006 16144
rect 1858 15952 1914 16008
rect 1950 15408 2006 15464
rect 1582 14456 1638 14512
rect 2778 18808 2834 18864
rect 570 3712 626 3768
rect 2502 16632 2558 16688
rect 2594 15680 2650 15736
rect 3238 18964 3294 19000
rect 3238 18944 3240 18964
rect 3240 18944 3292 18964
rect 3292 18944 3294 18964
rect 2226 12824 2282 12880
rect 3422 15816 3478 15872
rect 3882 15816 3938 15872
rect 3514 15000 3570 15056
rect 2778 14048 2834 14104
rect 1674 3440 1730 3496
rect 3238 9560 3294 9616
rect 3606 13504 3662 13560
rect 3514 12552 3570 12608
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4894 18400 4950 18456
rect 5262 18944 5318 19000
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 5814 19760 5870 19816
rect 5446 18672 5502 18728
rect 4066 16768 4122 16824
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 3422 11600 3478 11656
rect 2594 3848 2650 3904
rect 1950 3460 2006 3496
rect 1950 3440 1952 3460
rect 1952 3440 2004 3460
rect 2004 3440 2006 3460
rect 1766 3032 1822 3088
rect 2870 2760 2926 2816
rect 2778 2080 2834 2136
rect 3238 3596 3294 3632
rect 3238 3576 3240 3596
rect 3240 3576 3292 3596
rect 3292 3576 3294 3596
rect 3422 2932 3424 2952
rect 3424 2932 3476 2952
rect 3476 2932 3478 2952
rect 3422 2896 3478 2932
rect 3882 12164 3938 12200
rect 3882 12144 3884 12164
rect 3884 12144 3936 12164
rect 3936 12144 3938 12164
rect 3882 10648 3938 10704
rect 3882 10104 3938 10160
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4066 11076 4122 11112
rect 4066 11056 4068 11076
rect 4068 11056 4120 11076
rect 4120 11056 4122 11076
rect 4066 9696 4122 9752
rect 4250 8780 4252 8800
rect 4252 8780 4304 8800
rect 4304 8780 4306 8800
rect 4250 8744 4306 8780
rect 4066 8236 4068 8256
rect 4068 8236 4120 8256
rect 4120 8236 4122 8256
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4066 8200 4122 8236
rect 4066 7792 4122 7848
rect 3974 7248 4030 7304
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 3974 6296 4030 6352
rect 3974 5072 4030 5128
rect 4066 4936 4122 4992
rect 3974 4392 4030 4448
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 5814 17040 5870 17096
rect 5538 15680 5594 15736
rect 5722 12824 5778 12880
rect 5630 11872 5686 11928
rect 5722 9560 5778 9616
rect 5170 8472 5226 8528
rect 5078 7656 5134 7712
rect 5354 7948 5410 7984
rect 5354 7928 5356 7948
rect 5356 7928 5408 7948
rect 5408 7928 5410 7948
rect 4894 6296 4950 6352
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 3790 3032 3846 3088
rect 3146 2488 3202 2544
rect 3238 1536 3294 1592
rect 3146 584 3202 640
rect 4066 1128 4122 1184
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5998 16088 6054 16144
rect 5906 8744 5962 8800
rect 5814 8200 5870 8256
rect 6642 17312 6698 17368
rect 6274 11872 6330 11928
rect 6182 8608 6238 8664
rect 6182 6704 6238 6760
rect 5998 6196 6000 6216
rect 6000 6196 6052 6216
rect 6052 6196 6054 6216
rect 5998 6160 6054 6196
rect 5814 5752 5870 5808
rect 5906 4664 5962 4720
rect 5630 3304 5686 3360
rect 6182 3612 6184 3632
rect 6184 3612 6236 3632
rect 6236 3612 6238 3632
rect 6182 3576 6238 3612
rect 6274 2796 6276 2816
rect 6276 2796 6328 2816
rect 6328 2796 6330 2816
rect 6274 2760 6330 2796
rect 7102 16224 7158 16280
rect 7194 14728 7250 14784
rect 6918 13368 6974 13424
rect 6826 13232 6882 13288
rect 6734 12008 6790 12064
rect 6918 11600 6974 11656
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7654 19216 7710 19272
rect 7470 17448 7526 17504
rect 7378 17196 7434 17232
rect 7378 17176 7380 17196
rect 7380 17176 7432 17196
rect 7432 17176 7434 17196
rect 7378 16360 7434 16416
rect 7286 14184 7342 14240
rect 7378 12144 7434 12200
rect 7194 11736 7250 11792
rect 6550 8916 6552 8936
rect 6552 8916 6604 8936
rect 6604 8916 6606 8936
rect 6550 8880 6606 8916
rect 6918 9424 6974 9480
rect 6734 3168 6790 3224
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7746 17720 7802 17776
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7930 16496 7986 16552
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 8022 15272 8078 15328
rect 7838 15156 7894 15192
rect 7838 15136 7840 15156
rect 7840 15136 7892 15156
rect 7892 15136 7894 15156
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 8666 17856 8722 17912
rect 8666 16668 8668 16688
rect 8668 16668 8720 16688
rect 8720 16668 8722 16688
rect 8666 16632 8722 16668
rect 8390 15000 8446 15056
rect 8574 14592 8630 14648
rect 8482 14456 8538 14512
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7746 12280 7802 12336
rect 7654 11736 7710 11792
rect 7470 9696 7526 9752
rect 7194 8472 7250 8528
rect 7194 7812 7250 7848
rect 7194 7792 7196 7812
rect 7196 7792 7248 7812
rect 7248 7792 7250 7812
rect 7194 5208 7250 5264
rect 7378 5344 7434 5400
rect 7838 12144 7894 12200
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 8758 15272 8814 15328
rect 8942 16360 8998 16416
rect 9218 19252 9220 19272
rect 9220 19252 9272 19272
rect 9272 19252 9274 19272
rect 9218 19216 9274 19252
rect 9402 17856 9458 17912
rect 9218 16768 9274 16824
rect 8758 14456 8814 14512
rect 8758 14320 8814 14376
rect 8390 9832 8446 9888
rect 8390 9560 8446 9616
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8022 8744 8078 8800
rect 7746 8200 7802 8256
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 8298 9288 8354 9344
rect 8390 9152 8446 9208
rect 8942 14220 8944 14240
rect 8944 14220 8996 14240
rect 8996 14220 8998 14240
rect 8942 14184 8998 14220
rect 8666 9324 8668 9344
rect 8668 9324 8720 9344
rect 8720 9324 8722 9344
rect 8666 9288 8722 9324
rect 7838 7656 7894 7712
rect 7746 7248 7802 7304
rect 7470 5208 7526 5264
rect 7286 3848 7342 3904
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7930 5752 7986 5808
rect 7746 5516 7748 5536
rect 7748 5516 7800 5536
rect 7800 5516 7802 5536
rect 7746 5480 7802 5516
rect 8482 7384 8538 7440
rect 8298 5788 8300 5808
rect 8300 5788 8352 5808
rect 8352 5788 8354 5808
rect 8298 5752 8354 5788
rect 8390 5208 8446 5264
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 9586 19216 9642 19272
rect 9678 17584 9734 17640
rect 9586 16224 9642 16280
rect 9494 15988 9496 16008
rect 9496 15988 9548 16008
rect 9548 15988 9550 16008
rect 9494 15952 9550 15988
rect 10138 18536 10194 18592
rect 9770 15952 9826 16008
rect 9494 15000 9550 15056
rect 9310 14864 9366 14920
rect 9126 12144 9182 12200
rect 9126 11600 9182 11656
rect 9218 10804 9274 10840
rect 9218 10784 9220 10804
rect 9220 10784 9272 10804
rect 9272 10784 9274 10804
rect 9034 8472 9090 8528
rect 8850 7384 8906 7440
rect 9034 7656 9090 7712
rect 8942 7248 8998 7304
rect 8666 6296 8722 6352
rect 8666 6024 8722 6080
rect 8390 4936 8446 4992
rect 8574 4936 8630 4992
rect 8298 4800 8354 4856
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8574 4528 8630 4584
rect 8574 3576 8630 3632
rect 8850 5480 8906 5536
rect 9126 5480 9182 5536
rect 10138 15408 10194 15464
rect 9494 11872 9550 11928
rect 9678 11464 9734 11520
rect 9586 11228 9588 11248
rect 9588 11228 9640 11248
rect 9640 11228 9642 11248
rect 9586 11192 9642 11228
rect 9402 10376 9458 10432
rect 9402 8472 9458 8528
rect 9770 8336 9826 8392
rect 9770 8200 9826 8256
rect 9678 7520 9734 7576
rect 9770 7248 9826 7304
rect 9678 6840 9734 6896
rect 9494 6024 9550 6080
rect 9402 4936 9458 4992
rect 9954 11872 10010 11928
rect 10046 11328 10102 11384
rect 10322 17176 10378 17232
rect 10414 15680 10470 15736
rect 10322 15544 10378 15600
rect 10598 15544 10654 15600
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10414 12008 10470 12064
rect 10322 11056 10378 11112
rect 10046 8336 10102 8392
rect 10046 7656 10102 7712
rect 10046 7520 10102 7576
rect 10230 9288 10286 9344
rect 10230 5752 10286 5808
rect 10690 11872 10746 11928
rect 10506 11736 10562 11792
rect 11242 18808 11298 18864
rect 11610 19080 11666 19136
rect 11426 18944 11482 19000
rect 11610 18944 11666 19000
rect 11794 19116 11796 19136
rect 11796 19116 11848 19136
rect 11848 19116 11850 19136
rect 11794 19080 11850 19116
rect 10966 17992 11022 18048
rect 11058 17584 11114 17640
rect 10966 17448 11022 17504
rect 11150 17312 11206 17368
rect 11150 16940 11152 16960
rect 11152 16940 11204 16960
rect 11204 16940 11206 16960
rect 11150 16904 11206 16940
rect 11150 16496 11206 16552
rect 11150 15988 11152 16008
rect 11152 15988 11204 16008
rect 11204 15988 11206 16008
rect 11150 15952 11206 15988
rect 11150 15544 11206 15600
rect 11058 15136 11114 15192
rect 10782 10240 10838 10296
rect 10782 10104 10838 10160
rect 10598 8608 10654 8664
rect 10690 8472 10746 8528
rect 10506 8064 10562 8120
rect 10506 7656 10562 7712
rect 10230 4800 10286 4856
rect 9862 2508 9918 2544
rect 9862 2488 9864 2508
rect 9864 2488 9916 2508
rect 9916 2488 9918 2508
rect 10230 4392 10286 4448
rect 10322 4120 10378 4176
rect 10230 3848 10286 3904
rect 10138 3712 10194 3768
rect 10230 2624 10286 2680
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 12254 19352 12310 19408
rect 12162 18672 12218 18728
rect 12070 17992 12126 18048
rect 11886 17176 11942 17232
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11702 15544 11758 15600
rect 11702 15408 11758 15464
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 12162 17448 12218 17504
rect 12254 17332 12310 17368
rect 12254 17312 12256 17332
rect 12256 17312 12308 17332
rect 12308 17312 12310 17332
rect 12530 19080 12586 19136
rect 12438 17992 12494 18048
rect 12714 18536 12770 18592
rect 12806 17856 12862 17912
rect 11794 14592 11850 14648
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11426 13796 11482 13832
rect 11426 13776 11428 13796
rect 11428 13776 11480 13796
rect 11480 13776 11482 13796
rect 11426 13640 11482 13696
rect 11518 13404 11520 13424
rect 11520 13404 11572 13424
rect 11572 13404 11574 13424
rect 11518 13368 11574 13404
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11242 12280 11298 12336
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11886 14184 11942 14240
rect 12898 17584 12954 17640
rect 12622 15544 12678 15600
rect 12162 14320 12218 14376
rect 11886 12552 11942 12608
rect 11334 11636 11336 11656
rect 11336 11636 11388 11656
rect 11388 11636 11390 11656
rect 11334 11600 11390 11636
rect 11610 11192 11666 11248
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11334 10648 11390 10704
rect 11610 10376 11666 10432
rect 10966 10104 11022 10160
rect 11150 10104 11206 10160
rect 10966 9288 11022 9344
rect 10782 6160 10838 6216
rect 10598 5344 10654 5400
rect 10598 4800 10654 4856
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11702 9424 11758 9480
rect 11978 11872 12034 11928
rect 11978 11056 12034 11112
rect 11886 9288 11942 9344
rect 11794 9152 11850 9208
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11334 8336 11390 8392
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11334 5208 11390 5264
rect 10874 2644 10930 2680
rect 10874 2624 10876 2644
rect 10876 2624 10928 2644
rect 10928 2624 10930 2644
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12162 10784 12218 10840
rect 12346 12008 12402 12064
rect 12346 11464 12402 11520
rect 12162 7384 12218 7440
rect 12254 7112 12310 7168
rect 12162 6976 12218 7032
rect 12070 5888 12126 5944
rect 12070 5636 12126 5672
rect 12070 5616 12072 5636
rect 12072 5616 12124 5636
rect 12124 5616 12126 5636
rect 11150 2352 11206 2408
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 11886 2760 11942 2816
rect 12254 3576 12310 3632
rect 12254 2896 12310 2952
rect 12898 12860 12900 12880
rect 12900 12860 12952 12880
rect 12952 12860 12954 12880
rect 12898 12824 12954 12860
rect 12530 10240 12586 10296
rect 12530 9696 12586 9752
rect 13358 19080 13414 19136
rect 13358 14048 13414 14104
rect 13358 13812 13360 13832
rect 13360 13812 13412 13832
rect 13412 13812 13414 13832
rect 13358 13776 13414 13812
rect 12530 5888 12586 5944
rect 12622 5616 12678 5672
rect 12806 4664 12862 4720
rect 12806 4120 12862 4176
rect 12714 3984 12770 4040
rect 12622 3848 12678 3904
rect 13082 6296 13138 6352
rect 14002 19660 14004 19680
rect 14004 19660 14056 19680
rect 14056 19660 14058 19680
rect 14002 19624 14058 19660
rect 13910 18808 13966 18864
rect 13818 17176 13874 17232
rect 14002 18672 14058 18728
rect 14462 19352 14518 19408
rect 14002 17584 14058 17640
rect 14002 17040 14058 17096
rect 14186 16768 14242 16824
rect 13634 15408 13690 15464
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 15198 19216 15254 19272
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14830 18128 14886 18184
rect 15198 17992 15254 18048
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14646 15544 14702 15600
rect 14462 15272 14518 15328
rect 13450 12552 13506 12608
rect 14278 14320 14334 14376
rect 13910 13096 13966 13152
rect 14278 14048 14334 14104
rect 13910 12552 13966 12608
rect 14370 13640 14426 13696
rect 14370 12960 14426 13016
rect 15106 14884 15162 14920
rect 15106 14864 15108 14884
rect 15108 14864 15160 14884
rect 15160 14864 15162 14884
rect 14370 12688 14426 12744
rect 13818 11192 13874 11248
rect 14094 12144 14150 12200
rect 13634 10376 13690 10432
rect 13358 9016 13414 9072
rect 13266 7792 13322 7848
rect 13818 9016 13874 9072
rect 13726 6160 13782 6216
rect 14186 11600 14242 11656
rect 14186 9968 14242 10024
rect 13818 5788 13820 5808
rect 13820 5788 13872 5808
rect 13872 5788 13874 5808
rect 13818 5752 13874 5788
rect 13266 4256 13322 4312
rect 13082 3848 13138 3904
rect 13542 4664 13598 4720
rect 14462 12416 14518 12472
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14830 13812 14832 13832
rect 14832 13812 14884 13832
rect 14884 13812 14886 13832
rect 14830 13776 14886 13812
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14462 11076 14518 11112
rect 14462 11056 14464 11076
rect 14464 11056 14516 11076
rect 14516 11056 14518 11076
rect 14370 9696 14426 9752
rect 14278 9560 14334 9616
rect 14186 5616 14242 5672
rect 14278 3576 14334 3632
rect 14002 2644 14058 2680
rect 14002 2624 14004 2644
rect 14004 2624 14056 2644
rect 14056 2624 14058 2644
rect 14002 2508 14058 2544
rect 14002 2488 14004 2508
rect 14004 2488 14056 2508
rect 14056 2488 14058 2508
rect 14554 9560 14610 9616
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 15382 13912 15438 13968
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14922 9968 14978 10024
rect 14738 9560 14794 9616
rect 14554 9288 14610 9344
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 15290 9152 15346 9208
rect 15014 8492 15070 8528
rect 15014 8472 15016 8492
rect 15016 8472 15068 8492
rect 15068 8472 15070 8492
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 15382 8472 15438 8528
rect 15474 7928 15530 7984
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 16026 16360 16082 16416
rect 15750 8472 15806 8528
rect 15750 8200 15806 8256
rect 15566 7284 15568 7304
rect 15568 7284 15620 7304
rect 15620 7284 15622 7304
rect 15566 7248 15622 7284
rect 15934 10412 15936 10432
rect 15936 10412 15988 10432
rect 15988 10412 15990 10432
rect 15934 10376 15990 10412
rect 17958 21120 18014 21176
rect 16670 18536 16726 18592
rect 16394 17312 16450 17368
rect 16946 17076 16948 17096
rect 16948 17076 17000 17096
rect 17000 17076 17002 17096
rect 16946 17040 17002 17076
rect 16210 15680 16266 15736
rect 16394 15680 16450 15736
rect 16302 13776 16358 13832
rect 16486 14320 16542 14376
rect 16210 12552 16266 12608
rect 16394 12688 16450 12744
rect 16302 11892 16358 11928
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 17682 18808 17738 18864
rect 18050 18536 18106 18592
rect 17866 18264 17922 18320
rect 17130 15852 17132 15872
rect 17132 15852 17184 15872
rect 17184 15852 17186 15872
rect 17130 15816 17186 15852
rect 17130 14864 17186 14920
rect 17038 14592 17094 14648
rect 17038 14184 17094 14240
rect 16762 12688 16818 12744
rect 16670 12416 16726 12472
rect 16302 11872 16304 11892
rect 16304 11872 16356 11892
rect 16356 11872 16358 11892
rect 16394 11328 16450 11384
rect 16302 10784 16358 10840
rect 16486 9424 16542 9480
rect 16854 12144 16910 12200
rect 16762 11736 16818 11792
rect 16670 11620 16726 11656
rect 16670 11600 16672 11620
rect 16672 11600 16724 11620
rect 16724 11600 16726 11620
rect 15934 8336 15990 8392
rect 15658 6704 15714 6760
rect 15658 6604 15660 6624
rect 15660 6604 15712 6624
rect 15712 6604 15714 6624
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14922 4528 14978 4584
rect 14738 4256 14794 4312
rect 14922 4256 14978 4312
rect 15198 4004 15254 4040
rect 15198 3984 15200 4004
rect 15200 3984 15252 4004
rect 15252 3984 15254 4004
rect 14646 3440 14702 3496
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14830 3576 14886 3632
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 15658 6568 15714 6604
rect 15566 6296 15622 6352
rect 15934 6704 15990 6760
rect 16118 3984 16174 4040
rect 17406 15020 17462 15056
rect 17406 15000 17408 15020
rect 17408 15000 17460 15020
rect 17460 15000 17462 15020
rect 17314 12960 17370 13016
rect 17222 12552 17278 12608
rect 17314 12144 17370 12200
rect 16762 6568 16818 6624
rect 16670 6024 16726 6080
rect 16302 3168 16358 3224
rect 16578 4936 16634 4992
rect 16578 4120 16634 4176
rect 16578 2488 16634 2544
rect 17866 17312 17922 17368
rect 17958 17040 18014 17096
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18326 18284 18382 18320
rect 18326 18264 18328 18284
rect 18328 18264 18380 18284
rect 18380 18264 18382 18284
rect 18418 17856 18474 17912
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18786 17176 18842 17232
rect 18694 17040 18750 17096
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18786 16088 18842 16144
rect 17958 15000 18014 15056
rect 17498 12416 17554 12472
rect 17866 12688 17922 12744
rect 18050 14320 18106 14376
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18694 15408 18750 15464
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18602 13368 18658 13424
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18510 12688 18566 12744
rect 18050 12552 18106 12608
rect 17774 12008 17830 12064
rect 17590 11192 17646 11248
rect 17038 6840 17094 6896
rect 17958 10648 18014 10704
rect 17774 9560 17830 9616
rect 17406 8744 17462 8800
rect 17682 8608 17738 8664
rect 17406 7792 17462 7848
rect 17590 7792 17646 7848
rect 17222 6296 17278 6352
rect 17130 4256 17186 4312
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18694 13132 18696 13152
rect 18696 13132 18748 13152
rect 18748 13132 18750 13152
rect 18694 13096 18750 13132
rect 18694 11736 18750 11792
rect 18694 11500 18696 11520
rect 18696 11500 18748 11520
rect 18748 11500 18750 11520
rect 18694 11464 18750 11500
rect 18510 11056 18566 11112
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18510 9324 18512 9344
rect 18512 9324 18564 9344
rect 18564 9324 18566 9344
rect 18510 9288 18566 9324
rect 18510 9052 18512 9072
rect 18512 9052 18564 9072
rect 18564 9052 18566 9072
rect 18510 9016 18566 9052
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 17958 7792 18014 7848
rect 17958 7520 18014 7576
rect 17958 6840 18014 6896
rect 17498 6296 17554 6352
rect 17130 2508 17186 2544
rect 17130 2488 17132 2508
rect 17132 2488 17184 2508
rect 17184 2488 17186 2508
rect 17314 3032 17370 3088
rect 17498 5652 17500 5672
rect 17500 5652 17552 5672
rect 17552 5652 17554 5672
rect 17498 5616 17554 5652
rect 17958 6024 18014 6080
rect 17958 4392 18014 4448
rect 18326 8336 18382 8392
rect 18602 8336 18658 8392
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18510 7384 18566 7440
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18878 9444 18934 9480
rect 18878 9424 18880 9444
rect 18880 9424 18932 9444
rect 18932 9424 18934 9444
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18510 5108 18512 5128
rect 18512 5108 18564 5128
rect 18564 5108 18566 5128
rect 18510 5072 18566 5108
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18234 3440 18290 3496
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18418 3052 18474 3088
rect 18418 3032 18420 3052
rect 18420 3032 18472 3052
rect 18472 3032 18474 3052
rect 18326 2352 18382 2408
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 18694 3032 18750 3088
rect 18694 2760 18750 2816
rect 18786 2644 18842 2680
rect 18786 2624 18788 2644
rect 18788 2624 18840 2644
rect 18840 2624 18842 2644
rect 19890 22072 19946 22128
rect 19246 17992 19302 18048
rect 19338 17856 19394 17912
rect 19154 17212 19156 17232
rect 19156 17212 19208 17232
rect 19208 17212 19210 17232
rect 19154 17176 19210 17212
rect 19154 17076 19156 17096
rect 19156 17076 19208 17096
rect 19208 17076 19210 17096
rect 19154 17040 19210 17076
rect 19246 15952 19302 16008
rect 19246 13232 19302 13288
rect 19522 12980 19578 13016
rect 19522 12960 19524 12980
rect 19524 12960 19576 12980
rect 19576 12960 19578 12980
rect 19338 9424 19394 9480
rect 19154 8472 19210 8528
rect 19062 7384 19118 7440
rect 19154 2760 19210 2816
rect 19338 8472 19394 8528
rect 19338 8064 19394 8120
rect 19338 5752 19394 5808
rect 19890 17720 19946 17776
rect 20534 21664 20590 21720
rect 20258 19352 20314 19408
rect 19798 15952 19854 16008
rect 19706 13404 19708 13424
rect 19708 13404 19760 13424
rect 19760 13404 19762 13424
rect 19706 13368 19762 13404
rect 19706 12688 19762 12744
rect 20626 20712 20682 20768
rect 21086 20168 21142 20224
rect 20994 19760 21050 19816
rect 21086 19216 21142 19272
rect 21270 18808 21326 18864
rect 21086 18264 21142 18320
rect 22006 17876 22062 17912
rect 22006 17856 22008 17876
rect 22008 17856 22060 17876
rect 22060 17856 22062 17876
rect 20718 17584 20774 17640
rect 20442 16904 20498 16960
rect 20350 15952 20406 16008
rect 20074 14456 20130 14512
rect 19706 9560 19762 9616
rect 20074 9968 20130 10024
rect 20074 9560 20130 9616
rect 19982 9152 20038 9208
rect 19798 4684 19854 4720
rect 19798 4664 19800 4684
rect 19800 4664 19852 4684
rect 19852 4664 19854 4684
rect 20442 12960 20498 13016
rect 20442 11056 20498 11112
rect 20350 8336 20406 8392
rect 20166 5480 20222 5536
rect 20626 14456 20682 14512
rect 20994 17312 21050 17368
rect 21086 16360 21142 16416
rect 21454 15408 21510 15464
rect 21362 14048 21418 14104
rect 20626 10240 20682 10296
rect 20626 8492 20682 8528
rect 20626 8472 20628 8492
rect 20628 8472 20680 8492
rect 20680 8472 20682 8492
rect 20350 584 20406 640
rect 20534 5208 20590 5264
rect 20534 4800 20590 4856
rect 21270 13504 21326 13560
rect 21546 12552 21602 12608
rect 20626 1536 20682 1592
rect 20994 2796 20996 2816
rect 20996 2796 21048 2816
rect 21048 2796 21050 2816
rect 20994 2760 21050 2796
rect 21086 2488 21142 2544
rect 20994 2080 21050 2136
rect 3882 176 3938 232
rect 21730 8064 21786 8120
rect 22374 10104 22430 10160
rect 22374 9832 22430 9888
rect 22374 6024 22430 6080
rect 21730 1128 21786 1184
rect 22374 4392 22430 4448
rect 21454 176 21510 232
<< metal3 >>
rect 0 22674 480 22704
rect 1853 22674 1919 22677
rect 0 22672 1919 22674
rect 0 22616 1858 22672
rect 1914 22616 1919 22672
rect 0 22614 1919 22616
rect 0 22584 480 22614
rect 1853 22611 1919 22614
rect 20437 22674 20503 22677
rect 22520 22674 23000 22704
rect 20437 22672 23000 22674
rect 20437 22616 20442 22672
rect 20498 22616 23000 22672
rect 20437 22614 23000 22616
rect 20437 22611 20503 22614
rect 22520 22584 23000 22614
rect 0 22130 480 22160
rect 2865 22130 2931 22133
rect 0 22128 2931 22130
rect 0 22072 2870 22128
rect 2926 22072 2931 22128
rect 0 22070 2931 22072
rect 0 22040 480 22070
rect 2865 22067 2931 22070
rect 19885 22130 19951 22133
rect 22520 22130 23000 22160
rect 19885 22128 23000 22130
rect 19885 22072 19890 22128
rect 19946 22072 23000 22128
rect 19885 22070 23000 22072
rect 19885 22067 19951 22070
rect 22520 22040 23000 22070
rect 0 21722 480 21752
rect 2957 21722 3023 21725
rect 0 21720 3023 21722
rect 0 21664 2962 21720
rect 3018 21664 3023 21720
rect 0 21662 3023 21664
rect 0 21632 480 21662
rect 2957 21659 3023 21662
rect 20529 21722 20595 21725
rect 22520 21722 23000 21752
rect 20529 21720 23000 21722
rect 20529 21664 20534 21720
rect 20590 21664 23000 21720
rect 20529 21662 23000 21664
rect 20529 21659 20595 21662
rect 22520 21632 23000 21662
rect 0 21178 480 21208
rect 1945 21178 2011 21181
rect 0 21176 2011 21178
rect 0 21120 1950 21176
rect 2006 21120 2011 21176
rect 0 21118 2011 21120
rect 0 21088 480 21118
rect 1945 21115 2011 21118
rect 17953 21178 18019 21181
rect 22520 21178 23000 21208
rect 17953 21176 23000 21178
rect 17953 21120 17958 21176
rect 18014 21120 23000 21176
rect 17953 21118 23000 21120
rect 17953 21115 18019 21118
rect 22520 21088 23000 21118
rect 0 20770 480 20800
rect 2773 20770 2839 20773
rect 0 20768 2839 20770
rect 0 20712 2778 20768
rect 2834 20712 2839 20768
rect 0 20710 2839 20712
rect 0 20680 480 20710
rect 2773 20707 2839 20710
rect 20621 20770 20687 20773
rect 22520 20770 23000 20800
rect 20621 20768 23000 20770
rect 20621 20712 20626 20768
rect 20682 20712 23000 20768
rect 20621 20710 23000 20712
rect 20621 20707 20687 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22520 20680 23000 20710
rect 18270 20639 18590 20640
rect 0 20226 480 20256
rect 3049 20226 3115 20229
rect 0 20224 3115 20226
rect 0 20168 3054 20224
rect 3110 20168 3115 20224
rect 0 20166 3115 20168
rect 0 20136 480 20166
rect 3049 20163 3115 20166
rect 21081 20226 21147 20229
rect 22520 20226 23000 20256
rect 21081 20224 23000 20226
rect 21081 20168 21086 20224
rect 21142 20168 23000 20224
rect 21081 20166 23000 20168
rect 21081 20163 21147 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 22520 20136 23000 20166
rect 14805 20095 15125 20096
rect 0 19818 480 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 480 19758
rect 1853 19755 1919 19758
rect 2313 19818 2379 19821
rect 5809 19818 5875 19821
rect 2313 19816 5875 19818
rect 2313 19760 2318 19816
rect 2374 19760 5814 19816
rect 5870 19760 5875 19816
rect 2313 19758 5875 19760
rect 2313 19755 2379 19758
rect 5809 19755 5875 19758
rect 20989 19818 21055 19821
rect 22520 19818 23000 19848
rect 20989 19816 23000 19818
rect 20989 19760 20994 19816
rect 21050 19760 23000 19816
rect 20989 19758 23000 19760
rect 20989 19755 21055 19758
rect 22520 19728 23000 19758
rect 13854 19620 13860 19684
rect 13924 19682 13930 19684
rect 13997 19682 14063 19685
rect 13924 19680 14063 19682
rect 13924 19624 14002 19680
rect 14058 19624 14063 19680
rect 13924 19622 14063 19624
rect 13924 19620 13930 19622
rect 13997 19619 14063 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 12249 19410 12315 19413
rect 14457 19410 14523 19413
rect 12249 19408 14523 19410
rect 12249 19352 12254 19408
rect 12310 19352 14462 19408
rect 14518 19352 14523 19408
rect 12249 19350 14523 19352
rect 12249 19347 12315 19350
rect 14457 19347 14523 19350
rect 20253 19412 20319 19413
rect 20253 19408 20300 19412
rect 20364 19410 20370 19412
rect 20253 19352 20258 19408
rect 20253 19348 20300 19352
rect 20364 19350 20410 19410
rect 20364 19348 20370 19350
rect 20253 19347 20319 19348
rect 0 19274 480 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 480 19214
rect 1945 19211 2011 19214
rect 7649 19274 7715 19277
rect 9213 19274 9279 19277
rect 7649 19272 9279 19274
rect 7649 19216 7654 19272
rect 7710 19216 9218 19272
rect 9274 19216 9279 19272
rect 7649 19214 9279 19216
rect 7649 19211 7715 19214
rect 9213 19211 9279 19214
rect 9581 19274 9647 19277
rect 15193 19274 15259 19277
rect 9581 19272 15259 19274
rect 9581 19216 9586 19272
rect 9642 19216 15198 19272
rect 15254 19216 15259 19272
rect 9581 19214 15259 19216
rect 9581 19211 9647 19214
rect 15193 19211 15259 19214
rect 21081 19274 21147 19277
rect 22520 19274 23000 19304
rect 21081 19272 23000 19274
rect 21081 19216 21086 19272
rect 21142 19216 23000 19272
rect 21081 19214 23000 19216
rect 21081 19211 21147 19214
rect 22520 19184 23000 19214
rect 8334 19076 8340 19140
rect 8404 19138 8410 19140
rect 11605 19138 11671 19141
rect 11789 19140 11855 19141
rect 11789 19138 11836 19140
rect 8404 19136 11671 19138
rect 8404 19080 11610 19136
rect 11666 19080 11671 19136
rect 8404 19078 11671 19080
rect 11744 19136 11836 19138
rect 11744 19080 11794 19136
rect 11744 19078 11836 19080
rect 8404 19076 8410 19078
rect 11605 19075 11671 19078
rect 11789 19076 11836 19078
rect 11900 19076 11906 19140
rect 12525 19138 12591 19141
rect 13353 19138 13419 19141
rect 12525 19136 13419 19138
rect 12525 19080 12530 19136
rect 12586 19080 13358 19136
rect 13414 19080 13419 19136
rect 12525 19078 13419 19080
rect 11789 19075 11855 19076
rect 12525 19075 12591 19078
rect 13353 19075 13419 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 2037 19002 2103 19005
rect 3233 19002 3299 19005
rect 5257 19002 5323 19005
rect 2037 19000 5323 19002
rect 2037 18944 2042 19000
rect 2098 18944 3238 19000
rect 3294 18944 5262 19000
rect 5318 18944 5323 19000
rect 2037 18942 5323 18944
rect 2037 18939 2103 18942
rect 3233 18939 3299 18942
rect 5257 18939 5323 18942
rect 10910 18940 10916 19004
rect 10980 19002 10986 19004
rect 11421 19002 11487 19005
rect 10980 19000 11487 19002
rect 10980 18944 11426 19000
rect 11482 18944 11487 19000
rect 10980 18942 11487 18944
rect 10980 18940 10986 18942
rect 11421 18939 11487 18942
rect 11605 19002 11671 19005
rect 12382 19002 12388 19004
rect 11605 19000 12388 19002
rect 11605 18944 11610 19000
rect 11666 18944 12388 19000
rect 11605 18942 12388 18944
rect 11605 18939 11671 18942
rect 12382 18940 12388 18942
rect 12452 19002 12458 19004
rect 12452 18942 14106 19002
rect 12452 18940 12458 18942
rect 0 18866 480 18896
rect 2773 18866 2839 18869
rect 0 18864 2839 18866
rect 0 18808 2778 18864
rect 2834 18808 2839 18864
rect 0 18806 2839 18808
rect 0 18776 480 18806
rect 2773 18803 2839 18806
rect 11237 18866 11303 18869
rect 13905 18866 13971 18869
rect 11237 18864 13971 18866
rect 11237 18808 11242 18864
rect 11298 18808 13910 18864
rect 13966 18808 13971 18864
rect 11237 18806 13971 18808
rect 14046 18866 14106 18942
rect 17677 18866 17743 18869
rect 14046 18864 17743 18866
rect 14046 18808 17682 18864
rect 17738 18808 17743 18864
rect 14046 18806 17743 18808
rect 11237 18803 11303 18806
rect 13905 18803 13971 18806
rect 17677 18803 17743 18806
rect 21265 18866 21331 18869
rect 22520 18866 23000 18896
rect 21265 18864 23000 18866
rect 21265 18808 21270 18864
rect 21326 18808 23000 18864
rect 21265 18806 23000 18808
rect 21265 18803 21331 18806
rect 22520 18776 23000 18806
rect 5441 18730 5507 18733
rect 10726 18730 10732 18732
rect 5441 18728 10732 18730
rect 5441 18672 5446 18728
rect 5502 18672 10732 18728
rect 5441 18670 10732 18672
rect 5441 18667 5507 18670
rect 10726 18668 10732 18670
rect 10796 18668 10802 18732
rect 12157 18730 12223 18733
rect 13997 18730 14063 18733
rect 12157 18728 14063 18730
rect 12157 18672 12162 18728
rect 12218 18672 14002 18728
rect 14058 18672 14063 18728
rect 12157 18670 14063 18672
rect 12157 18667 12223 18670
rect 13997 18667 14063 18670
rect 10133 18594 10199 18597
rect 10358 18594 10364 18596
rect 10133 18592 10364 18594
rect 10133 18536 10138 18592
rect 10194 18536 10364 18592
rect 10133 18534 10364 18536
rect 10133 18531 10199 18534
rect 10358 18532 10364 18534
rect 10428 18532 10434 18596
rect 12709 18594 12775 18597
rect 16665 18594 16731 18597
rect 18045 18594 18111 18597
rect 12709 18592 18111 18594
rect 12709 18536 12714 18592
rect 12770 18536 16670 18592
rect 16726 18536 18050 18592
rect 18106 18536 18111 18592
rect 12709 18534 18111 18536
rect 12709 18531 12775 18534
rect 16665 18531 16731 18534
rect 18045 18531 18111 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 4889 18458 4955 18461
rect 8334 18458 8340 18460
rect 4889 18456 8340 18458
rect 4889 18400 4894 18456
rect 4950 18400 8340 18456
rect 4889 18398 8340 18400
rect 4889 18395 4955 18398
rect 8334 18396 8340 18398
rect 8404 18396 8410 18460
rect 0 18322 480 18352
rect 1485 18322 1551 18325
rect 0 18320 1551 18322
rect 0 18264 1490 18320
rect 1546 18264 1551 18320
rect 0 18262 1551 18264
rect 0 18232 480 18262
rect 1485 18259 1551 18262
rect 17861 18322 17927 18325
rect 18321 18322 18387 18325
rect 17861 18320 18387 18322
rect 17861 18264 17866 18320
rect 17922 18264 18326 18320
rect 18382 18264 18387 18320
rect 17861 18262 18387 18264
rect 17861 18259 17927 18262
rect 18321 18259 18387 18262
rect 21081 18322 21147 18325
rect 22520 18322 23000 18352
rect 21081 18320 23000 18322
rect 21081 18264 21086 18320
rect 21142 18264 23000 18320
rect 21081 18262 23000 18264
rect 21081 18259 21147 18262
rect 22520 18232 23000 18262
rect 14825 18186 14891 18189
rect 11240 18184 14891 18186
rect 11240 18128 14830 18184
rect 14886 18128 14891 18184
rect 11240 18126 14891 18128
rect 10961 18050 11027 18053
rect 11240 18050 11300 18126
rect 14825 18123 14891 18126
rect 10961 18048 11300 18050
rect 10961 17992 10966 18048
rect 11022 17992 11300 18048
rect 10961 17990 11300 17992
rect 12065 18050 12131 18053
rect 12433 18050 12499 18053
rect 12065 18048 12499 18050
rect 12065 17992 12070 18048
rect 12126 17992 12438 18048
rect 12494 17992 12499 18048
rect 12065 17990 12499 17992
rect 10961 17987 11027 17990
rect 12065 17987 12131 17990
rect 12433 17987 12499 17990
rect 15193 18050 15259 18053
rect 19241 18050 19307 18053
rect 15193 18048 19307 18050
rect 15193 17992 15198 18048
rect 15254 17992 19246 18048
rect 19302 17992 19307 18048
rect 15193 17990 19307 17992
rect 15193 17987 15259 17990
rect 19241 17987 19307 17990
rect 7874 17984 8194 17985
rect 0 17914 480 17944
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 1577 17914 1643 17917
rect 0 17912 1643 17914
rect 0 17856 1582 17912
rect 1638 17856 1643 17912
rect 0 17854 1643 17856
rect 0 17824 480 17854
rect 1577 17851 1643 17854
rect 8661 17914 8727 17917
rect 9397 17914 9463 17917
rect 12801 17914 12867 17917
rect 8661 17912 12867 17914
rect 8661 17856 8666 17912
rect 8722 17856 9402 17912
rect 9458 17856 12806 17912
rect 12862 17856 12867 17912
rect 8661 17854 12867 17856
rect 8661 17851 8727 17854
rect 9397 17851 9463 17854
rect 12801 17851 12867 17854
rect 18413 17914 18479 17917
rect 19333 17914 19399 17917
rect 18413 17912 19399 17914
rect 18413 17856 18418 17912
rect 18474 17856 19338 17912
rect 19394 17856 19399 17912
rect 18413 17854 19399 17856
rect 18413 17851 18479 17854
rect 19333 17851 19399 17854
rect 22001 17914 22067 17917
rect 22520 17914 23000 17944
rect 22001 17912 23000 17914
rect 22001 17856 22006 17912
rect 22062 17856 23000 17912
rect 22001 17854 23000 17856
rect 22001 17851 22067 17854
rect 22520 17824 23000 17854
rect 7598 17716 7604 17780
rect 7668 17778 7674 17780
rect 7741 17778 7807 17781
rect 19885 17778 19951 17781
rect 7668 17776 19951 17778
rect 7668 17720 7746 17776
rect 7802 17720 19890 17776
rect 19946 17720 19951 17776
rect 7668 17718 19951 17720
rect 7668 17716 7674 17718
rect 7741 17715 7807 17718
rect 19885 17715 19951 17718
rect 8518 17580 8524 17644
rect 8588 17642 8594 17644
rect 9673 17642 9739 17645
rect 8588 17640 9739 17642
rect 8588 17584 9678 17640
rect 9734 17584 9739 17640
rect 8588 17582 9739 17584
rect 8588 17580 8594 17582
rect 9673 17579 9739 17582
rect 11053 17642 11119 17645
rect 12893 17642 12959 17645
rect 13997 17642 14063 17645
rect 20713 17642 20779 17645
rect 11053 17640 14063 17642
rect 11053 17584 11058 17640
rect 11114 17584 12898 17640
rect 12954 17584 14002 17640
rect 14058 17584 14063 17640
rect 11053 17582 14063 17584
rect 11053 17579 11119 17582
rect 12893 17579 12959 17582
rect 13997 17579 14063 17582
rect 14184 17640 20779 17642
rect 14184 17584 20718 17640
rect 20774 17584 20779 17640
rect 14184 17582 20779 17584
rect 7465 17506 7531 17509
rect 10961 17506 11027 17509
rect 7465 17504 11027 17506
rect 7465 17448 7470 17504
rect 7526 17448 10966 17504
rect 11022 17448 11027 17504
rect 7465 17446 11027 17448
rect 7465 17443 7531 17446
rect 10961 17443 11027 17446
rect 12157 17506 12223 17509
rect 13670 17506 13676 17508
rect 12157 17504 13676 17506
rect 12157 17448 12162 17504
rect 12218 17448 13676 17504
rect 12157 17446 13676 17448
rect 12157 17443 12223 17446
rect 13670 17444 13676 17446
rect 13740 17506 13746 17508
rect 14184 17506 14244 17582
rect 20713 17579 20779 17582
rect 13740 17446 14244 17506
rect 13740 17444 13746 17446
rect 4409 17440 4729 17441
rect 0 17370 480 17400
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 480 17310
rect 1577 17307 1643 17310
rect 6637 17370 6703 17373
rect 8886 17370 8892 17372
rect 6637 17368 8892 17370
rect 6637 17312 6642 17368
rect 6698 17312 8892 17368
rect 6637 17310 8892 17312
rect 6637 17307 6703 17310
rect 8886 17308 8892 17310
rect 8956 17370 8962 17372
rect 11145 17370 11211 17373
rect 8956 17368 11211 17370
rect 8956 17312 11150 17368
rect 11206 17312 11211 17368
rect 8956 17310 11211 17312
rect 8956 17308 8962 17310
rect 11145 17307 11211 17310
rect 12249 17370 12315 17373
rect 16389 17370 16455 17373
rect 17861 17370 17927 17373
rect 12249 17368 17927 17370
rect 12249 17312 12254 17368
rect 12310 17312 16394 17368
rect 16450 17312 17866 17368
rect 17922 17312 17927 17368
rect 12249 17310 17927 17312
rect 12249 17307 12315 17310
rect 16389 17307 16455 17310
rect 17861 17307 17927 17310
rect 20989 17370 21055 17373
rect 22520 17370 23000 17400
rect 20989 17368 23000 17370
rect 20989 17312 20994 17368
rect 21050 17312 23000 17368
rect 20989 17310 23000 17312
rect 20989 17307 21055 17310
rect 22520 17280 23000 17310
rect 7373 17234 7439 17237
rect 10317 17234 10383 17237
rect 7373 17232 10383 17234
rect 7373 17176 7378 17232
rect 7434 17176 10322 17232
rect 10378 17176 10383 17232
rect 7373 17174 10383 17176
rect 7373 17171 7439 17174
rect 10317 17171 10383 17174
rect 11881 17234 11947 17237
rect 12566 17234 12572 17236
rect 11881 17232 12572 17234
rect 11881 17176 11886 17232
rect 11942 17176 12572 17232
rect 11881 17174 12572 17176
rect 11881 17171 11947 17174
rect 12566 17172 12572 17174
rect 12636 17172 12642 17236
rect 13813 17234 13879 17237
rect 14038 17234 14044 17236
rect 13813 17232 14044 17234
rect 13813 17176 13818 17232
rect 13874 17176 14044 17232
rect 13813 17174 14044 17176
rect 13813 17171 13879 17174
rect 14038 17172 14044 17174
rect 14108 17172 14114 17236
rect 18781 17234 18847 17237
rect 19149 17234 19215 17237
rect 18781 17232 19215 17234
rect 18781 17176 18786 17232
rect 18842 17176 19154 17232
rect 19210 17176 19215 17232
rect 18781 17174 19215 17176
rect 18781 17171 18847 17174
rect 19149 17171 19215 17174
rect 5809 17098 5875 17101
rect 9806 17098 9812 17100
rect 5809 17096 9812 17098
rect 5809 17040 5814 17096
rect 5870 17040 9812 17096
rect 5809 17038 9812 17040
rect 5809 17035 5875 17038
rect 9806 17036 9812 17038
rect 9876 17036 9882 17100
rect 10726 17036 10732 17100
rect 10796 17098 10802 17100
rect 13997 17098 14063 17101
rect 16941 17098 17007 17101
rect 10796 17096 14063 17098
rect 10796 17040 14002 17096
rect 14058 17040 14063 17096
rect 10796 17038 14063 17040
rect 10796 17036 10802 17038
rect 0 16962 480 16992
rect 1485 16962 1551 16965
rect 0 16960 1551 16962
rect 0 16904 1490 16960
rect 1546 16904 1551 16960
rect 0 16902 1551 16904
rect 9814 16962 9874 17036
rect 13997 17035 14063 17038
rect 14368 17096 17007 17098
rect 14368 17040 16946 17096
rect 17002 17040 17007 17096
rect 14368 17038 17007 17040
rect 11145 16962 11211 16965
rect 9814 16960 11211 16962
rect 9814 16904 11150 16960
rect 11206 16904 11211 16960
rect 9814 16902 11211 16904
rect 0 16872 480 16902
rect 1485 16899 1551 16902
rect 11145 16899 11211 16902
rect 12566 16900 12572 16964
rect 12636 16962 12642 16964
rect 14368 16962 14428 17038
rect 16941 17035 17007 17038
rect 17953 17098 18019 17101
rect 18086 17098 18092 17100
rect 17953 17096 18092 17098
rect 17953 17040 17958 17096
rect 18014 17040 18092 17096
rect 17953 17038 18092 17040
rect 17953 17035 18019 17038
rect 18086 17036 18092 17038
rect 18156 17036 18162 17100
rect 18689 17098 18755 17101
rect 19006 17098 19012 17100
rect 18689 17096 19012 17098
rect 18689 17040 18694 17096
rect 18750 17040 19012 17096
rect 18689 17038 19012 17040
rect 18689 17035 18755 17038
rect 19006 17036 19012 17038
rect 19076 17098 19082 17100
rect 19149 17098 19215 17101
rect 19076 17096 19215 17098
rect 19076 17040 19154 17096
rect 19210 17040 19215 17096
rect 19076 17038 19215 17040
rect 19076 17036 19082 17038
rect 19149 17035 19215 17038
rect 12636 16902 14428 16962
rect 20437 16962 20503 16965
rect 22520 16962 23000 16992
rect 20437 16960 23000 16962
rect 20437 16904 20442 16960
rect 20498 16904 23000 16960
rect 20437 16902 23000 16904
rect 12636 16900 12642 16902
rect 20437 16899 20503 16902
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 22520 16872 23000 16902
rect 14805 16831 15125 16832
rect 4061 16824 4127 16829
rect 9213 16828 9279 16829
rect 9213 16826 9260 16828
rect 4061 16768 4066 16824
rect 4122 16768 4127 16824
rect 4061 16763 4127 16768
rect 9168 16824 9260 16826
rect 9168 16768 9218 16824
rect 9168 16766 9260 16768
rect 9213 16764 9260 16766
rect 9324 16764 9330 16828
rect 10174 16764 10180 16828
rect 10244 16826 10250 16828
rect 14181 16826 14247 16829
rect 10244 16824 14247 16826
rect 10244 16768 14186 16824
rect 14242 16768 14247 16824
rect 10244 16766 14247 16768
rect 10244 16764 10250 16766
rect 9213 16763 9279 16764
rect 14181 16763 14247 16766
rect 2497 16690 2563 16693
rect 4064 16690 4124 16763
rect 8661 16690 8727 16693
rect 2497 16688 8727 16690
rect 2497 16632 2502 16688
rect 2558 16632 8666 16688
rect 8722 16632 8727 16688
rect 2497 16630 8727 16632
rect 2497 16627 2563 16630
rect 8661 16627 8727 16630
rect 1669 16554 1735 16557
rect 7414 16554 7420 16556
rect 1669 16552 7420 16554
rect 1669 16496 1674 16552
rect 1730 16496 7420 16552
rect 1669 16494 7420 16496
rect 1669 16491 1735 16494
rect 7414 16492 7420 16494
rect 7484 16554 7490 16556
rect 7925 16554 7991 16557
rect 7484 16552 7991 16554
rect 7484 16496 7930 16552
rect 7986 16496 7991 16552
rect 7484 16494 7991 16496
rect 7484 16492 7490 16494
rect 7925 16491 7991 16494
rect 11145 16554 11211 16557
rect 11145 16552 11852 16554
rect 11145 16496 11150 16552
rect 11206 16496 11852 16552
rect 11145 16494 11852 16496
rect 11145 16491 11211 16494
rect 0 16418 480 16448
rect 1669 16418 1735 16421
rect 0 16416 1735 16418
rect 0 16360 1674 16416
rect 1730 16360 1735 16416
rect 0 16358 1735 16360
rect 0 16328 480 16358
rect 1669 16355 1735 16358
rect 7373 16418 7439 16421
rect 8937 16418 9003 16421
rect 7373 16416 9003 16418
rect 7373 16360 7378 16416
rect 7434 16360 8942 16416
rect 8998 16360 9003 16416
rect 7373 16358 9003 16360
rect 11792 16418 11852 16494
rect 16021 16418 16087 16421
rect 11792 16416 16087 16418
rect 11792 16360 16026 16416
rect 16082 16360 16087 16416
rect 11792 16358 16087 16360
rect 7373 16355 7439 16358
rect 8937 16355 9003 16358
rect 16021 16355 16087 16358
rect 21081 16418 21147 16421
rect 22520 16418 23000 16448
rect 21081 16416 23000 16418
rect 21081 16360 21086 16416
rect 21142 16360 23000 16416
rect 21081 16358 23000 16360
rect 21081 16355 21147 16358
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 22520 16328 23000 16358
rect 18270 16287 18590 16288
rect 7097 16282 7163 16285
rect 9581 16282 9647 16285
rect 7097 16280 9647 16282
rect 7097 16224 7102 16280
rect 7158 16224 9586 16280
rect 9642 16224 9647 16280
rect 7097 16222 9647 16224
rect 7097 16219 7163 16222
rect 9581 16219 9647 16222
rect 1945 16146 2011 16149
rect 5993 16146 6059 16149
rect 1945 16144 6059 16146
rect 1945 16088 1950 16144
rect 2006 16088 5998 16144
rect 6054 16088 6059 16144
rect 1945 16086 6059 16088
rect 1945 16083 2011 16086
rect 5993 16083 6059 16086
rect 10358 16084 10364 16148
rect 10428 16146 10434 16148
rect 18781 16146 18847 16149
rect 10428 16144 18847 16146
rect 10428 16088 18786 16144
rect 18842 16088 18847 16144
rect 10428 16086 18847 16088
rect 10428 16084 10434 16086
rect 18781 16083 18847 16086
rect 0 16010 480 16040
rect 1853 16010 1919 16013
rect 9489 16010 9555 16013
rect 0 16008 1919 16010
rect 0 15952 1858 16008
rect 1914 15952 1919 16008
rect 0 15950 1919 15952
rect 0 15920 480 15950
rect 1853 15947 1919 15950
rect 5766 16008 9555 16010
rect 5766 15952 9494 16008
rect 9550 15952 9555 16008
rect 5766 15950 9555 15952
rect 3417 15874 3483 15877
rect 3877 15874 3943 15877
rect 5766 15874 5826 15950
rect 9489 15947 9555 15950
rect 9765 16010 9831 16013
rect 10542 16010 10548 16012
rect 9765 16008 10548 16010
rect 9765 15952 9770 16008
rect 9826 15952 10548 16008
rect 9765 15950 10548 15952
rect 9765 15947 9831 15950
rect 10542 15948 10548 15950
rect 10612 15948 10618 16012
rect 10910 15948 10916 16012
rect 10980 16010 10986 16012
rect 11145 16010 11211 16013
rect 10980 16008 11211 16010
rect 10980 15952 11150 16008
rect 11206 15952 11211 16008
rect 10980 15950 11211 15952
rect 10980 15948 10986 15950
rect 11145 15947 11211 15950
rect 11830 15948 11836 16012
rect 11900 16010 11906 16012
rect 19241 16010 19307 16013
rect 11900 16008 19307 16010
rect 11900 15952 19246 16008
rect 19302 15952 19307 16008
rect 11900 15950 19307 15952
rect 11900 15948 11906 15950
rect 19241 15947 19307 15950
rect 19374 15948 19380 16012
rect 19444 16010 19450 16012
rect 19793 16010 19859 16013
rect 19444 16008 19859 16010
rect 19444 15952 19798 16008
rect 19854 15952 19859 16008
rect 19444 15950 19859 15952
rect 19444 15948 19450 15950
rect 19793 15947 19859 15950
rect 20345 16010 20411 16013
rect 22520 16010 23000 16040
rect 20345 16008 23000 16010
rect 20345 15952 20350 16008
rect 20406 15952 23000 16008
rect 20345 15950 23000 15952
rect 20345 15947 20411 15950
rect 22520 15920 23000 15950
rect 3417 15872 5826 15874
rect 3417 15816 3422 15872
rect 3478 15816 3882 15872
rect 3938 15816 5826 15872
rect 3417 15814 5826 15816
rect 3417 15811 3483 15814
rect 3877 15811 3943 15814
rect 16982 15812 16988 15876
rect 17052 15874 17058 15876
rect 17125 15874 17191 15877
rect 17052 15872 17191 15874
rect 17052 15816 17130 15872
rect 17186 15816 17191 15872
rect 17052 15814 17191 15816
rect 17052 15812 17058 15814
rect 17125 15811 17191 15814
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 2589 15738 2655 15741
rect 5533 15738 5599 15741
rect 2589 15736 5599 15738
rect 2589 15680 2594 15736
rect 2650 15680 5538 15736
rect 5594 15680 5599 15736
rect 2589 15678 5599 15680
rect 2589 15675 2655 15678
rect 5533 15675 5599 15678
rect 10409 15738 10475 15741
rect 16205 15738 16271 15741
rect 16389 15738 16455 15741
rect 10409 15736 14290 15738
rect 10409 15680 10414 15736
rect 10470 15680 14290 15736
rect 10409 15678 14290 15680
rect 10409 15675 10475 15678
rect 10317 15602 10383 15605
rect 10593 15602 10659 15605
rect 11145 15602 11211 15605
rect 10317 15600 11211 15602
rect 10317 15544 10322 15600
rect 10378 15544 10598 15600
rect 10654 15544 11150 15600
rect 11206 15544 11211 15600
rect 10317 15542 11211 15544
rect 10317 15539 10383 15542
rect 10593 15539 10659 15542
rect 11145 15539 11211 15542
rect 11697 15602 11763 15605
rect 12617 15602 12683 15605
rect 14230 15604 14290 15678
rect 16205 15736 16455 15738
rect 16205 15680 16210 15736
rect 16266 15680 16394 15736
rect 16450 15680 16455 15736
rect 16205 15678 16455 15680
rect 16205 15675 16271 15678
rect 16389 15675 16455 15678
rect 11697 15600 12683 15602
rect 11697 15544 11702 15600
rect 11758 15544 12622 15600
rect 12678 15544 12683 15600
rect 11697 15542 12683 15544
rect 11697 15539 11763 15542
rect 12617 15539 12683 15542
rect 14222 15540 14228 15604
rect 14292 15602 14298 15604
rect 14641 15602 14707 15605
rect 14292 15600 14707 15602
rect 14292 15544 14646 15600
rect 14702 15544 14707 15600
rect 14292 15542 14707 15544
rect 14292 15540 14298 15542
rect 14641 15539 14707 15542
rect 0 15466 480 15496
rect 1945 15466 2011 15469
rect 0 15464 2011 15466
rect 0 15408 1950 15464
rect 2006 15408 2011 15464
rect 0 15406 2011 15408
rect 0 15376 480 15406
rect 1945 15403 2011 15406
rect 10133 15466 10199 15469
rect 11697 15466 11763 15469
rect 10133 15464 11763 15466
rect 10133 15408 10138 15464
rect 10194 15408 11702 15464
rect 11758 15408 11763 15464
rect 10133 15406 11763 15408
rect 10133 15403 10199 15406
rect 11697 15403 11763 15406
rect 13629 15466 13695 15469
rect 18689 15466 18755 15469
rect 13629 15464 18755 15466
rect 13629 15408 13634 15464
rect 13690 15408 18694 15464
rect 18750 15408 18755 15464
rect 13629 15406 18755 15408
rect 13629 15403 13695 15406
rect 18689 15403 18755 15406
rect 21449 15466 21515 15469
rect 22520 15466 23000 15496
rect 21449 15464 23000 15466
rect 21449 15408 21454 15464
rect 21510 15408 23000 15464
rect 21449 15406 23000 15408
rect 21449 15403 21515 15406
rect 22520 15376 23000 15406
rect 8017 15330 8083 15333
rect 8753 15330 8819 15333
rect 14457 15332 14523 15333
rect 8017 15328 8819 15330
rect 8017 15272 8022 15328
rect 8078 15272 8758 15328
rect 8814 15272 8819 15328
rect 8017 15270 8819 15272
rect 8017 15267 8083 15270
rect 8753 15267 8819 15270
rect 14406 15268 14412 15332
rect 14476 15330 14523 15332
rect 14476 15328 14568 15330
rect 14518 15272 14568 15328
rect 14476 15270 14568 15272
rect 14476 15268 14523 15270
rect 14457 15267 14523 15268
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 7833 15194 7899 15197
rect 11053 15194 11119 15197
rect 7833 15192 11119 15194
rect 7833 15136 7838 15192
rect 7894 15136 11058 15192
rect 11114 15136 11119 15192
rect 7833 15134 11119 15136
rect 7833 15131 7899 15134
rect 11053 15131 11119 15134
rect 0 15058 480 15088
rect 3509 15058 3575 15061
rect 0 15056 3575 15058
rect 0 15000 3514 15056
rect 3570 15000 3575 15056
rect 0 14998 3575 15000
rect 0 14968 480 14998
rect 3509 14995 3575 14998
rect 8385 15056 8451 15061
rect 8385 15000 8390 15056
rect 8446 15000 8451 15056
rect 8385 14995 8451 15000
rect 9070 14996 9076 15060
rect 9140 15058 9146 15060
rect 9489 15058 9555 15061
rect 9140 15056 9555 15058
rect 9140 15000 9494 15056
rect 9550 15000 9555 15056
rect 9140 14998 9555 15000
rect 9140 14996 9146 14998
rect 9489 14995 9555 14998
rect 14038 14996 14044 15060
rect 14108 15058 14114 15060
rect 17401 15058 17467 15061
rect 14108 15056 17467 15058
rect 14108 15000 17406 15056
rect 17462 15000 17467 15056
rect 14108 14998 17467 15000
rect 14108 14996 14114 14998
rect 17401 14995 17467 14998
rect 17953 15058 18019 15061
rect 22520 15058 23000 15088
rect 17953 15056 23000 15058
rect 17953 15000 17958 15056
rect 18014 15000 23000 15056
rect 17953 14998 23000 15000
rect 17953 14995 18019 14998
rect 8388 14922 8448 14995
rect 22520 14968 23000 14998
rect 9305 14922 9371 14925
rect 8388 14920 9371 14922
rect 8388 14864 9310 14920
rect 9366 14864 9371 14920
rect 8388 14862 9371 14864
rect 9305 14859 9371 14862
rect 15101 14922 15167 14925
rect 17125 14922 17191 14925
rect 15101 14920 17191 14922
rect 15101 14864 15106 14920
rect 15162 14864 17130 14920
rect 17186 14864 17191 14920
rect 15101 14862 17191 14864
rect 15101 14859 15167 14862
rect 17125 14859 17191 14862
rect 7189 14788 7255 14789
rect 7189 14784 7236 14788
rect 7300 14786 7306 14788
rect 7189 14728 7194 14784
rect 7189 14724 7236 14728
rect 7300 14726 7346 14786
rect 7300 14724 7306 14726
rect 7189 14723 7255 14724
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 8569 14650 8635 14653
rect 11789 14650 11855 14653
rect 8569 14648 11855 14650
rect 8569 14592 8574 14648
rect 8630 14592 11794 14648
rect 11850 14592 11855 14648
rect 8569 14590 11855 14592
rect 8569 14587 8635 14590
rect 11789 14587 11855 14590
rect 17033 14650 17099 14653
rect 17166 14650 17172 14652
rect 17033 14648 17172 14650
rect 17033 14592 17038 14648
rect 17094 14592 17172 14648
rect 17033 14590 17172 14592
rect 17033 14587 17099 14590
rect 17166 14588 17172 14590
rect 17236 14588 17242 14652
rect 0 14514 480 14544
rect 1577 14514 1643 14517
rect 0 14512 1643 14514
rect 0 14456 1582 14512
rect 1638 14456 1643 14512
rect 0 14454 1643 14456
rect 0 14424 480 14454
rect 1577 14451 1643 14454
rect 8477 14514 8543 14517
rect 8753 14514 8819 14517
rect 12198 14514 12204 14516
rect 8477 14512 8586 14514
rect 8477 14456 8482 14512
rect 8538 14456 8586 14512
rect 8477 14451 8586 14456
rect 8753 14512 12204 14514
rect 8753 14456 8758 14512
rect 8814 14456 12204 14512
rect 8753 14454 12204 14456
rect 8753 14451 8819 14454
rect 12198 14452 12204 14454
rect 12268 14514 12274 14516
rect 20069 14514 20135 14517
rect 12268 14512 20135 14514
rect 12268 14456 20074 14512
rect 20130 14456 20135 14512
rect 12268 14454 20135 14456
rect 12268 14452 12274 14454
rect 20069 14451 20135 14454
rect 20621 14514 20687 14517
rect 22520 14514 23000 14544
rect 20621 14512 23000 14514
rect 20621 14456 20626 14512
rect 20682 14456 23000 14512
rect 20621 14454 23000 14456
rect 20621 14451 20687 14454
rect 8526 14378 8586 14451
rect 22520 14424 23000 14454
rect 8753 14378 8819 14381
rect 8886 14378 8892 14380
rect 8526 14376 8892 14378
rect 8526 14320 8758 14376
rect 8814 14320 8892 14376
rect 8526 14318 8892 14320
rect 8753 14315 8819 14318
rect 8886 14316 8892 14318
rect 8956 14316 8962 14380
rect 12157 14378 12223 14381
rect 14273 14378 14339 14381
rect 12157 14376 14339 14378
rect 12157 14320 12162 14376
rect 12218 14320 14278 14376
rect 14334 14320 14339 14376
rect 12157 14318 14339 14320
rect 12157 14315 12223 14318
rect 14273 14315 14339 14318
rect 16481 14378 16547 14381
rect 18045 14378 18111 14381
rect 16481 14376 18111 14378
rect 16481 14320 16486 14376
rect 16542 14320 18050 14376
rect 18106 14320 18111 14376
rect 16481 14318 18111 14320
rect 16481 14315 16547 14318
rect 18045 14315 18111 14318
rect 7281 14242 7347 14245
rect 8937 14242 9003 14245
rect 7281 14240 9003 14242
rect 7281 14184 7286 14240
rect 7342 14184 8942 14240
rect 8998 14184 9003 14240
rect 7281 14182 9003 14184
rect 7281 14179 7347 14182
rect 8937 14179 9003 14182
rect 11881 14242 11947 14245
rect 13854 14242 13860 14244
rect 11881 14240 13860 14242
rect 11881 14184 11886 14240
rect 11942 14184 13860 14240
rect 11881 14182 13860 14184
rect 11881 14179 11947 14182
rect 13854 14180 13860 14182
rect 13924 14242 13930 14244
rect 17033 14242 17099 14245
rect 13924 14240 17099 14242
rect 13924 14184 17038 14240
rect 17094 14184 17099 14240
rect 13924 14182 17099 14184
rect 13924 14180 13930 14182
rect 17033 14179 17099 14182
rect 4409 14176 4729 14177
rect 0 14106 480 14136
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 2773 14106 2839 14109
rect 0 14104 2839 14106
rect 0 14048 2778 14104
rect 2834 14048 2839 14104
rect 0 14046 2839 14048
rect 0 14016 480 14046
rect 2773 14043 2839 14046
rect 13353 14106 13419 14109
rect 14273 14106 14339 14109
rect 13353 14104 14339 14106
rect 13353 14048 13358 14104
rect 13414 14048 14278 14104
rect 14334 14048 14339 14104
rect 13353 14046 14339 14048
rect 13353 14043 13419 14046
rect 14273 14043 14339 14046
rect 21357 14106 21423 14109
rect 22520 14106 23000 14136
rect 21357 14104 23000 14106
rect 21357 14048 21362 14104
rect 21418 14048 23000 14104
rect 21357 14046 23000 14048
rect 21357 14043 21423 14046
rect 22520 14016 23000 14046
rect 15377 13970 15443 13973
rect 12620 13968 15443 13970
rect 12620 13912 15382 13968
rect 15438 13912 15443 13968
rect 12620 13910 15443 13912
rect 11421 13834 11487 13837
rect 12620 13834 12680 13910
rect 15377 13907 15443 13910
rect 11421 13832 12680 13834
rect 11421 13776 11426 13832
rect 11482 13776 12680 13832
rect 11421 13774 12680 13776
rect 13353 13834 13419 13837
rect 14825 13834 14891 13837
rect 16297 13834 16363 13837
rect 13353 13832 16363 13834
rect 13353 13776 13358 13832
rect 13414 13776 14830 13832
rect 14886 13776 16302 13832
rect 16358 13776 16363 13832
rect 13353 13774 16363 13776
rect 11421 13771 11487 13774
rect 13353 13771 13419 13774
rect 14825 13771 14891 13774
rect 16297 13771 16363 13774
rect 11421 13698 11487 13701
rect 14365 13698 14431 13701
rect 11421 13696 14431 13698
rect 11421 13640 11426 13696
rect 11482 13640 14370 13696
rect 14426 13640 14431 13696
rect 11421 13638 14431 13640
rect 11421 13635 11487 13638
rect 14365 13635 14431 13638
rect 7874 13632 8194 13633
rect 0 13562 480 13592
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 3601 13562 3667 13565
rect 21265 13562 21331 13565
rect 22520 13562 23000 13592
rect 0 13560 3667 13562
rect 0 13504 3606 13560
rect 3662 13504 3667 13560
rect 0 13502 3667 13504
rect 0 13472 480 13502
rect 3601 13499 3667 13502
rect 11332 13502 12680 13562
rect 6913 13426 6979 13429
rect 11332 13426 11392 13502
rect 4248 13424 11392 13426
rect 4248 13368 6918 13424
rect 6974 13368 11392 13424
rect 4248 13366 11392 13368
rect 11513 13426 11579 13429
rect 12014 13426 12020 13428
rect 11513 13424 12020 13426
rect 11513 13368 11518 13424
rect 11574 13368 12020 13424
rect 11513 13366 12020 13368
rect 0 13154 480 13184
rect 4248 13154 4308 13366
rect 6913 13363 6979 13366
rect 11513 13363 11579 13366
rect 12014 13364 12020 13366
rect 12084 13364 12090 13428
rect 12620 13426 12680 13502
rect 21265 13560 23000 13562
rect 21265 13504 21270 13560
rect 21326 13504 23000 13560
rect 21265 13502 23000 13504
rect 21265 13499 21331 13502
rect 22520 13472 23000 13502
rect 18597 13426 18663 13429
rect 19701 13428 19767 13429
rect 19701 13426 19748 13428
rect 12620 13424 18663 13426
rect 12620 13368 18602 13424
rect 18658 13368 18663 13424
rect 12620 13366 18663 13368
rect 19656 13424 19748 13426
rect 19656 13368 19706 13424
rect 19656 13366 19748 13368
rect 18597 13363 18663 13366
rect 19701 13364 19748 13366
rect 19812 13364 19818 13428
rect 19701 13363 19767 13364
rect 6821 13290 6887 13293
rect 19241 13290 19307 13293
rect 6821 13288 19307 13290
rect 6821 13232 6826 13288
rect 6882 13232 19246 13288
rect 19302 13232 19307 13288
rect 6821 13230 19307 13232
rect 6821 13227 6887 13230
rect 19241 13227 19307 13230
rect 0 13094 4308 13154
rect 13905 13154 13971 13157
rect 18689 13154 18755 13157
rect 22520 13154 23000 13184
rect 13905 13152 18108 13154
rect 13905 13096 13910 13152
rect 13966 13096 18108 13152
rect 13905 13094 18108 13096
rect 0 13064 480 13094
rect 13905 13091 13971 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 14365 13018 14431 13021
rect 17309 13018 17375 13021
rect 14365 13016 17375 13018
rect 14365 12960 14370 13016
rect 14426 12960 17314 13016
rect 17370 12960 17375 13016
rect 14365 12958 17375 12960
rect 14365 12955 14431 12958
rect 17309 12955 17375 12958
rect 2221 12882 2287 12885
rect 5717 12882 5783 12885
rect 2221 12880 5783 12882
rect 2221 12824 2226 12880
rect 2282 12824 5722 12880
rect 5778 12824 5783 12880
rect 2221 12822 5783 12824
rect 2221 12819 2287 12822
rect 5717 12819 5783 12822
rect 12893 12882 12959 12885
rect 18048 12882 18108 13094
rect 18689 13152 23000 13154
rect 18689 13096 18694 13152
rect 18750 13096 23000 13152
rect 18689 13094 23000 13096
rect 18689 13091 18755 13094
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 22520 13064 23000 13094
rect 18270 13023 18590 13024
rect 19517 13018 19583 13021
rect 20437 13018 20503 13021
rect 19517 13016 20503 13018
rect 19517 12960 19522 13016
rect 19578 12960 20442 13016
rect 20498 12960 20503 13016
rect 19517 12958 20503 12960
rect 19517 12955 19583 12958
rect 20437 12955 20503 12958
rect 20294 12882 20300 12884
rect 12893 12880 16682 12882
rect 12893 12824 12898 12880
rect 12954 12824 16682 12880
rect 12893 12822 16682 12824
rect 18048 12822 20300 12882
rect 12893 12819 12959 12822
rect 14038 12684 14044 12748
rect 14108 12746 14114 12748
rect 14365 12746 14431 12749
rect 16389 12746 16455 12749
rect 14108 12744 14431 12746
rect 14108 12688 14370 12744
rect 14426 12688 14431 12744
rect 14108 12686 14431 12688
rect 14108 12684 14114 12686
rect 14365 12683 14431 12686
rect 14598 12744 16455 12746
rect 14598 12688 16394 12744
rect 16450 12688 16455 12744
rect 14598 12686 16455 12688
rect 0 12610 480 12640
rect 3509 12610 3575 12613
rect 0 12608 3575 12610
rect 0 12552 3514 12608
rect 3570 12552 3575 12608
rect 0 12550 3575 12552
rect 0 12520 480 12550
rect 3509 12547 3575 12550
rect 11881 12610 11947 12613
rect 12382 12610 12388 12612
rect 11881 12608 12388 12610
rect 11881 12552 11886 12608
rect 11942 12552 12388 12608
rect 11881 12550 12388 12552
rect 11881 12547 11947 12550
rect 12382 12548 12388 12550
rect 12452 12548 12458 12612
rect 13445 12610 13511 12613
rect 13905 12610 13971 12613
rect 14598 12610 14658 12686
rect 16389 12683 16455 12686
rect 16205 12612 16271 12613
rect 16205 12610 16252 12612
rect 13445 12608 14658 12610
rect 13445 12552 13450 12608
rect 13506 12552 13910 12608
rect 13966 12552 14658 12608
rect 13445 12550 14658 12552
rect 16160 12608 16252 12610
rect 16160 12552 16210 12608
rect 16160 12550 16252 12552
rect 13445 12547 13511 12550
rect 13905 12547 13971 12550
rect 16205 12548 16252 12550
rect 16316 12548 16322 12612
rect 16622 12610 16682 12822
rect 20294 12820 20300 12822
rect 20364 12820 20370 12884
rect 16757 12746 16823 12749
rect 17861 12746 17927 12749
rect 16757 12744 17927 12746
rect 16757 12688 16762 12744
rect 16818 12688 17866 12744
rect 17922 12688 17927 12744
rect 16757 12686 17927 12688
rect 16757 12683 16823 12686
rect 17861 12683 17927 12686
rect 18505 12746 18571 12749
rect 19701 12746 19767 12749
rect 18505 12744 19767 12746
rect 18505 12688 18510 12744
rect 18566 12688 19706 12744
rect 19762 12688 19767 12744
rect 18505 12686 19767 12688
rect 18505 12683 18571 12686
rect 19701 12683 19767 12686
rect 17217 12610 17283 12613
rect 16622 12608 17283 12610
rect 16622 12552 17222 12608
rect 17278 12552 17283 12608
rect 16622 12550 17283 12552
rect 16205 12547 16271 12548
rect 17217 12547 17283 12550
rect 17902 12548 17908 12612
rect 17972 12610 17978 12612
rect 18045 12610 18111 12613
rect 17972 12608 18111 12610
rect 17972 12552 18050 12608
rect 18106 12552 18111 12608
rect 17972 12550 18111 12552
rect 17972 12548 17978 12550
rect 18045 12547 18111 12550
rect 21541 12610 21607 12613
rect 22520 12610 23000 12640
rect 21541 12608 23000 12610
rect 21541 12552 21546 12608
rect 21602 12552 23000 12608
rect 21541 12550 23000 12552
rect 21541 12547 21607 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 22520 12520 23000 12550
rect 14805 12479 15125 12480
rect 10910 12412 10916 12476
rect 10980 12474 10986 12476
rect 14457 12474 14523 12477
rect 10980 12472 14523 12474
rect 10980 12416 14462 12472
rect 14518 12416 14523 12472
rect 10980 12414 14523 12416
rect 10980 12412 10986 12414
rect 11240 12341 11300 12414
rect 14457 12411 14523 12414
rect 16665 12474 16731 12477
rect 17493 12476 17559 12477
rect 16798 12474 16804 12476
rect 16665 12472 16804 12474
rect 16665 12416 16670 12472
rect 16726 12416 16804 12472
rect 16665 12414 16804 12416
rect 16665 12411 16731 12414
rect 16798 12412 16804 12414
rect 16868 12412 16874 12476
rect 17493 12472 17540 12476
rect 17604 12474 17610 12476
rect 17493 12416 17498 12472
rect 17493 12412 17540 12416
rect 17604 12414 17650 12474
rect 17604 12412 17610 12414
rect 17493 12411 17559 12412
rect 7230 12276 7236 12340
rect 7300 12338 7306 12340
rect 7741 12338 7807 12341
rect 7300 12336 7807 12338
rect 7300 12280 7746 12336
rect 7802 12280 7807 12336
rect 7300 12278 7807 12280
rect 7300 12276 7306 12278
rect 7741 12275 7807 12278
rect 11237 12336 11303 12341
rect 19190 12338 19196 12340
rect 11237 12280 11242 12336
rect 11298 12280 11303 12336
rect 11237 12275 11303 12280
rect 11424 12278 19196 12338
rect 0 12202 480 12232
rect 3877 12202 3943 12205
rect 0 12200 3943 12202
rect 0 12144 3882 12200
rect 3938 12144 3943 12200
rect 0 12142 3943 12144
rect 0 12112 480 12142
rect 3877 12139 3943 12142
rect 7373 12202 7439 12205
rect 7833 12202 7899 12205
rect 7373 12200 7899 12202
rect 7373 12144 7378 12200
rect 7434 12144 7838 12200
rect 7894 12144 7899 12200
rect 7373 12142 7899 12144
rect 7373 12139 7439 12142
rect 7833 12139 7899 12142
rect 9121 12202 9187 12205
rect 11424 12202 11484 12278
rect 19190 12276 19196 12278
rect 19260 12276 19266 12340
rect 9121 12200 11484 12202
rect 9121 12144 9126 12200
rect 9182 12144 11484 12200
rect 9121 12142 11484 12144
rect 14089 12202 14155 12205
rect 16849 12204 16915 12205
rect 14222 12202 14228 12204
rect 14089 12200 14228 12202
rect 14089 12144 14094 12200
rect 14150 12144 14228 12200
rect 14089 12142 14228 12144
rect 9121 12139 9187 12142
rect 14089 12139 14155 12142
rect 14222 12140 14228 12142
rect 14292 12140 14298 12204
rect 16798 12140 16804 12204
rect 16868 12202 16915 12204
rect 17309 12202 17375 12205
rect 17534 12202 17540 12204
rect 16868 12200 16960 12202
rect 16910 12144 16960 12200
rect 16868 12142 16960 12144
rect 17309 12200 17540 12202
rect 17309 12144 17314 12200
rect 17370 12144 17540 12200
rect 17309 12142 17540 12144
rect 16868 12140 16915 12142
rect 16849 12139 16915 12140
rect 17309 12139 17375 12142
rect 17534 12140 17540 12142
rect 17604 12140 17610 12204
rect 22520 12202 23000 12232
rect 17910 12142 23000 12202
rect 6729 12066 6795 12069
rect 10409 12068 10475 12069
rect 10174 12066 10180 12068
rect 6729 12064 10180 12066
rect 6729 12008 6734 12064
rect 6790 12008 10180 12064
rect 6729 12006 10180 12008
rect 6729 12003 6795 12006
rect 10174 12004 10180 12006
rect 10244 12004 10250 12068
rect 10358 12004 10364 12068
rect 10428 12066 10475 12068
rect 12341 12066 12407 12069
rect 17769 12066 17835 12069
rect 10428 12064 10520 12066
rect 10470 12008 10520 12064
rect 10428 12006 10520 12008
rect 12341 12064 17835 12066
rect 12341 12008 12346 12064
rect 12402 12008 17774 12064
rect 17830 12008 17835 12064
rect 12341 12006 17835 12008
rect 10428 12004 10475 12006
rect 10409 12003 10475 12004
rect 12341 12003 12407 12006
rect 17769 12003 17835 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 5625 11930 5691 11933
rect 6269 11930 6335 11933
rect 9489 11930 9555 11933
rect 5625 11928 9555 11930
rect 5625 11872 5630 11928
rect 5686 11872 6274 11928
rect 6330 11872 9494 11928
rect 9550 11872 9555 11928
rect 5625 11870 9555 11872
rect 5625 11867 5691 11870
rect 6269 11867 6335 11870
rect 9489 11867 9555 11870
rect 9949 11930 10015 11933
rect 10685 11930 10751 11933
rect 9949 11928 10751 11930
rect 9949 11872 9954 11928
rect 10010 11872 10690 11928
rect 10746 11872 10751 11928
rect 9949 11870 10751 11872
rect 9949 11867 10015 11870
rect 10685 11867 10751 11870
rect 11973 11930 12039 11933
rect 16297 11930 16363 11933
rect 17910 11930 17970 12142
rect 22520 12112 23000 12142
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 11973 11928 16363 11930
rect 11973 11872 11978 11928
rect 12034 11872 16302 11928
rect 16358 11872 16363 11928
rect 11973 11870 16363 11872
rect 11973 11867 12039 11870
rect 16297 11867 16363 11870
rect 16760 11870 17970 11930
rect 16760 11797 16820 11870
rect 7189 11794 7255 11797
rect 7649 11794 7715 11797
rect 7189 11792 7715 11794
rect 7189 11736 7194 11792
rect 7250 11736 7654 11792
rect 7710 11736 7715 11792
rect 7189 11734 7715 11736
rect 7189 11731 7255 11734
rect 7649 11731 7715 11734
rect 10501 11794 10567 11797
rect 14406 11794 14412 11796
rect 10501 11792 14412 11794
rect 10501 11736 10506 11792
rect 10562 11736 14412 11792
rect 10501 11734 14412 11736
rect 10501 11731 10567 11734
rect 14406 11732 14412 11734
rect 14476 11794 14482 11796
rect 16757 11794 16823 11797
rect 14476 11792 16823 11794
rect 14476 11736 16762 11792
rect 16818 11736 16823 11792
rect 14476 11734 16823 11736
rect 14476 11732 14482 11734
rect 16757 11731 16823 11734
rect 18689 11794 18755 11797
rect 20294 11794 20300 11796
rect 18689 11792 20300 11794
rect 18689 11736 18694 11792
rect 18750 11736 20300 11792
rect 18689 11734 20300 11736
rect 18689 11731 18755 11734
rect 20294 11732 20300 11734
rect 20364 11732 20370 11796
rect 0 11658 480 11688
rect 3417 11658 3483 11661
rect 0 11656 3483 11658
rect 0 11600 3422 11656
rect 3478 11600 3483 11656
rect 0 11598 3483 11600
rect 0 11568 480 11598
rect 3417 11595 3483 11598
rect 6913 11658 6979 11661
rect 9121 11658 9187 11661
rect 11329 11658 11395 11661
rect 6913 11656 11395 11658
rect 6913 11600 6918 11656
rect 6974 11600 9126 11656
rect 9182 11600 11334 11656
rect 11390 11600 11395 11656
rect 6913 11598 11395 11600
rect 6913 11595 6979 11598
rect 9121 11595 9187 11598
rect 11329 11595 11395 11598
rect 14181 11658 14247 11661
rect 16665 11658 16731 11661
rect 22520 11658 23000 11688
rect 14181 11656 15578 11658
rect 14181 11600 14186 11656
rect 14242 11600 15578 11656
rect 14181 11598 15578 11600
rect 14181 11595 14247 11598
rect 9673 11522 9739 11525
rect 12341 11522 12407 11525
rect 12566 11522 12572 11524
rect 9673 11520 12572 11522
rect 9673 11464 9678 11520
rect 9734 11464 12346 11520
rect 12402 11464 12572 11520
rect 9673 11462 12572 11464
rect 9673 11459 9739 11462
rect 12341 11459 12407 11462
rect 12566 11460 12572 11462
rect 12636 11460 12642 11524
rect 15518 11522 15578 11598
rect 16665 11656 23000 11658
rect 16665 11600 16670 11656
rect 16726 11600 23000 11656
rect 16665 11598 23000 11600
rect 16665 11595 16731 11598
rect 22520 11568 23000 11598
rect 18689 11522 18755 11525
rect 15518 11520 18755 11522
rect 15518 11464 18694 11520
rect 18750 11464 18755 11520
rect 15518 11462 18755 11464
rect 18689 11459 18755 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 9806 11324 9812 11388
rect 9876 11386 9882 11388
rect 10041 11386 10107 11389
rect 9876 11384 10107 11386
rect 9876 11328 10046 11384
rect 10102 11328 10107 11384
rect 9876 11326 10107 11328
rect 9876 11324 9882 11326
rect 10041 11323 10107 11326
rect 16246 11324 16252 11388
rect 16316 11386 16322 11388
rect 16389 11386 16455 11389
rect 16316 11384 16455 11386
rect 16316 11328 16394 11384
rect 16450 11328 16455 11384
rect 16316 11326 16455 11328
rect 16316 11324 16322 11326
rect 16389 11323 16455 11326
rect 9438 11188 9444 11252
rect 9508 11250 9514 11252
rect 9581 11250 9647 11253
rect 9508 11248 9647 11250
rect 9508 11192 9586 11248
rect 9642 11192 9647 11248
rect 9508 11190 9647 11192
rect 9508 11188 9514 11190
rect 9581 11187 9647 11190
rect 10358 11188 10364 11252
rect 10428 11250 10434 11252
rect 11605 11250 11671 11253
rect 10428 11248 11671 11250
rect 10428 11192 11610 11248
rect 11666 11192 11671 11248
rect 10428 11190 11671 11192
rect 10428 11188 10434 11190
rect 11605 11187 11671 11190
rect 13813 11250 13879 11253
rect 17585 11250 17651 11253
rect 13813 11248 17651 11250
rect 13813 11192 13818 11248
rect 13874 11192 17590 11248
rect 17646 11192 17651 11248
rect 13813 11190 17651 11192
rect 13813 11187 13879 11190
rect 17585 11187 17651 11190
rect 18086 11188 18092 11252
rect 18156 11250 18162 11252
rect 18156 11190 20730 11250
rect 18156 11188 18162 11190
rect 0 11114 480 11144
rect 4061 11114 4127 11117
rect 0 11112 4127 11114
rect 0 11056 4066 11112
rect 4122 11056 4127 11112
rect 0 11054 4127 11056
rect 0 11024 480 11054
rect 4061 11051 4127 11054
rect 9622 11052 9628 11116
rect 9692 11114 9698 11116
rect 10317 11114 10383 11117
rect 9692 11112 10383 11114
rect 9692 11056 10322 11112
rect 10378 11056 10383 11112
rect 9692 11054 10383 11056
rect 9692 11052 9698 11054
rect 10317 11051 10383 11054
rect 11973 11114 12039 11117
rect 12198 11114 12204 11116
rect 11973 11112 12204 11114
rect 11973 11056 11978 11112
rect 12034 11056 12204 11112
rect 11973 11054 12204 11056
rect 11973 11051 12039 11054
rect 12198 11052 12204 11054
rect 12268 11052 12274 11116
rect 14457 11114 14523 11117
rect 18505 11114 18571 11117
rect 14457 11112 18571 11114
rect 14457 11056 14462 11112
rect 14518 11056 18510 11112
rect 18566 11056 18571 11112
rect 14457 11054 18571 11056
rect 14457 11051 14523 11054
rect 18505 11051 18571 11054
rect 20437 11116 20503 11117
rect 20437 11112 20484 11116
rect 20548 11114 20554 11116
rect 20670 11114 20730 11190
rect 22520 11114 23000 11144
rect 20437 11056 20442 11112
rect 20437 11052 20484 11056
rect 20548 11054 20594 11114
rect 20670 11054 23000 11114
rect 20548 11052 20554 11054
rect 20437 11051 20503 11052
rect 22520 11024 23000 11054
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 9213 10844 9279 10845
rect 9213 10842 9260 10844
rect 9168 10840 9260 10842
rect 9168 10784 9218 10840
rect 9168 10782 9260 10784
rect 9213 10780 9260 10782
rect 9324 10780 9330 10844
rect 12157 10842 12223 10845
rect 16297 10842 16363 10845
rect 12157 10840 16363 10842
rect 12157 10784 12162 10840
rect 12218 10784 16302 10840
rect 16358 10784 16363 10840
rect 12157 10782 16363 10784
rect 9213 10779 9279 10780
rect 12157 10779 12223 10782
rect 16297 10779 16363 10782
rect 0 10706 480 10736
rect 3877 10706 3943 10709
rect 0 10704 3943 10706
rect 0 10648 3882 10704
rect 3938 10648 3943 10704
rect 0 10646 3943 10648
rect 0 10616 480 10646
rect 3877 10643 3943 10646
rect 10726 10644 10732 10708
rect 10796 10706 10802 10708
rect 11329 10706 11395 10709
rect 10796 10704 11395 10706
rect 10796 10648 11334 10704
rect 11390 10648 11395 10704
rect 10796 10646 11395 10648
rect 10796 10644 10802 10646
rect 11329 10643 11395 10646
rect 17953 10706 18019 10709
rect 22520 10706 23000 10736
rect 17953 10704 23000 10706
rect 17953 10648 17958 10704
rect 18014 10648 23000 10704
rect 17953 10646 23000 10648
rect 17953 10643 18019 10646
rect 22520 10616 23000 10646
rect 9397 10436 9463 10437
rect 9397 10434 9444 10436
rect 9352 10432 9444 10434
rect 9352 10376 9402 10432
rect 9352 10374 9444 10376
rect 9397 10372 9444 10374
rect 9508 10372 9514 10436
rect 11605 10434 11671 10437
rect 13629 10434 13695 10437
rect 11605 10432 13695 10434
rect 11605 10376 11610 10432
rect 11666 10376 13634 10432
rect 13690 10376 13695 10432
rect 11605 10374 13695 10376
rect 9397 10371 9463 10372
rect 11605 10371 11671 10374
rect 13629 10371 13695 10374
rect 15929 10434 15995 10437
rect 16982 10434 16988 10436
rect 15929 10432 16988 10434
rect 15929 10376 15934 10432
rect 15990 10376 16988 10432
rect 15929 10374 16988 10376
rect 15929 10371 15995 10374
rect 16982 10372 16988 10374
rect 17052 10372 17058 10436
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 10777 10298 10843 10301
rect 12525 10298 12591 10301
rect 10777 10296 12591 10298
rect 10777 10240 10782 10296
rect 10838 10240 12530 10296
rect 12586 10240 12591 10296
rect 10777 10238 12591 10240
rect 10777 10235 10843 10238
rect 12525 10235 12591 10238
rect 19190 10236 19196 10300
rect 19260 10298 19266 10300
rect 20621 10298 20687 10301
rect 19260 10296 20687 10298
rect 19260 10240 20626 10296
rect 20682 10240 20687 10296
rect 19260 10238 20687 10240
rect 19260 10236 19266 10238
rect 20621 10235 20687 10238
rect 0 10162 480 10192
rect 3877 10162 3943 10165
rect 0 10160 3943 10162
rect 0 10104 3882 10160
rect 3938 10104 3943 10160
rect 0 10102 3943 10104
rect 0 10072 480 10102
rect 3877 10099 3943 10102
rect 10542 10100 10548 10164
rect 10612 10162 10618 10164
rect 10777 10162 10843 10165
rect 10612 10160 10843 10162
rect 10612 10104 10782 10160
rect 10838 10104 10843 10160
rect 10612 10102 10843 10104
rect 10612 10100 10618 10102
rect 10777 10099 10843 10102
rect 10961 10162 11027 10165
rect 11145 10162 11211 10165
rect 10961 10160 11211 10162
rect 10961 10104 10966 10160
rect 11022 10104 11150 10160
rect 11206 10104 11211 10160
rect 10961 10102 11211 10104
rect 10961 10099 11027 10102
rect 11145 10099 11211 10102
rect 22369 10162 22435 10165
rect 22520 10162 23000 10192
rect 22369 10160 23000 10162
rect 22369 10104 22374 10160
rect 22430 10104 23000 10160
rect 22369 10102 23000 10104
rect 22369 10099 22435 10102
rect 22520 10072 23000 10102
rect 13670 9964 13676 10028
rect 13740 10026 13746 10028
rect 14181 10026 14247 10029
rect 13740 10024 14247 10026
rect 13740 9968 14186 10024
rect 14242 9968 14247 10024
rect 13740 9966 14247 9968
rect 13740 9964 13746 9966
rect 14181 9963 14247 9966
rect 14917 10026 14983 10029
rect 14917 10024 19626 10026
rect 14917 9968 14922 10024
rect 14978 9968 19626 10024
rect 14917 9966 19626 9968
rect 14917 9963 14983 9966
rect 8385 9892 8451 9893
rect 8334 9890 8340 9892
rect 8294 9830 8340 9890
rect 8404 9888 8451 9892
rect 19566 9890 19626 9966
rect 19742 9964 19748 10028
rect 19812 10026 19818 10028
rect 20069 10026 20135 10029
rect 19812 10024 20135 10026
rect 19812 9968 20074 10024
rect 20130 9968 20135 10024
rect 19812 9966 20135 9968
rect 19812 9964 19818 9966
rect 20069 9963 20135 9966
rect 22369 9890 22435 9893
rect 8446 9832 8451 9888
rect 8334 9828 8340 9830
rect 8404 9828 8451 9832
rect 8385 9827 8451 9828
rect 11792 9830 18108 9890
rect 19566 9888 22435 9890
rect 19566 9832 22374 9888
rect 22430 9832 22435 9888
rect 19566 9830 22435 9832
rect 4409 9824 4729 9825
rect 0 9754 480 9784
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 4061 9754 4127 9757
rect 7465 9756 7531 9757
rect 0 9752 4127 9754
rect 0 9696 4066 9752
rect 4122 9696 4127 9752
rect 0 9694 4127 9696
rect 0 9664 480 9694
rect 4061 9691 4127 9694
rect 7414 9692 7420 9756
rect 7484 9754 7531 9756
rect 7484 9752 7576 9754
rect 7526 9696 7576 9752
rect 7484 9694 7576 9696
rect 7484 9692 7531 9694
rect 7465 9691 7531 9692
rect 3233 9618 3299 9621
rect 5717 9618 5783 9621
rect 3233 9616 5783 9618
rect 3233 9560 3238 9616
rect 3294 9560 5722 9616
rect 5778 9560 5783 9616
rect 3233 9558 5783 9560
rect 3233 9555 3299 9558
rect 5717 9555 5783 9558
rect 8385 9618 8451 9621
rect 11792 9618 11852 9830
rect 12525 9754 12591 9757
rect 14365 9754 14431 9757
rect 12525 9752 14431 9754
rect 12525 9696 12530 9752
rect 12586 9696 14370 9752
rect 14426 9696 14431 9752
rect 12525 9694 14431 9696
rect 12525 9691 12591 9694
rect 14365 9691 14431 9694
rect 8385 9616 11852 9618
rect 8385 9560 8390 9616
rect 8446 9560 11852 9616
rect 8385 9558 11852 9560
rect 14273 9616 14339 9621
rect 14273 9560 14278 9616
rect 14334 9560 14339 9616
rect 8385 9555 8451 9558
rect 14273 9555 14339 9560
rect 14549 9618 14615 9621
rect 14733 9618 14799 9621
rect 14549 9616 16820 9618
rect 14549 9560 14554 9616
rect 14610 9560 14738 9616
rect 14794 9560 16820 9616
rect 14549 9558 16820 9560
rect 14549 9555 14615 9558
rect 14733 9555 14799 9558
rect 6913 9482 6979 9485
rect 8518 9482 8524 9484
rect 6913 9480 8524 9482
rect 6913 9424 6918 9480
rect 6974 9424 8524 9480
rect 6913 9422 8524 9424
rect 6913 9419 6979 9422
rect 8518 9420 8524 9422
rect 8588 9420 8594 9484
rect 8702 9420 8708 9484
rect 8772 9482 8778 9484
rect 11697 9482 11763 9485
rect 8772 9480 11763 9482
rect 8772 9424 11702 9480
rect 11758 9424 11763 9480
rect 8772 9422 11763 9424
rect 14276 9482 14336 9555
rect 16481 9484 16547 9485
rect 14276 9422 15256 9482
rect 8772 9420 8778 9422
rect 11697 9419 11763 9422
rect 8293 9346 8359 9349
rect 8518 9346 8524 9348
rect 8293 9344 8524 9346
rect 8293 9288 8298 9344
rect 8354 9288 8524 9344
rect 8293 9286 8524 9288
rect 8293 9283 8359 9286
rect 8518 9284 8524 9286
rect 8588 9284 8594 9348
rect 8661 9346 8727 9349
rect 10225 9346 10291 9349
rect 10961 9346 11027 9349
rect 11881 9348 11947 9349
rect 11830 9346 11836 9348
rect 8661 9344 10291 9346
rect 8661 9288 8666 9344
rect 8722 9288 10230 9344
rect 10286 9288 10291 9344
rect 8661 9286 10291 9288
rect 8661 9283 8727 9286
rect 10225 9283 10291 9286
rect 10366 9344 11027 9346
rect 10366 9288 10966 9344
rect 11022 9288 11027 9344
rect 10366 9286 11027 9288
rect 11790 9286 11836 9346
rect 11900 9344 11947 9348
rect 14549 9346 14615 9349
rect 11942 9288 11947 9344
rect 7874 9280 8194 9281
rect 0 9210 480 9240
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 8385 9212 8451 9213
rect 0 9150 2836 9210
rect 0 9120 480 9150
rect 2776 9074 2836 9150
rect 8334 9148 8340 9212
rect 8404 9210 8451 9212
rect 8404 9208 8496 9210
rect 8446 9152 8496 9208
rect 8404 9150 8496 9152
rect 8404 9148 8451 9150
rect 8385 9147 8451 9148
rect 10366 9076 10426 9286
rect 10961 9283 11027 9286
rect 11830 9284 11836 9286
rect 11900 9284 11947 9288
rect 11881 9283 11947 9284
rect 12160 9344 14615 9346
rect 12160 9288 14554 9344
rect 14610 9288 14615 9344
rect 12160 9286 14615 9288
rect 15196 9346 15256 9422
rect 16430 9420 16436 9484
rect 16500 9482 16547 9484
rect 16760 9482 16820 9558
rect 17166 9556 17172 9620
rect 17236 9618 17242 9620
rect 17769 9618 17835 9621
rect 17236 9616 17835 9618
rect 17236 9560 17774 9616
rect 17830 9560 17835 9616
rect 17236 9558 17835 9560
rect 18048 9618 18108 9830
rect 22369 9827 22435 9830
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 18822 9692 18828 9756
rect 18892 9754 18898 9756
rect 22520 9754 23000 9784
rect 18892 9694 23000 9754
rect 18892 9692 18898 9694
rect 18830 9618 18890 9692
rect 22520 9664 23000 9694
rect 18048 9558 18890 9618
rect 17236 9556 17242 9558
rect 17769 9555 17835 9558
rect 19374 9556 19380 9620
rect 19444 9618 19450 9620
rect 19701 9618 19767 9621
rect 20069 9620 20135 9621
rect 20069 9618 20116 9620
rect 19444 9616 19767 9618
rect 19444 9560 19706 9616
rect 19762 9560 19767 9616
rect 19444 9558 19767 9560
rect 20024 9616 20116 9618
rect 20024 9560 20074 9616
rect 20024 9558 20116 9560
rect 19444 9556 19450 9558
rect 19701 9555 19767 9558
rect 20069 9556 20116 9558
rect 20180 9556 20186 9620
rect 20069 9555 20135 9556
rect 18873 9482 18939 9485
rect 16500 9480 16592 9482
rect 16542 9424 16592 9480
rect 16500 9422 16592 9424
rect 16760 9480 18939 9482
rect 16760 9424 18878 9480
rect 18934 9424 18939 9480
rect 16760 9422 18939 9424
rect 16500 9420 16547 9422
rect 16481 9419 16547 9420
rect 18873 9419 18939 9422
rect 19006 9420 19012 9484
rect 19076 9482 19082 9484
rect 19333 9482 19399 9485
rect 19076 9480 19399 9482
rect 19076 9424 19338 9480
rect 19394 9424 19399 9480
rect 19076 9422 19399 9424
rect 19076 9420 19082 9422
rect 19333 9419 19399 9422
rect 18505 9346 18571 9349
rect 15196 9344 18571 9346
rect 15196 9288 18510 9344
rect 18566 9288 18571 9344
rect 15196 9286 18571 9288
rect 11789 9210 11855 9213
rect 12160 9210 12220 9286
rect 14549 9283 14615 9286
rect 18505 9283 18571 9286
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 11789 9208 12220 9210
rect 11789 9152 11794 9208
rect 11850 9152 12220 9208
rect 11789 9150 12220 9152
rect 15285 9210 15351 9213
rect 15510 9210 15516 9212
rect 15285 9208 15516 9210
rect 15285 9152 15290 9208
rect 15346 9152 15516 9208
rect 15285 9150 15516 9152
rect 11789 9147 11855 9150
rect 15285 9147 15351 9150
rect 15510 9148 15516 9150
rect 15580 9148 15586 9212
rect 19977 9210 20043 9213
rect 22520 9210 23000 9240
rect 19977 9208 23000 9210
rect 19977 9152 19982 9208
rect 20038 9152 23000 9208
rect 19977 9150 23000 9152
rect 19977 9147 20043 9150
rect 22520 9120 23000 9150
rect 10358 9074 10364 9076
rect 2776 9014 10364 9074
rect 10358 9012 10364 9014
rect 10428 9012 10434 9076
rect 13353 9072 13419 9077
rect 13353 9016 13358 9072
rect 13414 9016 13419 9072
rect 13353 9011 13419 9016
rect 13813 9074 13879 9077
rect 18505 9074 18571 9077
rect 13813 9072 18571 9074
rect 13813 9016 13818 9072
rect 13874 9016 18510 9072
rect 18566 9016 18571 9072
rect 13813 9014 18571 9016
rect 13813 9011 13879 9014
rect 18505 9011 18571 9014
rect 19198 9014 20178 9074
rect 6545 8938 6611 8941
rect 13356 8938 13416 9011
rect 6545 8936 13416 8938
rect 6545 8880 6550 8936
rect 6606 8880 13416 8936
rect 6545 8878 13416 8880
rect 6545 8875 6611 8878
rect 0 8802 480 8832
rect 4245 8802 4311 8805
rect 0 8800 4311 8802
rect 0 8744 4250 8800
rect 4306 8744 4311 8800
rect 0 8742 4311 8744
rect 0 8712 480 8742
rect 4245 8739 4311 8742
rect 5901 8802 5967 8805
rect 8017 8802 8083 8805
rect 9806 8802 9812 8804
rect 5901 8800 9812 8802
rect 5901 8744 5906 8800
rect 5962 8744 8022 8800
rect 8078 8744 9812 8800
rect 5901 8742 9812 8744
rect 5901 8739 5967 8742
rect 8017 8739 8083 8742
rect 9806 8740 9812 8742
rect 9876 8740 9882 8804
rect 13356 8802 13416 8878
rect 16430 8876 16436 8940
rect 16500 8938 16506 8940
rect 19198 8938 19258 9014
rect 16500 8878 19258 8938
rect 16500 8876 16506 8878
rect 17401 8802 17467 8805
rect 13356 8800 17467 8802
rect 13356 8744 17406 8800
rect 17462 8744 17467 8800
rect 13356 8742 17467 8744
rect 20118 8802 20178 9014
rect 22520 8802 23000 8832
rect 20118 8742 23000 8802
rect 17401 8739 17467 8742
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 22520 8712 23000 8742
rect 18270 8671 18590 8672
rect 6177 8666 6243 8669
rect 10593 8666 10659 8669
rect 17677 8666 17743 8669
rect 6177 8664 10659 8666
rect 6177 8608 6182 8664
rect 6238 8608 10598 8664
rect 10654 8608 10659 8664
rect 6177 8606 10659 8608
rect 6177 8603 6243 8606
rect 10593 8603 10659 8606
rect 11884 8664 17743 8666
rect 11884 8608 17682 8664
rect 17738 8608 17743 8664
rect 11884 8606 17743 8608
rect 5165 8530 5231 8533
rect 7189 8530 7255 8533
rect 8702 8530 8708 8532
rect 5165 8528 8708 8530
rect 5165 8472 5170 8528
rect 5226 8472 7194 8528
rect 7250 8472 8708 8528
rect 5165 8470 8708 8472
rect 5165 8467 5231 8470
rect 7189 8467 7255 8470
rect 8702 8468 8708 8470
rect 8772 8468 8778 8532
rect 9029 8530 9095 8533
rect 9397 8530 9463 8533
rect 9029 8528 9463 8530
rect 9029 8472 9034 8528
rect 9090 8472 9402 8528
rect 9458 8472 9463 8528
rect 9029 8470 9463 8472
rect 9029 8467 9095 8470
rect 9397 8467 9463 8470
rect 10685 8530 10751 8533
rect 11884 8530 11944 8606
rect 17677 8603 17743 8606
rect 10685 8528 11944 8530
rect 10685 8472 10690 8528
rect 10746 8472 11944 8528
rect 10685 8470 11944 8472
rect 15009 8530 15075 8533
rect 15377 8530 15443 8533
rect 15745 8530 15811 8533
rect 19149 8530 19215 8533
rect 15009 8528 19215 8530
rect 15009 8472 15014 8528
rect 15070 8472 15382 8528
rect 15438 8472 15750 8528
rect 15806 8472 19154 8528
rect 19210 8472 19215 8528
rect 15009 8470 19215 8472
rect 10685 8467 10751 8470
rect 15009 8467 15075 8470
rect 15377 8467 15443 8470
rect 15745 8467 15811 8470
rect 19149 8467 19215 8470
rect 19333 8530 19399 8533
rect 20621 8530 20687 8533
rect 19333 8528 20687 8530
rect 19333 8472 19338 8528
rect 19394 8472 20626 8528
rect 20682 8472 20687 8528
rect 19333 8470 20687 8472
rect 19333 8467 19399 8470
rect 20621 8467 20687 8470
rect 8518 8332 8524 8396
rect 8588 8394 8594 8396
rect 9765 8394 9831 8397
rect 8588 8392 9831 8394
rect 8588 8336 9770 8392
rect 9826 8336 9831 8392
rect 8588 8334 9831 8336
rect 8588 8332 8594 8334
rect 9765 8331 9831 8334
rect 10041 8394 10107 8397
rect 11329 8394 11395 8397
rect 15929 8394 15995 8397
rect 10041 8392 11395 8394
rect 10041 8336 10046 8392
rect 10102 8336 11334 8392
rect 11390 8336 11395 8392
rect 10041 8334 11395 8336
rect 10041 8331 10107 8334
rect 11329 8331 11395 8334
rect 11470 8392 15995 8394
rect 11470 8336 15934 8392
rect 15990 8336 15995 8392
rect 11470 8334 15995 8336
rect 0 8258 480 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 480 8198
rect 4061 8195 4127 8198
rect 5809 8258 5875 8261
rect 7741 8258 7807 8261
rect 5809 8256 7807 8258
rect 5809 8200 5814 8256
rect 5870 8200 7746 8256
rect 7802 8200 7807 8256
rect 5809 8198 7807 8200
rect 5809 8195 5875 8198
rect 7741 8195 7807 8198
rect 9765 8258 9831 8261
rect 11470 8258 11530 8334
rect 15929 8331 15995 8334
rect 17902 8332 17908 8396
rect 17972 8394 17978 8396
rect 18321 8394 18387 8397
rect 17972 8392 18387 8394
rect 17972 8336 18326 8392
rect 18382 8336 18387 8392
rect 17972 8334 18387 8336
rect 17972 8332 17978 8334
rect 18321 8331 18387 8334
rect 18597 8394 18663 8397
rect 19190 8394 19196 8396
rect 18597 8392 19196 8394
rect 18597 8336 18602 8392
rect 18658 8336 19196 8392
rect 18597 8334 19196 8336
rect 18597 8331 18663 8334
rect 19190 8332 19196 8334
rect 19260 8332 19266 8396
rect 20110 8332 20116 8396
rect 20180 8394 20186 8396
rect 20345 8394 20411 8397
rect 20180 8392 20411 8394
rect 20180 8336 20350 8392
rect 20406 8336 20411 8392
rect 20180 8334 20411 8336
rect 20180 8332 20186 8334
rect 20345 8331 20411 8334
rect 9765 8256 11530 8258
rect 9765 8200 9770 8256
rect 9826 8200 11530 8256
rect 9765 8198 11530 8200
rect 15745 8258 15811 8261
rect 22520 8258 23000 8288
rect 15745 8256 23000 8258
rect 15745 8200 15750 8256
rect 15806 8200 23000 8256
rect 15745 8198 23000 8200
rect 9765 8195 9831 8198
rect 15745 8195 15811 8198
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 22520 8168 23000 8198
rect 14805 8127 15125 8128
rect 10501 8122 10567 8125
rect 13854 8122 13860 8124
rect 10501 8120 13860 8122
rect 10501 8064 10506 8120
rect 10562 8064 13860 8120
rect 10501 8062 13860 8064
rect 10501 8059 10567 8062
rect 13854 8060 13860 8062
rect 13924 8060 13930 8124
rect 19333 8122 19399 8125
rect 21725 8122 21791 8125
rect 19333 8120 21791 8122
rect 19333 8064 19338 8120
rect 19394 8064 21730 8120
rect 21786 8064 21791 8120
rect 19333 8062 21791 8064
rect 19333 8059 19399 8062
rect 21725 8059 21791 8062
rect 5349 7986 5415 7989
rect 15469 7986 15535 7989
rect 5349 7984 15535 7986
rect 5349 7928 5354 7984
rect 5410 7928 15474 7984
rect 15530 7928 15535 7984
rect 5349 7926 15535 7928
rect 5349 7923 5415 7926
rect 15469 7923 15535 7926
rect 0 7850 480 7880
rect 4061 7850 4127 7853
rect 0 7848 4127 7850
rect 0 7792 4066 7848
rect 4122 7792 4127 7848
rect 0 7790 4127 7792
rect 0 7760 480 7790
rect 4061 7787 4127 7790
rect 7189 7850 7255 7853
rect 13261 7850 13327 7853
rect 7189 7848 13327 7850
rect 7189 7792 7194 7848
rect 7250 7792 13266 7848
rect 13322 7792 13327 7848
rect 7189 7790 13327 7792
rect 7189 7787 7255 7790
rect 13261 7787 13327 7790
rect 17401 7850 17467 7853
rect 17585 7850 17651 7853
rect 17401 7848 17651 7850
rect 17401 7792 17406 7848
rect 17462 7792 17590 7848
rect 17646 7792 17651 7848
rect 17401 7790 17651 7792
rect 17401 7787 17467 7790
rect 17585 7787 17651 7790
rect 17953 7850 18019 7853
rect 22520 7850 23000 7880
rect 17953 7848 23000 7850
rect 17953 7792 17958 7848
rect 18014 7792 23000 7848
rect 17953 7790 23000 7792
rect 17953 7787 18019 7790
rect 22520 7760 23000 7790
rect 5073 7714 5139 7717
rect 7833 7714 7899 7717
rect 9029 7716 9095 7717
rect 9029 7714 9076 7716
rect 5073 7712 7899 7714
rect 5073 7656 5078 7712
rect 5134 7656 7838 7712
rect 7894 7656 7899 7712
rect 5073 7654 7899 7656
rect 8948 7712 9076 7714
rect 9140 7714 9146 7716
rect 10041 7714 10107 7717
rect 9140 7712 10107 7714
rect 8948 7656 9034 7712
rect 9140 7656 10046 7712
rect 10102 7656 10107 7712
rect 8948 7654 9076 7656
rect 5073 7651 5139 7654
rect 7833 7651 7899 7654
rect 9029 7652 9076 7654
rect 9140 7654 10107 7656
rect 9140 7652 9146 7654
rect 9029 7651 9095 7652
rect 10041 7651 10107 7654
rect 10358 7652 10364 7716
rect 10428 7714 10434 7716
rect 10501 7714 10567 7717
rect 10428 7712 10567 7714
rect 10428 7656 10506 7712
rect 10562 7656 10567 7712
rect 10428 7654 10567 7656
rect 10428 7652 10434 7654
rect 10501 7651 10567 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 9673 7578 9739 7581
rect 10041 7578 10107 7581
rect 17953 7578 18019 7581
rect 9673 7576 10107 7578
rect 9673 7520 9678 7576
rect 9734 7520 10046 7576
rect 10102 7520 10107 7576
rect 9673 7518 10107 7520
rect 9673 7515 9739 7518
rect 10041 7515 10107 7518
rect 11838 7576 18019 7578
rect 11838 7520 17958 7576
rect 18014 7520 18019 7576
rect 11838 7518 18019 7520
rect 8477 7442 8543 7445
rect 8845 7442 8911 7445
rect 11838 7442 11898 7518
rect 17953 7515 18019 7518
rect 8477 7440 8770 7442
rect 8477 7384 8482 7440
rect 8538 7384 8770 7440
rect 8477 7382 8770 7384
rect 8477 7379 8543 7382
rect 0 7306 480 7336
rect 3969 7306 4035 7309
rect 0 7304 4035 7306
rect 0 7248 3974 7304
rect 4030 7248 4035 7304
rect 0 7246 4035 7248
rect 0 7216 480 7246
rect 3969 7243 4035 7246
rect 7741 7306 7807 7309
rect 8710 7306 8770 7382
rect 8845 7440 11898 7442
rect 8845 7384 8850 7440
rect 8906 7384 11898 7440
rect 8845 7382 11898 7384
rect 12157 7442 12223 7445
rect 18505 7442 18571 7445
rect 19057 7442 19123 7445
rect 12157 7440 17556 7442
rect 12157 7384 12162 7440
rect 12218 7384 17556 7440
rect 12157 7382 17556 7384
rect 8845 7379 8911 7382
rect 12157 7379 12223 7382
rect 8937 7306 9003 7309
rect 9765 7306 9831 7309
rect 15561 7306 15627 7309
rect 7741 7304 8586 7306
rect 7741 7248 7746 7304
rect 7802 7248 8586 7304
rect 7741 7246 8586 7248
rect 8710 7304 9690 7306
rect 8710 7248 8942 7304
rect 8998 7248 9690 7304
rect 8710 7246 9690 7248
rect 7741 7243 7807 7246
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 8526 7034 8586 7246
rect 8937 7243 9003 7246
rect 9630 7170 9690 7246
rect 9765 7304 15627 7306
rect 9765 7248 9770 7304
rect 9826 7248 15566 7304
rect 15622 7248 15627 7304
rect 9765 7246 15627 7248
rect 17496 7306 17556 7382
rect 18505 7440 19123 7442
rect 18505 7384 18510 7440
rect 18566 7384 19062 7440
rect 19118 7384 19123 7440
rect 18505 7382 19123 7384
rect 18505 7379 18571 7382
rect 19057 7379 19123 7382
rect 22520 7306 23000 7336
rect 17496 7246 23000 7306
rect 9765 7243 9831 7246
rect 15561 7243 15627 7246
rect 22520 7216 23000 7246
rect 12249 7170 12315 7173
rect 9630 7168 12315 7170
rect 9630 7112 12254 7168
rect 12310 7112 12315 7168
rect 9630 7110 12315 7112
rect 12249 7107 12315 7110
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 12157 7034 12223 7037
rect 8526 7032 12223 7034
rect 8526 6976 12162 7032
rect 12218 6976 12223 7032
rect 8526 6974 12223 6976
rect 12157 6971 12223 6974
rect 0 6898 480 6928
rect 9673 6898 9739 6901
rect 17033 6898 17099 6901
rect 0 6896 9739 6898
rect 0 6840 9678 6896
rect 9734 6840 9739 6896
rect 0 6838 9739 6840
rect 0 6808 480 6838
rect 9673 6835 9739 6838
rect 13310 6896 17099 6898
rect 13310 6840 17038 6896
rect 17094 6840 17099 6896
rect 13310 6838 17099 6840
rect 6177 6762 6243 6765
rect 13310 6762 13370 6838
rect 17033 6835 17099 6838
rect 17953 6898 18019 6901
rect 22520 6898 23000 6928
rect 17953 6896 23000 6898
rect 17953 6840 17958 6896
rect 18014 6840 23000 6896
rect 17953 6838 23000 6840
rect 17953 6835 18019 6838
rect 22520 6808 23000 6838
rect 6177 6760 13370 6762
rect 6177 6704 6182 6760
rect 6238 6704 13370 6760
rect 6177 6702 13370 6704
rect 15653 6762 15719 6765
rect 15929 6762 15995 6765
rect 15653 6760 15995 6762
rect 15653 6704 15658 6760
rect 15714 6704 15934 6760
rect 15990 6704 15995 6760
rect 15653 6702 15995 6704
rect 6177 6699 6243 6702
rect 15653 6699 15719 6702
rect 15929 6699 15995 6702
rect 15653 6626 15719 6629
rect 16757 6626 16823 6629
rect 15653 6624 16823 6626
rect 15653 6568 15658 6624
rect 15714 6568 16762 6624
rect 16818 6568 16823 6624
rect 15653 6566 16823 6568
rect 15653 6563 15719 6566
rect 16757 6563 16823 6566
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6354 480 6384
rect 3969 6354 4035 6357
rect 0 6352 4035 6354
rect 0 6296 3974 6352
rect 4030 6296 4035 6352
rect 0 6294 4035 6296
rect 0 6264 480 6294
rect 3969 6291 4035 6294
rect 4889 6354 4955 6357
rect 8661 6354 8727 6357
rect 4889 6352 8727 6354
rect 4889 6296 4894 6352
rect 4950 6296 8666 6352
rect 8722 6296 8727 6352
rect 4889 6294 8727 6296
rect 4889 6291 4955 6294
rect 8661 6291 8727 6294
rect 12014 6292 12020 6356
rect 12084 6354 12090 6356
rect 13077 6354 13143 6357
rect 12084 6352 13143 6354
rect 12084 6296 13082 6352
rect 13138 6296 13143 6352
rect 12084 6294 13143 6296
rect 12084 6292 12090 6294
rect 13077 6291 13143 6294
rect 15561 6354 15627 6357
rect 17217 6354 17283 6357
rect 15561 6352 17283 6354
rect 15561 6296 15566 6352
rect 15622 6296 17222 6352
rect 17278 6296 17283 6352
rect 15561 6294 17283 6296
rect 15561 6291 15627 6294
rect 17217 6291 17283 6294
rect 17493 6354 17559 6357
rect 22520 6354 23000 6384
rect 17493 6352 23000 6354
rect 17493 6296 17498 6352
rect 17554 6296 23000 6352
rect 17493 6294 23000 6296
rect 17493 6291 17559 6294
rect 22520 6264 23000 6294
rect 5993 6218 6059 6221
rect 10777 6218 10843 6221
rect 13721 6218 13787 6221
rect 5993 6216 13787 6218
rect 5993 6160 5998 6216
rect 6054 6160 10782 6216
rect 10838 6160 13726 6216
rect 13782 6160 13787 6216
rect 5993 6158 13787 6160
rect 5993 6155 6059 6158
rect 10777 6155 10843 6158
rect 13721 6155 13787 6158
rect 13854 6156 13860 6220
rect 13924 6218 13930 6220
rect 13924 6158 16682 6218
rect 13924 6156 13930 6158
rect 16622 6085 16682 6158
rect 8661 6082 8727 6085
rect 9489 6082 9555 6085
rect 8661 6080 9555 6082
rect 8661 6024 8666 6080
rect 8722 6024 9494 6080
rect 9550 6024 9555 6080
rect 8661 6022 9555 6024
rect 16622 6080 16731 6085
rect 16622 6024 16670 6080
rect 16726 6024 16731 6080
rect 16622 6022 16731 6024
rect 8661 6019 8727 6022
rect 9489 6019 9555 6022
rect 16665 6019 16731 6022
rect 17953 6082 18019 6085
rect 22369 6082 22435 6085
rect 17953 6080 22435 6082
rect 17953 6024 17958 6080
rect 18014 6024 22374 6080
rect 22430 6024 22435 6080
rect 17953 6022 22435 6024
rect 17953 6019 18019 6022
rect 22369 6019 22435 6022
rect 7874 6016 8194 6017
rect 0 5946 480 5976
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 12065 5946 12131 5949
rect 12525 5946 12591 5949
rect 22520 5946 23000 5976
rect 0 5886 5688 5946
rect 0 5856 480 5886
rect 5628 5674 5688 5886
rect 12065 5944 12591 5946
rect 12065 5888 12070 5944
rect 12126 5888 12530 5944
rect 12586 5888 12591 5944
rect 12065 5886 12591 5888
rect 12065 5883 12131 5886
rect 12525 5883 12591 5886
rect 19566 5886 23000 5946
rect 5809 5810 5875 5813
rect 7925 5810 7991 5813
rect 5809 5808 7991 5810
rect 5809 5752 5814 5808
rect 5870 5752 7930 5808
rect 7986 5752 7991 5808
rect 5809 5750 7991 5752
rect 5809 5747 5875 5750
rect 7925 5747 7991 5750
rect 8293 5810 8359 5813
rect 10225 5810 10291 5813
rect 8293 5808 10291 5810
rect 8293 5752 8298 5808
rect 8354 5752 10230 5808
rect 10286 5752 10291 5808
rect 8293 5750 10291 5752
rect 8293 5747 8359 5750
rect 10225 5747 10291 5750
rect 13813 5810 13879 5813
rect 19333 5812 19399 5813
rect 19333 5810 19380 5812
rect 13813 5808 19074 5810
rect 13813 5752 13818 5808
rect 13874 5752 19074 5808
rect 13813 5750 19074 5752
rect 19288 5808 19380 5810
rect 19288 5752 19338 5808
rect 19288 5750 19380 5752
rect 13813 5747 13879 5750
rect 7598 5674 7604 5676
rect 5628 5614 7604 5674
rect 7598 5612 7604 5614
rect 7668 5674 7674 5676
rect 12065 5674 12131 5677
rect 12617 5674 12683 5677
rect 7668 5614 11162 5674
rect 7668 5612 7674 5614
rect 7741 5538 7807 5541
rect 8845 5538 8911 5541
rect 9121 5538 9187 5541
rect 7741 5536 9187 5538
rect 7741 5480 7746 5536
rect 7802 5480 8850 5536
rect 8906 5480 9126 5536
rect 9182 5480 9187 5536
rect 7741 5478 9187 5480
rect 7741 5475 7807 5478
rect 8845 5475 8911 5478
rect 9121 5475 9187 5478
rect 4409 5472 4729 5473
rect 0 5402 480 5432
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 7373 5402 7439 5405
rect 10593 5402 10659 5405
rect 0 5342 4170 5402
rect 0 5312 480 5342
rect 4110 5266 4170 5342
rect 7373 5400 10659 5402
rect 7373 5344 7378 5400
rect 7434 5344 10598 5400
rect 10654 5344 10659 5400
rect 7373 5342 10659 5344
rect 7373 5339 7439 5342
rect 10593 5339 10659 5342
rect 7189 5266 7255 5269
rect 4110 5264 7255 5266
rect 4110 5208 7194 5264
rect 7250 5208 7255 5264
rect 4110 5206 7255 5208
rect 7189 5203 7255 5206
rect 7465 5266 7531 5269
rect 8385 5266 8451 5269
rect 7465 5264 8451 5266
rect 7465 5208 7470 5264
rect 7526 5208 8390 5264
rect 8446 5208 8451 5264
rect 7465 5206 8451 5208
rect 11102 5266 11162 5614
rect 12065 5672 12683 5674
rect 12065 5616 12070 5672
rect 12126 5616 12622 5672
rect 12678 5616 12683 5672
rect 12065 5614 12683 5616
rect 12065 5611 12131 5614
rect 12617 5611 12683 5614
rect 14181 5674 14247 5677
rect 17493 5674 17559 5677
rect 19014 5674 19074 5750
rect 19333 5748 19380 5750
rect 19444 5748 19450 5812
rect 19333 5747 19399 5748
rect 19566 5674 19626 5886
rect 22520 5856 23000 5886
rect 14181 5672 17559 5674
rect 14181 5616 14186 5672
rect 14242 5616 17498 5672
rect 17554 5616 17559 5672
rect 14181 5614 17559 5616
rect 14181 5611 14247 5614
rect 17493 5611 17559 5614
rect 18094 5614 18844 5674
rect 19014 5614 19626 5674
rect 12198 5476 12204 5540
rect 12268 5538 12274 5540
rect 18094 5538 18154 5614
rect 12268 5478 18154 5538
rect 18784 5538 18844 5614
rect 20161 5538 20227 5541
rect 18784 5536 20227 5538
rect 18784 5480 20166 5536
rect 20222 5480 20227 5536
rect 18784 5478 20227 5480
rect 12268 5476 12274 5478
rect 20161 5475 20227 5478
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 22520 5402 23000 5432
rect 22326 5342 23000 5402
rect 11329 5266 11395 5269
rect 17902 5266 17908 5268
rect 11102 5264 11395 5266
rect 11102 5208 11334 5264
rect 11390 5208 11395 5264
rect 11102 5206 11395 5208
rect 7465 5203 7531 5206
rect 8385 5203 8451 5206
rect 11329 5203 11395 5206
rect 14414 5206 17908 5266
rect 3969 5130 4035 5133
rect 12014 5130 12020 5132
rect 3969 5128 12020 5130
rect 3969 5072 3974 5128
rect 4030 5072 12020 5128
rect 3969 5070 12020 5072
rect 3969 5067 4035 5070
rect 12014 5068 12020 5070
rect 12084 5068 12090 5132
rect 0 4994 480 5024
rect 4061 4994 4127 4997
rect 0 4992 4127 4994
rect 0 4936 4066 4992
rect 4122 4936 4127 4992
rect 0 4934 4127 4936
rect 0 4904 480 4934
rect 4061 4931 4127 4934
rect 8385 4994 8451 4997
rect 8569 4994 8635 4997
rect 8385 4992 8635 4994
rect 8385 4936 8390 4992
rect 8446 4936 8574 4992
rect 8630 4936 8635 4992
rect 8385 4934 8635 4936
rect 8385 4931 8451 4934
rect 8569 4931 8635 4934
rect 9397 4994 9463 4997
rect 14414 4994 14474 5206
rect 17902 5204 17908 5206
rect 17972 5204 17978 5268
rect 20529 5266 20595 5269
rect 22326 5266 22386 5342
rect 22520 5312 23000 5342
rect 20529 5264 22386 5266
rect 20529 5208 20534 5264
rect 20590 5208 22386 5264
rect 20529 5206 22386 5208
rect 20529 5203 20595 5206
rect 18505 5130 18571 5133
rect 9397 4992 14474 4994
rect 9397 4936 9402 4992
rect 9458 4936 14474 4992
rect 9397 4934 14474 4936
rect 14552 5128 18571 5130
rect 14552 5072 18510 5128
rect 18566 5072 18571 5128
rect 14552 5070 18571 5072
rect 9397 4931 9463 4934
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 8293 4858 8359 4861
rect 10225 4858 10291 4861
rect 8293 4856 10291 4858
rect 8293 4800 8298 4856
rect 8354 4800 10230 4856
rect 10286 4800 10291 4856
rect 8293 4798 10291 4800
rect 8293 4795 8359 4798
rect 10225 4795 10291 4798
rect 10593 4858 10659 4861
rect 14552 4858 14612 5070
rect 18505 5067 18571 5070
rect 16573 4994 16639 4997
rect 19006 4994 19012 4996
rect 16573 4992 19012 4994
rect 16573 4936 16578 4992
rect 16634 4936 19012 4992
rect 16573 4934 19012 4936
rect 16573 4931 16639 4934
rect 19006 4932 19012 4934
rect 19076 4994 19082 4996
rect 22520 4994 23000 5024
rect 19076 4934 23000 4994
rect 19076 4932 19082 4934
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 22520 4904 23000 4934
rect 14805 4863 15125 4864
rect 10593 4856 14612 4858
rect 10593 4800 10598 4856
rect 10654 4800 14612 4856
rect 10593 4798 14612 4800
rect 10593 4795 10659 4798
rect 17902 4796 17908 4860
rect 17972 4858 17978 4860
rect 20529 4858 20595 4861
rect 17972 4856 20595 4858
rect 17972 4800 20534 4856
rect 20590 4800 20595 4856
rect 17972 4798 20595 4800
rect 17972 4796 17978 4798
rect 20529 4795 20595 4798
rect 5901 4722 5967 4725
rect 12801 4722 12867 4725
rect 5901 4720 12867 4722
rect 5901 4664 5906 4720
rect 5962 4664 12806 4720
rect 12862 4664 12867 4720
rect 5901 4662 12867 4664
rect 5901 4659 5967 4662
rect 12801 4659 12867 4662
rect 13537 4722 13603 4725
rect 19793 4722 19859 4725
rect 13537 4720 19859 4722
rect 13537 4664 13542 4720
rect 13598 4664 19798 4720
rect 19854 4664 19859 4720
rect 13537 4662 19859 4664
rect 13537 4659 13603 4662
rect 19793 4659 19859 4662
rect 8569 4586 8635 4589
rect 14917 4586 14983 4589
rect 8569 4584 14983 4586
rect 8569 4528 8574 4584
rect 8630 4528 14922 4584
rect 14978 4528 14983 4584
rect 8569 4526 14983 4528
rect 8569 4523 8635 4526
rect 14917 4523 14983 4526
rect 0 4450 480 4480
rect 3969 4450 4035 4453
rect 10225 4452 10291 4453
rect 10174 4450 10180 4452
rect 0 4448 4035 4450
rect 0 4392 3974 4448
rect 4030 4392 4035 4448
rect 0 4390 4035 4392
rect 10134 4390 10180 4450
rect 10244 4448 10291 4452
rect 17953 4450 18019 4453
rect 10286 4392 10291 4448
rect 0 4360 480 4390
rect 3969 4387 4035 4390
rect 10174 4388 10180 4390
rect 10244 4388 10291 4392
rect 10225 4387 10291 4388
rect 11838 4448 18019 4450
rect 11838 4392 17958 4448
rect 18014 4392 18019 4448
rect 11838 4390 18019 4392
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 10317 4178 10383 4181
rect 11838 4178 11898 4390
rect 17953 4387 18019 4390
rect 22369 4450 22435 4453
rect 22520 4450 23000 4480
rect 22369 4448 23000 4450
rect 22369 4392 22374 4448
rect 22430 4392 23000 4448
rect 22369 4390 23000 4392
rect 22369 4387 22435 4390
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22520 4360 23000 4390
rect 18270 4319 18590 4320
rect 13261 4314 13327 4317
rect 14733 4314 14799 4317
rect 13261 4312 14799 4314
rect 13261 4256 13266 4312
rect 13322 4256 14738 4312
rect 14794 4256 14799 4312
rect 13261 4254 14799 4256
rect 13261 4251 13327 4254
rect 14733 4251 14799 4254
rect 14917 4314 14983 4317
rect 17125 4314 17191 4317
rect 14917 4312 17191 4314
rect 14917 4256 14922 4312
rect 14978 4256 17130 4312
rect 17186 4256 17191 4312
rect 14917 4254 17191 4256
rect 14917 4251 14983 4254
rect 17125 4251 17191 4254
rect 10317 4176 11898 4178
rect 10317 4120 10322 4176
rect 10378 4120 11898 4176
rect 10317 4118 11898 4120
rect 12801 4178 12867 4181
rect 16573 4178 16639 4181
rect 12801 4176 16639 4178
rect 12801 4120 12806 4176
rect 12862 4120 16578 4176
rect 16634 4120 16639 4176
rect 12801 4118 16639 4120
rect 10317 4115 10383 4118
rect 12801 4115 12867 4118
rect 16573 4115 16639 4118
rect 0 4042 480 4072
rect 12709 4042 12775 4045
rect 15193 4042 15259 4045
rect 0 4040 15259 4042
rect 0 3984 12714 4040
rect 12770 3984 15198 4040
rect 15254 3984 15259 4040
rect 0 3982 15259 3984
rect 0 3952 480 3982
rect 12709 3979 12775 3982
rect 15193 3979 15259 3982
rect 16113 4042 16179 4045
rect 22520 4042 23000 4072
rect 16113 4040 23000 4042
rect 16113 3984 16118 4040
rect 16174 3984 23000 4040
rect 16113 3982 23000 3984
rect 16113 3979 16179 3982
rect 22520 3952 23000 3982
rect 2589 3906 2655 3909
rect 7281 3906 7347 3909
rect 2589 3904 7347 3906
rect 2589 3848 2594 3904
rect 2650 3848 7286 3904
rect 7342 3848 7347 3904
rect 2589 3846 7347 3848
rect 2589 3843 2655 3846
rect 7281 3843 7347 3846
rect 10225 3906 10291 3909
rect 12198 3906 12204 3908
rect 10225 3904 12204 3906
rect 10225 3848 10230 3904
rect 10286 3848 12204 3904
rect 10225 3846 12204 3848
rect 10225 3843 10291 3846
rect 12198 3844 12204 3846
rect 12268 3844 12274 3908
rect 12617 3906 12683 3909
rect 13077 3906 13143 3909
rect 12617 3904 13143 3906
rect 12617 3848 12622 3904
rect 12678 3848 13082 3904
rect 13138 3848 13143 3904
rect 12617 3846 13143 3848
rect 12617 3843 12683 3846
rect 13077 3843 13143 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 565 3770 631 3773
rect 10133 3770 10199 3773
rect 565 3768 7666 3770
rect 565 3712 570 3768
rect 626 3712 7666 3768
rect 565 3710 7666 3712
rect 565 3707 631 3710
rect 3233 3634 3299 3637
rect 6177 3634 6243 3637
rect 3233 3632 6243 3634
rect 3233 3576 3238 3632
rect 3294 3576 6182 3632
rect 6238 3576 6243 3632
rect 3233 3574 6243 3576
rect 7606 3634 7666 3710
rect 10133 3768 14704 3770
rect 10133 3712 10138 3768
rect 10194 3712 14704 3768
rect 10133 3710 14704 3712
rect 10133 3707 10199 3710
rect 8569 3634 8635 3637
rect 7606 3632 8635 3634
rect 7606 3576 8574 3632
rect 8630 3576 8635 3632
rect 7606 3574 8635 3576
rect 3233 3571 3299 3574
rect 6177 3571 6243 3574
rect 8569 3571 8635 3574
rect 12249 3634 12315 3637
rect 14273 3634 14339 3637
rect 12249 3632 14339 3634
rect 12249 3576 12254 3632
rect 12310 3576 14278 3632
rect 14334 3576 14339 3632
rect 12249 3574 14339 3576
rect 14644 3634 14704 3710
rect 14825 3634 14891 3637
rect 16430 3634 16436 3636
rect 14644 3632 16436 3634
rect 14644 3576 14830 3632
rect 14886 3576 16436 3632
rect 14644 3574 16436 3576
rect 12249 3571 12315 3574
rect 14273 3571 14339 3574
rect 14825 3571 14891 3574
rect 16430 3572 16436 3574
rect 16500 3572 16506 3636
rect 0 3498 480 3528
rect 1669 3498 1735 3501
rect 0 3496 1735 3498
rect 0 3440 1674 3496
rect 1730 3440 1735 3496
rect 0 3438 1735 3440
rect 0 3408 480 3438
rect 1669 3435 1735 3438
rect 1945 3498 2011 3501
rect 14641 3498 14707 3501
rect 1945 3496 14707 3498
rect 1945 3440 1950 3496
rect 2006 3440 14646 3496
rect 14702 3440 14707 3496
rect 1945 3438 14707 3440
rect 1945 3435 2011 3438
rect 14641 3435 14707 3438
rect 18229 3498 18295 3501
rect 22520 3498 23000 3528
rect 18229 3496 23000 3498
rect 18229 3440 18234 3496
rect 18290 3440 23000 3496
rect 18229 3438 23000 3440
rect 18229 3435 18295 3438
rect 22520 3408 23000 3438
rect 5625 3362 5691 3365
rect 10542 3362 10548 3364
rect 5625 3360 10548 3362
rect 5625 3304 5630 3360
rect 5686 3304 10548 3360
rect 5625 3302 10548 3304
rect 5625 3299 5691 3302
rect 10542 3300 10548 3302
rect 10612 3300 10618 3364
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 6729 3226 6795 3229
rect 6729 3224 9874 3226
rect 6729 3168 6734 3224
rect 6790 3168 9874 3224
rect 6729 3166 9874 3168
rect 6729 3163 6795 3166
rect 0 3090 480 3120
rect 1761 3090 1827 3093
rect 0 3088 1827 3090
rect 0 3032 1766 3088
rect 1822 3032 1827 3088
rect 0 3030 1827 3032
rect 0 3000 480 3030
rect 1761 3027 1827 3030
rect 3785 3090 3851 3093
rect 9622 3090 9628 3092
rect 3785 3088 9628 3090
rect 3785 3032 3790 3088
rect 3846 3032 9628 3088
rect 3785 3030 9628 3032
rect 3785 3027 3851 3030
rect 9622 3028 9628 3030
rect 9692 3028 9698 3092
rect 9814 3090 9874 3166
rect 12014 3164 12020 3228
rect 12084 3226 12090 3228
rect 15510 3226 15516 3228
rect 12084 3166 15516 3226
rect 12084 3164 12090 3166
rect 15510 3164 15516 3166
rect 15580 3226 15586 3228
rect 16297 3226 16363 3229
rect 15580 3224 16363 3226
rect 15580 3168 16302 3224
rect 16358 3168 16363 3224
rect 15580 3166 16363 3168
rect 15580 3164 15586 3166
rect 16297 3163 16363 3166
rect 17309 3090 17375 3093
rect 9814 3088 17375 3090
rect 9814 3032 17314 3088
rect 17370 3032 17375 3088
rect 9814 3030 17375 3032
rect 17309 3027 17375 3030
rect 18086 3028 18092 3092
rect 18156 3090 18162 3092
rect 18413 3090 18479 3093
rect 18156 3088 18479 3090
rect 18156 3032 18418 3088
rect 18474 3032 18479 3088
rect 18156 3030 18479 3032
rect 18156 3028 18162 3030
rect 18413 3027 18479 3030
rect 18689 3090 18755 3093
rect 22520 3090 23000 3120
rect 18689 3088 23000 3090
rect 18689 3032 18694 3088
rect 18750 3032 23000 3088
rect 18689 3030 23000 3032
rect 18689 3027 18755 3030
rect 22520 3000 23000 3030
rect 3417 2954 3483 2957
rect 12249 2954 12315 2957
rect 3417 2952 12315 2954
rect 3417 2896 3422 2952
rect 3478 2896 12254 2952
rect 12310 2896 12315 2952
rect 3417 2894 12315 2896
rect 3417 2891 3483 2894
rect 11884 2821 11944 2894
rect 12249 2891 12315 2894
rect 2865 2818 2931 2821
rect 6269 2818 6335 2821
rect 2865 2816 6335 2818
rect 2865 2760 2870 2816
rect 2926 2760 6274 2816
rect 6330 2760 6335 2816
rect 2865 2758 6335 2760
rect 2865 2755 2931 2758
rect 6269 2755 6335 2758
rect 11881 2816 11947 2821
rect 11881 2760 11886 2816
rect 11942 2760 11947 2816
rect 11881 2755 11947 2760
rect 18689 2818 18755 2821
rect 18822 2818 18828 2820
rect 18689 2816 18828 2818
rect 18689 2760 18694 2816
rect 18750 2760 18828 2816
rect 18689 2758 18828 2760
rect 18689 2755 18755 2758
rect 18822 2756 18828 2758
rect 18892 2756 18898 2820
rect 19149 2818 19215 2821
rect 20989 2818 21055 2821
rect 19149 2816 21055 2818
rect 19149 2760 19154 2816
rect 19210 2760 20994 2816
rect 21050 2760 21055 2816
rect 19149 2758 21055 2760
rect 19149 2755 19215 2758
rect 20989 2755 21055 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 10225 2682 10291 2685
rect 10869 2682 10935 2685
rect 10225 2680 10935 2682
rect 10225 2624 10230 2680
rect 10286 2624 10874 2680
rect 10930 2624 10935 2680
rect 10225 2622 10935 2624
rect 10225 2619 10291 2622
rect 10869 2619 10935 2622
rect 13854 2620 13860 2684
rect 13924 2682 13930 2684
rect 13997 2682 14063 2685
rect 13924 2680 14063 2682
rect 13924 2624 14002 2680
rect 14058 2624 14063 2680
rect 13924 2622 14063 2624
rect 13924 2620 13930 2622
rect 13997 2619 14063 2622
rect 18781 2682 18847 2685
rect 19006 2682 19012 2684
rect 18781 2680 19012 2682
rect 18781 2624 18786 2680
rect 18842 2624 19012 2680
rect 18781 2622 19012 2624
rect 18781 2619 18847 2622
rect 19006 2620 19012 2622
rect 19076 2620 19082 2684
rect 0 2546 480 2576
rect 3141 2546 3207 2549
rect 9857 2548 9923 2549
rect 0 2544 3207 2546
rect 0 2488 3146 2544
rect 3202 2488 3207 2544
rect 0 2486 3207 2488
rect 0 2456 480 2486
rect 3141 2483 3207 2486
rect 9806 2484 9812 2548
rect 9876 2546 9923 2548
rect 13997 2546 14063 2549
rect 16573 2546 16639 2549
rect 9876 2544 16639 2546
rect 9918 2488 14002 2544
rect 14058 2488 16578 2544
rect 16634 2488 16639 2544
rect 9876 2486 16639 2488
rect 9876 2484 9923 2486
rect 9857 2483 9923 2484
rect 13997 2483 14063 2486
rect 16573 2483 16639 2486
rect 17125 2546 17191 2549
rect 20478 2546 20484 2548
rect 17125 2544 20484 2546
rect 17125 2488 17130 2544
rect 17186 2488 20484 2544
rect 17125 2486 20484 2488
rect 17125 2483 17191 2486
rect 20478 2484 20484 2486
rect 20548 2484 20554 2548
rect 21081 2546 21147 2549
rect 22520 2546 23000 2576
rect 21081 2544 23000 2546
rect 21081 2488 21086 2544
rect 21142 2488 23000 2544
rect 21081 2486 23000 2488
rect 21081 2483 21147 2486
rect 22520 2456 23000 2486
rect 11145 2410 11211 2413
rect 18321 2410 18387 2413
rect 11145 2408 18387 2410
rect 11145 2352 11150 2408
rect 11206 2352 18326 2408
rect 18382 2352 18387 2408
rect 11145 2350 18387 2352
rect 11145 2347 11211 2350
rect 18321 2347 18387 2350
rect 4409 2208 4729 2209
rect 0 2138 480 2168
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 2048 480 2078
rect 2773 2075 2839 2078
rect 20989 2138 21055 2141
rect 22520 2138 23000 2168
rect 20989 2136 23000 2138
rect 20989 2080 20994 2136
rect 21050 2080 23000 2136
rect 20989 2078 23000 2080
rect 20989 2075 21055 2078
rect 22520 2048 23000 2078
rect 0 1594 480 1624
rect 3233 1594 3299 1597
rect 0 1592 3299 1594
rect 0 1536 3238 1592
rect 3294 1536 3299 1592
rect 0 1534 3299 1536
rect 0 1504 480 1534
rect 3233 1531 3299 1534
rect 20621 1594 20687 1597
rect 22520 1594 23000 1624
rect 20621 1592 23000 1594
rect 20621 1536 20626 1592
rect 20682 1536 23000 1592
rect 20621 1534 23000 1536
rect 20621 1531 20687 1534
rect 22520 1504 23000 1534
rect 0 1186 480 1216
rect 4061 1186 4127 1189
rect 0 1184 4127 1186
rect 0 1128 4066 1184
rect 4122 1128 4127 1184
rect 0 1126 4127 1128
rect 0 1096 480 1126
rect 4061 1123 4127 1126
rect 21725 1186 21791 1189
rect 22520 1186 23000 1216
rect 21725 1184 23000 1186
rect 21725 1128 21730 1184
rect 21786 1128 23000 1184
rect 21725 1126 23000 1128
rect 21725 1123 21791 1126
rect 22520 1096 23000 1126
rect 0 642 480 672
rect 3141 642 3207 645
rect 0 640 3207 642
rect 0 584 3146 640
rect 3202 584 3207 640
rect 0 582 3207 584
rect 0 552 480 582
rect 3141 579 3207 582
rect 20345 642 20411 645
rect 22520 642 23000 672
rect 20345 640 23000 642
rect 20345 584 20350 640
rect 20406 584 23000 640
rect 20345 582 23000 584
rect 20345 579 20411 582
rect 22520 552 23000 582
rect 0 234 480 264
rect 3877 234 3943 237
rect 0 232 3943 234
rect 0 176 3882 232
rect 3938 176 3943 232
rect 0 174 3943 176
rect 0 144 480 174
rect 3877 171 3943 174
rect 21449 234 21515 237
rect 22520 234 23000 264
rect 21449 232 23000 234
rect 21449 176 21454 232
rect 21510 176 23000 232
rect 21449 174 23000 176
rect 21449 171 21515 174
rect 22520 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 13860 19620 13924 19684
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 20300 19408 20364 19412
rect 20300 19352 20314 19408
rect 20314 19352 20364 19408
rect 20300 19348 20364 19352
rect 8340 19076 8404 19140
rect 11836 19136 11900 19140
rect 11836 19080 11850 19136
rect 11850 19080 11900 19136
rect 11836 19076 11900 19080
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 10916 18940 10980 19004
rect 12388 18940 12452 19004
rect 10732 18668 10796 18732
rect 10364 18532 10428 18596
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 8340 18396 8404 18460
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 7604 17716 7668 17780
rect 8524 17580 8588 17644
rect 13676 17444 13740 17508
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 8892 17308 8956 17372
rect 12572 17172 12636 17236
rect 14044 17172 14108 17236
rect 9812 17036 9876 17100
rect 10732 17036 10796 17100
rect 12572 16900 12636 16964
rect 18092 17036 18156 17100
rect 19012 17036 19076 17100
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 9260 16824 9324 16828
rect 9260 16768 9274 16824
rect 9274 16768 9324 16824
rect 9260 16764 9324 16768
rect 10180 16764 10244 16828
rect 7420 16492 7484 16556
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 10364 16084 10428 16148
rect 10548 15948 10612 16012
rect 10916 15948 10980 16012
rect 11836 15948 11900 16012
rect 19380 15948 19444 16012
rect 16988 15812 17052 15876
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 14228 15540 14292 15604
rect 14412 15328 14476 15332
rect 14412 15272 14462 15328
rect 14462 15272 14476 15328
rect 14412 15268 14476 15272
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 9076 14996 9140 15060
rect 14044 14996 14108 15060
rect 7236 14784 7300 14788
rect 7236 14728 7250 14784
rect 7250 14728 7300 14784
rect 7236 14724 7300 14728
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 17172 14588 17236 14652
rect 12204 14452 12268 14516
rect 8892 14316 8956 14380
rect 13860 14180 13924 14244
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 12020 13364 12084 13428
rect 19748 13424 19812 13428
rect 19748 13368 19762 13424
rect 19762 13368 19812 13424
rect 19748 13364 19812 13368
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 14044 12684 14108 12748
rect 12388 12548 12452 12612
rect 16252 12608 16316 12612
rect 16252 12552 16266 12608
rect 16266 12552 16316 12608
rect 16252 12548 16316 12552
rect 20300 12820 20364 12884
rect 17908 12548 17972 12612
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 10916 12412 10980 12476
rect 16804 12412 16868 12476
rect 17540 12472 17604 12476
rect 17540 12416 17554 12472
rect 17554 12416 17604 12472
rect 17540 12412 17604 12416
rect 7236 12276 7300 12340
rect 19196 12276 19260 12340
rect 14228 12140 14292 12204
rect 16804 12200 16868 12204
rect 16804 12144 16854 12200
rect 16854 12144 16868 12200
rect 16804 12140 16868 12144
rect 17540 12140 17604 12204
rect 10180 12004 10244 12068
rect 10364 12064 10428 12068
rect 10364 12008 10414 12064
rect 10414 12008 10428 12064
rect 10364 12004 10428 12008
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 14412 11732 14476 11796
rect 20300 11732 20364 11796
rect 12572 11460 12636 11524
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 9812 11324 9876 11388
rect 16252 11324 16316 11388
rect 9444 11188 9508 11252
rect 10364 11188 10428 11252
rect 18092 11188 18156 11252
rect 9628 11052 9692 11116
rect 12204 11052 12268 11116
rect 20484 11112 20548 11116
rect 20484 11056 20498 11112
rect 20498 11056 20548 11112
rect 20484 11052 20548 11056
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 9260 10840 9324 10844
rect 9260 10784 9274 10840
rect 9274 10784 9324 10840
rect 9260 10780 9324 10784
rect 10732 10644 10796 10708
rect 9444 10432 9508 10436
rect 9444 10376 9458 10432
rect 9458 10376 9508 10432
rect 9444 10372 9508 10376
rect 16988 10372 17052 10436
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 19196 10236 19260 10300
rect 10548 10100 10612 10164
rect 13676 9964 13740 10028
rect 8340 9888 8404 9892
rect 19748 9964 19812 10028
rect 8340 9832 8390 9888
rect 8390 9832 8404 9888
rect 8340 9828 8404 9832
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 7420 9752 7484 9756
rect 7420 9696 7470 9752
rect 7470 9696 7484 9752
rect 7420 9692 7484 9696
rect 8524 9420 8588 9484
rect 8708 9420 8772 9484
rect 8524 9284 8588 9348
rect 11836 9344 11900 9348
rect 11836 9288 11886 9344
rect 11886 9288 11900 9344
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 8340 9208 8404 9212
rect 8340 9152 8390 9208
rect 8390 9152 8404 9208
rect 8340 9148 8404 9152
rect 11836 9284 11900 9288
rect 16436 9480 16500 9484
rect 17172 9556 17236 9620
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 18828 9692 18892 9756
rect 19380 9556 19444 9620
rect 20116 9616 20180 9620
rect 20116 9560 20130 9616
rect 20130 9560 20180 9616
rect 20116 9556 20180 9560
rect 16436 9424 16486 9480
rect 16486 9424 16500 9480
rect 16436 9420 16500 9424
rect 19012 9420 19076 9484
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 15516 9148 15580 9212
rect 10364 9012 10428 9076
rect 9812 8740 9876 8804
rect 16436 8876 16500 8940
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 8708 8468 8772 8532
rect 8524 8332 8588 8396
rect 17908 8332 17972 8396
rect 19196 8332 19260 8396
rect 20116 8332 20180 8396
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 13860 8060 13924 8124
rect 9076 7712 9140 7716
rect 9076 7656 9090 7712
rect 9090 7656 9140 7712
rect 9076 7652 9140 7656
rect 10364 7652 10428 7716
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 12020 6292 12084 6356
rect 13860 6156 13924 6220
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 19380 5808 19444 5812
rect 19380 5752 19394 5808
rect 19394 5752 19444 5808
rect 7604 5612 7668 5676
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 19380 5748 19444 5752
rect 12204 5476 12268 5540
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 12020 5068 12084 5132
rect 17908 5204 17972 5268
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 19012 4932 19076 4996
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 17908 4796 17972 4860
rect 10180 4448 10244 4452
rect 10180 4392 10230 4448
rect 10230 4392 10244 4448
rect 10180 4388 10244 4392
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 12204 3844 12268 3908
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 16436 3572 16500 3636
rect 10548 3300 10612 3364
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 9628 3028 9692 3092
rect 12020 3164 12084 3228
rect 15516 3164 15580 3228
rect 18092 3028 18156 3092
rect 18828 2756 18892 2820
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 13860 2620 13924 2684
rect 19012 2620 19076 2684
rect 9812 2544 9876 2548
rect 9812 2488 9862 2544
rect 9862 2488 9876 2544
rect 9812 2484 9876 2488
rect 20484 2484 20548 2548
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 13859 19684 13925 19685
rect 13859 19620 13860 19684
rect 13924 19620 13925 19684
rect 13859 19619 13925 19620
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 8339 19140 8405 19141
rect 8339 19076 8340 19140
rect 8404 19076 8405 19140
rect 8339 19075 8405 19076
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 8342 18461 8402 19075
rect 10915 19004 10981 19005
rect 10915 18940 10916 19004
rect 10980 18940 10981 19004
rect 10915 18939 10981 18940
rect 10731 18732 10797 18733
rect 10731 18668 10732 18732
rect 10796 18668 10797 18732
rect 10731 18667 10797 18668
rect 10363 18596 10429 18597
rect 10363 18532 10364 18596
rect 10428 18532 10429 18596
rect 10363 18531 10429 18532
rect 8339 18460 8405 18461
rect 8339 18396 8340 18460
rect 8404 18396 8405 18460
rect 8339 18395 8405 18396
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7603 17780 7669 17781
rect 7603 17716 7604 17780
rect 7668 17716 7669 17780
rect 7603 17715 7669 17716
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 7419 16556 7485 16557
rect 7419 16492 7420 16556
rect 7484 16492 7485 16556
rect 7419 16491 7485 16492
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 7235 14788 7301 14789
rect 7235 14724 7236 14788
rect 7300 14724 7301 14788
rect 7235 14723 7301 14724
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 7238 12341 7298 14723
rect 7235 12340 7301 12341
rect 7235 12276 7236 12340
rect 7300 12276 7301 12340
rect 7235 12275 7301 12276
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 7422 9757 7482 16491
rect 7419 9756 7485 9757
rect 7419 9692 7420 9756
rect 7484 9692 7485 9756
rect 7419 9691 7485 9692
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 7606 5677 7666 17715
rect 7874 16896 8195 17920
rect 8523 17644 8589 17645
rect 8523 17580 8524 17644
rect 8588 17580 8589 17644
rect 8523 17579 8589 17580
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 8339 9892 8405 9893
rect 8339 9828 8340 9892
rect 8404 9828 8405 9892
rect 8339 9827 8405 9828
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 8342 9213 8402 9827
rect 8526 9485 8586 17579
rect 8891 17372 8957 17373
rect 8891 17308 8892 17372
rect 8956 17308 8957 17372
rect 8891 17307 8957 17308
rect 8894 14381 8954 17307
rect 9811 17100 9877 17101
rect 9811 17036 9812 17100
rect 9876 17036 9877 17100
rect 9811 17035 9877 17036
rect 9259 16828 9325 16829
rect 9259 16764 9260 16828
rect 9324 16764 9325 16828
rect 9259 16763 9325 16764
rect 9075 15060 9141 15061
rect 9075 14996 9076 15060
rect 9140 14996 9141 15060
rect 9075 14995 9141 14996
rect 8891 14380 8957 14381
rect 8891 14316 8892 14380
rect 8956 14316 8957 14380
rect 8891 14315 8957 14316
rect 8523 9484 8589 9485
rect 8523 9420 8524 9484
rect 8588 9420 8589 9484
rect 8523 9419 8589 9420
rect 8707 9484 8773 9485
rect 8707 9420 8708 9484
rect 8772 9420 8773 9484
rect 8707 9419 8773 9420
rect 8523 9348 8589 9349
rect 8523 9284 8524 9348
rect 8588 9284 8589 9348
rect 8523 9283 8589 9284
rect 8339 9212 8405 9213
rect 8339 9148 8340 9212
rect 8404 9148 8405 9212
rect 8339 9147 8405 9148
rect 8526 8397 8586 9283
rect 8710 8533 8770 9419
rect 8707 8532 8773 8533
rect 8707 8468 8708 8532
rect 8772 8468 8773 8532
rect 8707 8467 8773 8468
rect 8523 8396 8589 8397
rect 8523 8332 8524 8396
rect 8588 8332 8589 8396
rect 8523 8331 8589 8332
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 9078 7717 9138 14995
rect 9262 10845 9322 16763
rect 9814 11389 9874 17035
rect 10179 16828 10245 16829
rect 10179 16764 10180 16828
rect 10244 16764 10245 16828
rect 10179 16763 10245 16764
rect 10182 12069 10242 16763
rect 10366 16149 10426 18531
rect 10734 17101 10794 18667
rect 10731 17100 10797 17101
rect 10731 17036 10732 17100
rect 10796 17036 10797 17100
rect 10731 17035 10797 17036
rect 10363 16148 10429 16149
rect 10363 16084 10364 16148
rect 10428 16084 10429 16148
rect 10363 16083 10429 16084
rect 10366 12069 10426 16083
rect 10547 16012 10613 16013
rect 10547 15948 10548 16012
rect 10612 15948 10613 16012
rect 10547 15947 10613 15948
rect 10179 12068 10245 12069
rect 10179 12004 10180 12068
rect 10244 12004 10245 12068
rect 10179 12003 10245 12004
rect 10363 12068 10429 12069
rect 10363 12004 10364 12068
rect 10428 12004 10429 12068
rect 10363 12003 10429 12004
rect 9811 11388 9877 11389
rect 9811 11324 9812 11388
rect 9876 11324 9877 11388
rect 9811 11323 9877 11324
rect 9443 11252 9509 11253
rect 9443 11188 9444 11252
rect 9508 11188 9509 11252
rect 9443 11187 9509 11188
rect 9259 10844 9325 10845
rect 9259 10780 9260 10844
rect 9324 10780 9325 10844
rect 9259 10779 9325 10780
rect 9446 10437 9506 11187
rect 9627 11116 9693 11117
rect 9627 11052 9628 11116
rect 9692 11052 9693 11116
rect 9627 11051 9693 11052
rect 9443 10436 9509 10437
rect 9443 10372 9444 10436
rect 9508 10372 9509 10436
rect 9443 10371 9509 10372
rect 9075 7716 9141 7717
rect 9075 7652 9076 7716
rect 9140 7652 9141 7716
rect 9075 7651 9141 7652
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7603 5676 7669 5677
rect 7603 5612 7604 5676
rect 7668 5612 7669 5676
rect 7603 5611 7669 5612
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 9630 3093 9690 11051
rect 9811 8804 9877 8805
rect 9811 8740 9812 8804
rect 9876 8740 9877 8804
rect 9811 8739 9877 8740
rect 9627 3092 9693 3093
rect 9627 3028 9628 3092
rect 9692 3028 9693 3092
rect 9627 3027 9693 3028
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 9814 2549 9874 8739
rect 10182 4453 10242 12003
rect 10363 11252 10429 11253
rect 10363 11188 10364 11252
rect 10428 11188 10429 11252
rect 10363 11187 10429 11188
rect 10366 10026 10426 11187
rect 10550 10165 10610 15947
rect 10734 10709 10794 17035
rect 10918 16013 10978 18939
rect 11340 18528 11660 19552
rect 11835 19140 11901 19141
rect 11835 19076 11836 19140
rect 11900 19076 11901 19140
rect 11835 19075 11901 19076
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 10915 16012 10981 16013
rect 10915 15948 10916 16012
rect 10980 15948 10981 16012
rect 10915 15947 10981 15948
rect 10918 12477 10978 15947
rect 11340 15264 11660 16288
rect 11838 16013 11898 19075
rect 12387 19004 12453 19005
rect 12387 18940 12388 19004
rect 12452 18940 12453 19004
rect 12387 18939 12453 18940
rect 11835 16012 11901 16013
rect 11835 15948 11836 16012
rect 11900 15948 11901 16012
rect 11835 15947 11901 15948
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 10915 12476 10981 12477
rect 10915 12412 10916 12476
rect 10980 12412 10981 12476
rect 10915 12411 10981 12412
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 10731 10708 10797 10709
rect 10731 10644 10732 10708
rect 10796 10644 10797 10708
rect 10731 10643 10797 10644
rect 10547 10164 10613 10165
rect 10547 10100 10548 10164
rect 10612 10100 10613 10164
rect 10547 10099 10613 10100
rect 10366 9966 10610 10026
rect 10363 9076 10429 9077
rect 10363 9012 10364 9076
rect 10428 9012 10429 9076
rect 10363 9011 10429 9012
rect 10366 7717 10426 9011
rect 10363 7716 10429 7717
rect 10363 7652 10364 7716
rect 10428 7652 10429 7716
rect 10363 7651 10429 7652
rect 10179 4452 10245 4453
rect 10179 4388 10180 4452
rect 10244 4388 10245 4452
rect 10179 4387 10245 4388
rect 10550 3365 10610 9966
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11838 9349 11898 15947
rect 12203 14516 12269 14517
rect 12203 14452 12204 14516
rect 12268 14452 12269 14516
rect 12203 14451 12269 14452
rect 12019 13428 12085 13429
rect 12019 13364 12020 13428
rect 12084 13364 12085 13428
rect 12019 13363 12085 13364
rect 11835 9348 11901 9349
rect 11835 9284 11836 9348
rect 11900 9284 11901 9348
rect 11835 9283 11901 9284
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 12022 6357 12082 13363
rect 12206 11117 12266 14451
rect 12390 12613 12450 18939
rect 13675 17508 13741 17509
rect 13675 17444 13676 17508
rect 13740 17444 13741 17508
rect 13675 17443 13741 17444
rect 12571 17236 12637 17237
rect 12571 17172 12572 17236
rect 12636 17172 12637 17236
rect 12571 17171 12637 17172
rect 12574 16965 12634 17171
rect 12571 16964 12637 16965
rect 12571 16900 12572 16964
rect 12636 16900 12637 16964
rect 12571 16899 12637 16900
rect 12387 12612 12453 12613
rect 12387 12548 12388 12612
rect 12452 12548 12453 12612
rect 12387 12547 12453 12548
rect 12574 11525 12634 16899
rect 12571 11524 12637 11525
rect 12571 11460 12572 11524
rect 12636 11460 12637 11524
rect 12571 11459 12637 11460
rect 12203 11116 12269 11117
rect 12203 11052 12204 11116
rect 12268 11052 12269 11116
rect 12203 11051 12269 11052
rect 13678 10029 13738 17443
rect 13862 14245 13922 19619
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14043 17236 14109 17237
rect 14043 17172 14044 17236
rect 14108 17172 14109 17236
rect 14043 17171 14109 17172
rect 14046 15061 14106 17171
rect 14805 16896 15125 17920
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 20299 19412 20365 19413
rect 20299 19348 20300 19412
rect 20364 19348 20365 19412
rect 20299 19347 20365 19348
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18091 17100 18157 17101
rect 18091 17036 18092 17100
rect 18156 17036 18157 17100
rect 18091 17035 18157 17036
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 16987 15876 17053 15877
rect 16987 15812 16988 15876
rect 17052 15812 17053 15876
rect 16987 15811 17053 15812
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14227 15604 14293 15605
rect 14227 15540 14228 15604
rect 14292 15540 14293 15604
rect 14227 15539 14293 15540
rect 14043 15060 14109 15061
rect 14043 14996 14044 15060
rect 14108 14996 14109 15060
rect 14043 14995 14109 14996
rect 13859 14244 13925 14245
rect 13859 14180 13860 14244
rect 13924 14180 13925 14244
rect 13859 14179 13925 14180
rect 14046 12749 14106 14995
rect 14043 12748 14109 12749
rect 14043 12684 14044 12748
rect 14108 12684 14109 12748
rect 14043 12683 14109 12684
rect 14230 12205 14290 15539
rect 14411 15332 14477 15333
rect 14411 15268 14412 15332
rect 14476 15268 14477 15332
rect 14411 15267 14477 15268
rect 14227 12204 14293 12205
rect 14227 12140 14228 12204
rect 14292 12140 14293 12204
rect 14227 12139 14293 12140
rect 14414 11797 14474 15267
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 16251 12612 16317 12613
rect 16251 12548 16252 12612
rect 16316 12548 16317 12612
rect 16251 12547 16317 12548
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14411 11796 14477 11797
rect 14411 11732 14412 11796
rect 14476 11732 14477 11796
rect 14411 11731 14477 11732
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 16254 11389 16314 12547
rect 16803 12476 16869 12477
rect 16803 12412 16804 12476
rect 16868 12412 16869 12476
rect 16803 12411 16869 12412
rect 16806 12205 16866 12411
rect 16803 12204 16869 12205
rect 16803 12140 16804 12204
rect 16868 12140 16869 12204
rect 16803 12139 16869 12140
rect 16251 11388 16317 11389
rect 16251 11324 16252 11388
rect 16316 11324 16317 11388
rect 16251 11323 16317 11324
rect 16990 10437 17050 15811
rect 17171 14652 17237 14653
rect 17171 14588 17172 14652
rect 17236 14588 17237 14652
rect 17171 14587 17237 14588
rect 16987 10436 17053 10437
rect 16987 10372 16988 10436
rect 17052 10372 17053 10436
rect 16987 10371 17053 10372
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 13675 10028 13741 10029
rect 13675 9964 13676 10028
rect 13740 9964 13741 10028
rect 13675 9963 13741 9964
rect 14805 9280 15125 10304
rect 17174 9621 17234 14587
rect 17907 12612 17973 12613
rect 17907 12548 17908 12612
rect 17972 12548 17973 12612
rect 17907 12547 17973 12548
rect 17539 12476 17605 12477
rect 17539 12412 17540 12476
rect 17604 12412 17605 12476
rect 17539 12411 17605 12412
rect 17542 12205 17602 12411
rect 17539 12204 17605 12205
rect 17539 12140 17540 12204
rect 17604 12140 17605 12204
rect 17539 12139 17605 12140
rect 17171 9620 17237 9621
rect 17171 9556 17172 9620
rect 17236 9556 17237 9620
rect 17171 9555 17237 9556
rect 16435 9484 16501 9485
rect 16435 9420 16436 9484
rect 16500 9420 16501 9484
rect 16435 9419 16501 9420
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 15515 9212 15581 9213
rect 15515 9148 15516 9212
rect 15580 9148 15581 9212
rect 15515 9147 15581 9148
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 13859 8124 13925 8125
rect 13859 8060 13860 8124
rect 13924 8060 13925 8124
rect 13859 8059 13925 8060
rect 12019 6356 12085 6357
rect 12019 6292 12020 6356
rect 12084 6292 12085 6356
rect 12019 6291 12085 6292
rect 13862 6221 13922 8059
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 13859 6220 13925 6221
rect 13859 6156 13860 6220
rect 13924 6156 13925 6220
rect 13859 6155 13925 6156
rect 12203 5540 12269 5541
rect 12203 5476 12204 5540
rect 12268 5476 12269 5540
rect 12203 5475 12269 5476
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 12019 5132 12085 5133
rect 12019 5068 12020 5132
rect 12084 5068 12085 5132
rect 12019 5067 12085 5068
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 10547 3364 10613 3365
rect 10547 3300 10548 3364
rect 10612 3300 10613 3364
rect 10547 3299 10613 3300
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9811 2548 9877 2549
rect 9811 2484 9812 2548
rect 9876 2484 9877 2548
rect 9811 2483 9877 2484
rect 11340 2208 11660 3232
rect 12022 3229 12082 5067
rect 12206 3909 12266 5475
rect 12203 3908 12269 3909
rect 12203 3844 12204 3908
rect 12268 3844 12269 3908
rect 12203 3843 12269 3844
rect 12019 3228 12085 3229
rect 12019 3164 12020 3228
rect 12084 3164 12085 3228
rect 12019 3163 12085 3164
rect 13862 2685 13922 6155
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 15518 3229 15578 9147
rect 16438 8941 16498 9419
rect 16435 8940 16501 8941
rect 16435 8876 16436 8940
rect 16500 8876 16501 8940
rect 16435 8875 16501 8876
rect 16438 3637 16498 8875
rect 17910 8397 17970 12547
rect 18094 11253 18154 17035
rect 18270 16352 18590 17376
rect 19011 17100 19077 17101
rect 19011 17036 19012 17100
rect 19076 17036 19077 17100
rect 19011 17035 19077 17036
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 14176 18590 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 12000 18590 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18091 11252 18157 11253
rect 18091 11188 18092 11252
rect 18156 11188 18157 11252
rect 18091 11187 18157 11188
rect 17907 8396 17973 8397
rect 17907 8332 17908 8396
rect 17972 8332 17973 8396
rect 17907 8331 17973 8332
rect 17907 5268 17973 5269
rect 17907 5204 17908 5268
rect 17972 5204 17973 5268
rect 17907 5203 17973 5204
rect 17910 4861 17970 5203
rect 17907 4860 17973 4861
rect 17907 4796 17908 4860
rect 17972 4796 17973 4860
rect 17907 4795 17973 4796
rect 16435 3636 16501 3637
rect 16435 3572 16436 3636
rect 16500 3572 16501 3636
rect 16435 3571 16501 3572
rect 15515 3228 15581 3229
rect 15515 3164 15516 3228
rect 15580 3164 15581 3228
rect 15515 3163 15581 3164
rect 18094 3093 18154 11187
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 9824 18590 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 8736 18590 9760
rect 18827 9756 18893 9757
rect 18827 9692 18828 9756
rect 18892 9692 18893 9756
rect 18827 9691 18893 9692
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 3296 18590 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18091 3092 18157 3093
rect 18091 3028 18092 3092
rect 18156 3028 18157 3092
rect 18091 3027 18157 3028
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 13859 2684 13925 2685
rect 13859 2620 13860 2684
rect 13924 2620 13925 2684
rect 13859 2619 13925 2620
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 2128 15125 2688
rect 18270 2208 18590 3232
rect 18830 2821 18890 9691
rect 19014 9485 19074 17035
rect 19379 16012 19445 16013
rect 19379 15948 19380 16012
rect 19444 15948 19445 16012
rect 19379 15947 19445 15948
rect 19195 12340 19261 12341
rect 19195 12276 19196 12340
rect 19260 12338 19261 12340
rect 19382 12338 19442 15947
rect 19747 13428 19813 13429
rect 19747 13364 19748 13428
rect 19812 13364 19813 13428
rect 19747 13363 19813 13364
rect 19260 12278 19442 12338
rect 19260 12276 19261 12278
rect 19195 12275 19261 12276
rect 19195 10300 19261 10301
rect 19195 10236 19196 10300
rect 19260 10236 19261 10300
rect 19195 10235 19261 10236
rect 19011 9484 19077 9485
rect 19011 9420 19012 9484
rect 19076 9420 19077 9484
rect 19011 9419 19077 9420
rect 19198 8397 19258 10235
rect 19750 10029 19810 13363
rect 20302 12885 20362 19347
rect 20299 12884 20365 12885
rect 20299 12820 20300 12884
rect 20364 12820 20365 12884
rect 20299 12819 20365 12820
rect 20302 11797 20362 12819
rect 20299 11796 20365 11797
rect 20299 11732 20300 11796
rect 20364 11732 20365 11796
rect 20299 11731 20365 11732
rect 20483 11116 20549 11117
rect 20483 11052 20484 11116
rect 20548 11052 20549 11116
rect 20483 11051 20549 11052
rect 19747 10028 19813 10029
rect 19747 9964 19748 10028
rect 19812 9964 19813 10028
rect 19747 9963 19813 9964
rect 19379 9620 19445 9621
rect 19379 9556 19380 9620
rect 19444 9556 19445 9620
rect 19379 9555 19445 9556
rect 20115 9620 20181 9621
rect 20115 9556 20116 9620
rect 20180 9556 20181 9620
rect 20115 9555 20181 9556
rect 19195 8396 19261 8397
rect 19195 8332 19196 8396
rect 19260 8332 19261 8396
rect 19195 8331 19261 8332
rect 19382 5813 19442 9555
rect 20118 8397 20178 9555
rect 20115 8396 20181 8397
rect 20115 8332 20116 8396
rect 20180 8332 20181 8396
rect 20115 8331 20181 8332
rect 19379 5812 19445 5813
rect 19379 5748 19380 5812
rect 19444 5748 19445 5812
rect 19379 5747 19445 5748
rect 19011 4996 19077 4997
rect 19011 4932 19012 4996
rect 19076 4932 19077 4996
rect 19011 4931 19077 4932
rect 18827 2820 18893 2821
rect 18827 2756 18828 2820
rect 18892 2756 18893 2820
rect 18827 2755 18893 2756
rect 19014 2685 19074 4931
rect 19011 2684 19077 2685
rect 19011 2620 19012 2684
rect 19076 2620 19077 2684
rect 19011 2619 19077 2620
rect 20486 2549 20546 11051
rect 20483 2548 20549 2549
rect 20483 2484 20484 2548
rect 20548 2484 20549 2548
rect 20483 2483 20549 2484
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1604681595
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1604681595
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 8648 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1604681595
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_75 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_81
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _110_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10396 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1604681595
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1604681595
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14444 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1604681595
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_163
timestamp 1604681595
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1604681595
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1604681595
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19320 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1604681595
transform 1 0 21252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1604681595
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7912 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9752 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11408 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_110
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_121
timestamp 1604681595
transform 1 0 12236 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_143
timestamp 1604681595
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1604681595
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17572 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16560 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_167
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1604681595
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1604681595
transform 1 0 18124 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_198
timestamp 1604681595
transform 1 0 19320 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1604681595
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1604681595
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_34
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1604681595
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1604681595
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_111
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13708 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 14536 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16928 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_168
timestamp 1604681595
transform 1 0 16560 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18400 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_20
timestamp 1604681595
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4324 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_25
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8188 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_86
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_4_113
timestamp 1604681595
transform 1 0 11500 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14260 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15824 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1604681595
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19412 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_198
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_208
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_18
timestamp 1604681595
transform 1 0 2760 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3128 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_38
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1604681595
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1604681595
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 9660 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1604681595
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1604681595
transform 1 0 11500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 12696 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_130
timestamp 1604681595
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_141
timestamp 1604681595
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1604681595
transform 1 0 18124 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_174
timestamp 1604681595
transform 1 0 17112 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1604681595
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_194
timestamp 1604681595
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_205
timestamp 1604681595
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20332 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1604681595
transform 1 0 21160 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1604681595
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1840 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_24
timestamp 1604681595
transform 1 0 3312 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1604681595
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp 1604681595
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1604681595
transform 1 0 6072 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5520 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_53
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1604681595
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7268 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1604681595
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_76
timestamp 1604681595
transform 1 0 8096 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9936 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9568 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp 1604681595
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1604681595
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp 1604681595
transform 1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1604681595
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_106
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604681595
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12880 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_144
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_150
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1604681595
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 14996 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15364 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_171
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_182
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 18032 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_187
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18492 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1604681595
transform 1 0 20056 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_205
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 21068 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1604681595
transform 1 0 21252 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_215
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1604681595
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_25
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1604681595
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp 1604681595
transform 1 0 5428 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1604681595
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10672 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12328 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1604681595
transform 1 0 13156 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_140
timestamp 1604681595
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 15548 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1604681595
transform 1 0 17112 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_172
timestamp 1604681595
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_183
timestamp 1604681595
transform 1 0 17940 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 20148 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1604681595
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_218
timestamp 1604681595
transform 1 0 21160 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1604681595
transform 1 0 21528 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1604681595
transform 1 0 3312 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1604681595
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_33
timestamp 1604681595
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_56
timestamp 1604681595
transform 1 0 6256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1604681595
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7452 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_68
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10672 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13432 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 15364 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_150
timestamp 1604681595
transform 1 0 14904 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18676 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_207
timestamp 1604681595
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1604681595
transform 1 0 20332 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_218
timestamp 1604681595
transform 1 0 21160 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1604681595
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp 1604681595
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_51
timestamp 1604681595
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_55
timestamp 1604681595
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8280 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1604681595
transform 1 0 9936 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_116
timestamp 1604681595
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1604681595
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12696 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_142
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17940 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1604681595
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_192
timestamp 1604681595
transform 1 0 18768 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_24
timestamp 1604681595
transform 1 0 3312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5244 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp 1604681595
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_145
timestamp 1604681595
transform 1 0 14444 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 14996 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_163
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_192
timestamp 1604681595
transform 1 0 18768 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1604681595
transform 1 0 19688 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1840 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_24
timestamp 1604681595
transform 1 0 3312 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604681595
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6072 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1604681595
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_74
timestamp 1604681595
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1604681595
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12328 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_111
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_119
timestamp 1604681595
transform 1 0 12052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17388 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_174
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_204
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1604681595
transform 1 0 21160 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1604681595
transform 1 0 21528 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1604681595
transform 1 0 2852 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1604681595
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_21
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_40
timestamp 1604681595
transform 1 0 4784 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6532 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 1604681595
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_57
timestamp 1604681595
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_82
timestamp 1604681595
transform 1 0 8648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12236 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10948 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_116
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 14444 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_148
timestamp 1604681595
transform 1 0 14720 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1604681595
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16928 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1604681595
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_181
timestamp 1604681595
transform 1 0 17756 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_200
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 20424 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1604681595
transform 1 0 21252 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1604681595
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1604681595
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_18
timestamp 1604681595
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_29
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_76
timestamp 1604681595
transform 1 0 8096 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1604681595
transform 1 0 10488 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10856 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14444 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_143
timestamp 1604681595
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1604681595
transform 1 0 15272 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1604681595
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_197
timestamp 1604681595
transform 1 0 19228 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 20976 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_214
timestamp 1604681595
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1604681595
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5796 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1604681595
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_76
timestamp 1604681595
transform 1 0 8096 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10304 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12144 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1604681595
transform 1 0 17112 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_195
timestamp 1604681595
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1604681595
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_12
timestamp 1604681595
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 6256 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5244 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1604681595
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9476 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_100
timestamp 1604681595
transform 1 0 10304 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20056 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_204
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_52
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_78
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_117
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13708 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_135
timestamp 1604681595
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_146
timestamp 1604681595
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1604681595
transform 1 0 15732 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_179
timestamp 1604681595
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19504 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1604681595
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4324 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1604681595
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_42
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1604681595
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1604681595
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1604681595
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6348 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8372 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1604681595
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11132 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12144 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_107
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_117
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 13340 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13708 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 13432 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_151
timestamp 1604681595
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_146
timestamp 1604681595
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 14720 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16284 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 16284 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_174
timestamp 1604681595
transform 1 0 17112 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_180
timestamp 1604681595
transform 1 0 17664 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18400 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19780 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19688 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1604681595
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_201
timestamp 1604681595
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20700 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1604681595
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1604681595
transform 1 0 21252 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1604681595
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_18
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3036 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_37
timestamp 1604681595
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7084 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_21_81
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1604681595
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11132 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1604681595
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13340 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 13064 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1604681595
transform 1 0 12696 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15180 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1604681595
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1604681595
transform 1 0 20056 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_204
timestamp 1604681595
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2300 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 3312 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_22
timestamp 1604681595
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_28
timestamp 1604681595
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1604681595
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_83
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11776 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1604681595
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13984 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1604681595
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_22_174
timestamp 1604681595
transform 1 0 17112 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_180
timestamp 1604681595
transform 1 0 17664 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19780 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_201
timestamp 1604681595
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1604681595
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 1656 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1604681595
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_18
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5244 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1604681595
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1604681595
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_83
timestamp 1604681595
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10488 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1604681595
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_96
timestamp 1604681595
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1604681595
transform 1 0 14076 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1604681595
transform 1 0 13708 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15824 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_150
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1604681595
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 17480 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_176
timestamp 1604681595
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19688 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1604681595
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_211
timestamp 1604681595
transform 1 0 20516 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1604681595
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 1472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1604681595
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_8
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1604681595
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5428 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1604681595
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_81
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_108
timestamp 1604681595
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1604681595
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_137
timestamp 1604681595
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1604681595
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_163
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 16560 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1604681595
transform 1 0 16468 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_195
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1604681595
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_20
timestamp 1604681595
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5704 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_43
timestamp 1604681595
transform 1 0 5060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 1604681595
transform 1 0 5612 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6900 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1604681595
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1604681595
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14076 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1604681595
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_150
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1604681595
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1604681595
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1604681595
transform 1 0 19320 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_197
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_207
timestamp 1604681595
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20332 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1604681595
transform 1 0 21160 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1604681595
transform 1 0 21528 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_17
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1604681595
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1604681595
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1604681595
transform 1 0 4324 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_34
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6164 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_52
timestamp 1604681595
transform 1 0 5888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_49
timestamp 1604681595
transform 1 0 5612 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_64
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9844 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_104
timestamp 1604681595
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 11684 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10856 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1604681595
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1604681595
transform 1 0 12696 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_139
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 14720 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_146
timestamp 1604681595
transform 1 0 14536 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_158
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17296 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18308 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_174
timestamp 1604681595
transform 1 0 17112 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_185
timestamp 1604681595
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1604681595
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1604681595
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18400 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19320 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_196
timestamp 1604681595
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_207
timestamp 1604681595
transform 1 0 20148 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604681595
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1604681595
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1604681595
transform 1 0 21252 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2944 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5336 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_45
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_62
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1604681595
transform 1 0 7452 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_78
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_89
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11316 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1604681595
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_120
timestamp 1604681595
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_143
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1604681595
transform 1 0 17112 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_187
timestamp 1604681595
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1604681595
transform 1 0 18492 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1604681595
transform 1 0 19780 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_198
timestamp 1604681595
transform 1 0 19320 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1604681595
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 1604681595
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_46
timestamp 1604681595
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_73
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_83
timestamp 1604681595
transform 1 0 8740 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12512 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11040 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1604681595
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1604681595
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1604681595
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_133
timestamp 1604681595
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_150
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_155
timestamp 1604681595
transform 1 0 15364 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_163
timestamp 1604681595
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_174
timestamp 1604681595
transform 1 0 17112 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604681595
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18400 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_197
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_207
timestamp 1604681595
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 21068 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20332 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1604681595
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 1656 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1604681595
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5704 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5060 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1604681595
transform 1 0 6716 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_49
timestamp 1604681595
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1604681595
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 7912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8372 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6900 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_72
timestamp 1604681595
transform 1 0 7728 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1604681595
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1604681595
transform 1 0 11684 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12236 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 1604681595
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_119
timestamp 1604681595
transform 1 0 12052 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_137
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1604681595
transform 1 0 14720 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1604681595
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17204 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_174
timestamp 1604681595
transform 1 0 17112 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_181
timestamp 1604681595
transform 1 0 17756 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_191
timestamp 1604681595
transform 1 0 18676 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_199
timestamp 1604681595
transform 1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1604681595
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5704 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_78
timestamp 1604681595
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9568 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_89
timestamp 1604681595
transform 1 0 9292 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_108
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14076 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1604681595
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15916 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15088 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_150
timestamp 1604681595
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_158
timestamp 1604681595
transform 1 0 15640 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1604681595
transform 1 0 16652 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_167
timestamp 1604681595
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_173
timestamp 1604681595
transform 1 0 17020 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 19688 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_188
timestamp 1604681595
transform 1 0 18400 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1604681595
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1604681595
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1604681595
transform 1 0 21160 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1604681595
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604681595
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_17
timestamp 1604681595
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4324 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5980 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_51
timestamp 1604681595
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7636 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_69
timestamp 1604681595
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_87
timestamp 1604681595
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1604681595
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11960 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_116
timestamp 1604681595
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1604681595
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1604681595
transform 1 0 16284 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15548 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1604681595
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 16836 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1604681595
transform 1 0 17572 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_169
timestamp 1604681595
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp 1604681595
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_183
timestamp 1604681595
transform 1 0 17940 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 19136 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1604681595
transform 1 0 18492 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_200
timestamp 1604681595
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1604681595
transform 1 0 21252 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1604681595
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_17
timestamp 1604681595
transform 1 0 2668 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_29
timestamp 1604681595
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_48
timestamp 1604681595
transform 1 0 5520 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7360 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_63
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_67
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1604681595
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_88
timestamp 1604681595
transform 1 0 9200 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_92
timestamp 1604681595
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 11316 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_109
timestamp 1604681595
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_134
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_142
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1604681595
transform 1 0 14812 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_148
timestamp 1604681595
transform 1 0 14720 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_153
timestamp 1604681595
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1604681595
transform 1 0 16100 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1604681595
transform 1 0 16468 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_183
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_187
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 19320 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_195
timestamp 1604681595
transform 1 0 19044 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_202
timestamp 1604681595
transform 1 0 19688 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 20516 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1030 0 1086 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2410 0 2466 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 4250 0 4306 480 6 ccff_head
port 8 nsew default input
rlabel metal2 s 4710 0 4766 480 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 22520 3952 23000 4072 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 22520 8712 23000 8832 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 22520 9120 23000 9240 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 22520 9664 23000 9784 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 22520 10072 23000 10192 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 22520 10616 23000 10736 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 22520 11024 23000 11144 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 22520 11568 23000 11688 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 22520 12112 23000 12232 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 22520 12520 23000 12640 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 22520 13064 23000 13184 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 22520 4360 23000 4480 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 22520 4904 23000 5024 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 22520 5312 23000 5432 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 22520 5856 23000 5976 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 22520 6264 23000 6384 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 22520 6808 23000 6928 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 22520 7216 23000 7336 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 22520 7760 23000 7880 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 22520 8168 23000 8288 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 22520 13472 23000 13592 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 22520 18232 23000 18352 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 22520 18776 23000 18896 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 22520 19184 23000 19304 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 22520 19728 23000 19848 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 22520 20136 23000 20256 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 22520 20680 23000 20800 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 22520 21088 23000 21208 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 22520 21632 23000 21752 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 22520 22040 23000 22160 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 22520 22584 23000 22704 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 22520 14016 23000 14136 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 22520 14424 23000 14544 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 22520 14968 23000 15088 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 22520 15376 23000 15496 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 22520 15920 23000 16040 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 22520 16328 23000 16448 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 22520 16872 23000 16992 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 22520 17280 23000 17400 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 22520 17824 23000 17944 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 12346 0 12402 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 19982 0 20038 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 22282 0 22338 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal2 s 3974 22520 4030 23000 6 chany_top_in[0]
port 130 nsew default input
rlabel metal2 s 8758 22520 8814 23000 6 chany_top_in[10]
port 131 nsew default input
rlabel metal2 s 9218 22520 9274 23000 6 chany_top_in[11]
port 132 nsew default input
rlabel metal2 s 9770 22520 9826 23000 6 chany_top_in[12]
port 133 nsew default input
rlabel metal2 s 10230 22520 10286 23000 6 chany_top_in[13]
port 134 nsew default input
rlabel metal2 s 10690 22520 10746 23000 6 chany_top_in[14]
port 135 nsew default input
rlabel metal2 s 11150 22520 11206 23000 6 chany_top_in[15]
port 136 nsew default input
rlabel metal2 s 11702 22520 11758 23000 6 chany_top_in[16]
port 137 nsew default input
rlabel metal2 s 12162 22520 12218 23000 6 chany_top_in[17]
port 138 nsew default input
rlabel metal2 s 12622 22520 12678 23000 6 chany_top_in[18]
port 139 nsew default input
rlabel metal2 s 13082 22520 13138 23000 6 chany_top_in[19]
port 140 nsew default input
rlabel metal2 s 4434 22520 4490 23000 6 chany_top_in[1]
port 141 nsew default input
rlabel metal2 s 4986 22520 5042 23000 6 chany_top_in[2]
port 142 nsew default input
rlabel metal2 s 5446 22520 5502 23000 6 chany_top_in[3]
port 143 nsew default input
rlabel metal2 s 5906 22520 5962 23000 6 chany_top_in[4]
port 144 nsew default input
rlabel metal2 s 6366 22520 6422 23000 6 chany_top_in[5]
port 145 nsew default input
rlabel metal2 s 6826 22520 6882 23000 6 chany_top_in[6]
port 146 nsew default input
rlabel metal2 s 7378 22520 7434 23000 6 chany_top_in[7]
port 147 nsew default input
rlabel metal2 s 7838 22520 7894 23000 6 chany_top_in[8]
port 148 nsew default input
rlabel metal2 s 8298 22520 8354 23000 6 chany_top_in[9]
port 149 nsew default input
rlabel metal2 s 13542 22520 13598 23000 6 chany_top_out[0]
port 150 nsew default tristate
rlabel metal2 s 18326 22520 18382 23000 6 chany_top_out[10]
port 151 nsew default tristate
rlabel metal2 s 18878 22520 18934 23000 6 chany_top_out[11]
port 152 nsew default tristate
rlabel metal2 s 19338 22520 19394 23000 6 chany_top_out[12]
port 153 nsew default tristate
rlabel metal2 s 19798 22520 19854 23000 6 chany_top_out[13]
port 154 nsew default tristate
rlabel metal2 s 20258 22520 20314 23000 6 chany_top_out[14]
port 155 nsew default tristate
rlabel metal2 s 20718 22520 20774 23000 6 chany_top_out[15]
port 156 nsew default tristate
rlabel metal2 s 21270 22520 21326 23000 6 chany_top_out[16]
port 157 nsew default tristate
rlabel metal2 s 21730 22520 21786 23000 6 chany_top_out[17]
port 158 nsew default tristate
rlabel metal2 s 22190 22520 22246 23000 6 chany_top_out[18]
port 159 nsew default tristate
rlabel metal2 s 22650 22520 22706 23000 6 chany_top_out[19]
port 160 nsew default tristate
rlabel metal2 s 14094 22520 14150 23000 6 chany_top_out[1]
port 161 nsew default tristate
rlabel metal2 s 14554 22520 14610 23000 6 chany_top_out[2]
port 162 nsew default tristate
rlabel metal2 s 15014 22520 15070 23000 6 chany_top_out[3]
port 163 nsew default tristate
rlabel metal2 s 15474 22520 15530 23000 6 chany_top_out[4]
port 164 nsew default tristate
rlabel metal2 s 15934 22520 15990 23000 6 chany_top_out[5]
port 165 nsew default tristate
rlabel metal2 s 16486 22520 16542 23000 6 chany_top_out[6]
port 166 nsew default tristate
rlabel metal2 s 16946 22520 17002 23000 6 chany_top_out[7]
port 167 nsew default tristate
rlabel metal2 s 17406 22520 17462 23000 6 chany_top_out[8]
port 168 nsew default tristate
rlabel metal2 s 17866 22520 17922 23000 6 chany_top_out[9]
port 169 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 170 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 171 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_36_
port 172 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 173 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_38_
port 174 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 175 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_40_
port 176 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 177 nsew default input
rlabel metal2 s 3790 0 3846 480 6 prog_clk
port 178 nsew default input
rlabel metal3 s 22520 144 23000 264 6 right_bottom_grid_pin_34_
port 179 nsew default input
rlabel metal3 s 22520 552 23000 672 6 right_bottom_grid_pin_35_
port 180 nsew default input
rlabel metal3 s 22520 1096 23000 1216 6 right_bottom_grid_pin_36_
port 181 nsew default input
rlabel metal3 s 22520 1504 23000 1624 6 right_bottom_grid_pin_37_
port 182 nsew default input
rlabel metal3 s 22520 2048 23000 2168 6 right_bottom_grid_pin_38_
port 183 nsew default input
rlabel metal3 s 22520 2456 23000 2576 6 right_bottom_grid_pin_39_
port 184 nsew default input
rlabel metal3 s 22520 3000 23000 3120 6 right_bottom_grid_pin_40_
port 185 nsew default input
rlabel metal3 s 22520 3408 23000 3528 6 right_bottom_grid_pin_41_
port 186 nsew default input
rlabel metal2 s 202 22520 258 23000 6 top_left_grid_pin_42_
port 187 nsew default input
rlabel metal2 s 662 22520 718 23000 6 top_left_grid_pin_43_
port 188 nsew default input
rlabel metal2 s 1122 22520 1178 23000 6 top_left_grid_pin_44_
port 189 nsew default input
rlabel metal2 s 1582 22520 1638 23000 6 top_left_grid_pin_45_
port 190 nsew default input
rlabel metal2 s 2042 22520 2098 23000 6 top_left_grid_pin_46_
port 191 nsew default input
rlabel metal2 s 2594 22520 2650 23000 6 top_left_grid_pin_47_
port 192 nsew default input
rlabel metal2 s 3054 22520 3110 23000 6 top_left_grid_pin_48_
port 193 nsew default input
rlabel metal2 s 3514 22520 3570 23000 6 top_left_grid_pin_49_
port 194 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 195 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 196 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
