magic
tech sky130A
magscale 1 2
timestamp 1606226928
<< locali >>
rect 17785 19227 17819 19465
rect 5825 18683 5859 18921
rect 9505 18819 9539 18921
rect 19073 18683 19107 18785
rect 12173 18071 12207 18241
rect 13461 18139 13495 18309
rect 16405 15351 16439 15453
rect 6101 14875 6135 14977
rect 7665 14807 7699 14909
rect 8677 14807 8711 15113
rect 15669 14807 15703 14977
rect 15761 14943 15795 15113
rect 12265 12631 12299 12937
rect 13829 12631 13863 12937
rect 17785 12767 17819 12869
rect 6009 12223 6043 12325
rect 4261 11611 4295 11781
rect 3893 10999 3927 11169
rect 11805 10115 11839 10217
rect 7665 9911 7699 10081
rect 10241 9367 10275 9537
rect 13369 9435 13403 9605
rect 16865 9503 16899 9673
rect 4905 8483 4939 8585
rect 14565 8347 14599 8517
<< viali >>
rect 1961 20009 1995 20043
rect 12173 20009 12207 20043
rect 14105 20009 14139 20043
rect 15025 20009 15059 20043
rect 15853 20009 15887 20043
rect 16405 20009 16439 20043
rect 17141 20009 17175 20043
rect 17877 20009 17911 20043
rect 20177 20009 20211 20043
rect 20729 20009 20763 20043
rect 1777 19873 1811 19907
rect 2335 19873 2369 19907
rect 2881 19873 2915 19907
rect 3433 19873 3467 19907
rect 11989 19873 12023 19907
rect 13093 19873 13127 19907
rect 13185 19873 13219 19907
rect 13921 19873 13955 19907
rect 14841 19873 14875 19907
rect 15669 19873 15703 19907
rect 16221 19873 16255 19907
rect 16957 19873 16991 19907
rect 17693 19873 17727 19907
rect 18337 19873 18371 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 13369 19805 13403 19839
rect 18521 19805 18555 19839
rect 19625 19737 19659 19771
rect 2513 19669 2547 19703
rect 3065 19669 3099 19703
rect 3617 19669 3651 19703
rect 12725 19669 12759 19703
rect 1961 19465 1995 19499
rect 3709 19465 3743 19499
rect 4261 19465 4295 19499
rect 16957 19465 16991 19499
rect 17785 19465 17819 19499
rect 18061 19465 18095 19499
rect 11713 19329 11747 19363
rect 15761 19329 15795 19363
rect 17601 19329 17635 19363
rect 1777 19261 1811 19295
rect 2605 19261 2639 19295
rect 3525 19261 3559 19295
rect 4077 19261 4111 19295
rect 4629 19261 4663 19295
rect 10517 19261 10551 19295
rect 11437 19261 11471 19295
rect 12449 19261 12483 19295
rect 13185 19261 13219 19295
rect 16129 19261 16163 19295
rect 16405 19261 16439 19295
rect 18613 19329 18647 19363
rect 19073 19261 19107 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 10793 19193 10827 19227
rect 12725 19193 12759 19227
rect 13452 19193 13486 19227
rect 17417 19193 17451 19227
rect 17785 19193 17819 19227
rect 18521 19193 18555 19227
rect 19349 19193 19383 19227
rect 2789 19125 2823 19159
rect 4813 19125 4847 19159
rect 14565 19125 14599 19159
rect 15117 19125 15151 19159
rect 15485 19125 15519 19159
rect 15577 19125 15611 19159
rect 17325 19125 17359 19159
rect 18429 19125 18463 19159
rect 20177 19125 20211 19159
rect 20729 19125 20763 19159
rect 1961 18921 1995 18955
rect 2513 18921 2547 18955
rect 5825 18921 5859 18955
rect 8309 18921 8343 18955
rect 9505 18921 9539 18955
rect 13461 18921 13495 18955
rect 15485 18921 15519 18955
rect 20453 18921 20487 18955
rect 3249 18853 3283 18887
rect 1777 18785 1811 18819
rect 2329 18785 2363 18819
rect 2973 18785 3007 18819
rect 4813 18717 4847 18751
rect 16190 18853 16224 18887
rect 6285 18785 6319 18819
rect 9505 18785 9539 18819
rect 10333 18785 10367 18819
rect 11529 18785 11563 18819
rect 12081 18785 12115 18819
rect 12348 18785 12382 18819
rect 13737 18785 13771 18819
rect 14565 18785 14599 18819
rect 15301 18785 15335 18819
rect 17601 18785 17635 18819
rect 17868 18785 17902 18819
rect 19073 18785 19107 18819
rect 19257 18785 19291 18819
rect 20269 18785 20303 18819
rect 6377 18717 6411 18751
rect 6469 18717 6503 18751
rect 8401 18717 8435 18751
rect 8585 18717 8619 18751
rect 10425 18717 10459 18751
rect 10609 18717 10643 18751
rect 11069 18717 11103 18751
rect 14657 18717 14691 18751
rect 14841 18717 14875 18751
rect 15945 18717 15979 18751
rect 19533 18717 19567 18751
rect 20913 18717 20947 18751
rect 5825 18649 5859 18683
rect 9965 18649 9999 18683
rect 11713 18649 11747 18683
rect 14197 18649 14231 18683
rect 17325 18649 17359 18683
rect 18981 18649 19015 18683
rect 19073 18649 19107 18683
rect 5917 18581 5951 18615
rect 7941 18581 7975 18615
rect 1777 18377 1811 18411
rect 3065 18377 3099 18411
rect 6837 18377 6871 18411
rect 11069 18377 11103 18411
rect 12541 18377 12575 18411
rect 15945 18377 15979 18411
rect 16497 18377 16531 18411
rect 17049 18377 17083 18411
rect 17601 18377 17635 18411
rect 18061 18377 18095 18411
rect 19625 18377 19659 18411
rect 5641 18309 5675 18343
rect 13461 18309 13495 18343
rect 20913 18309 20947 18343
rect 7297 18241 7331 18275
rect 7481 18241 7515 18275
rect 9689 18241 9723 18275
rect 11989 18241 12023 18275
rect 12173 18241 12207 18275
rect 13001 18241 13035 18275
rect 13185 18241 13219 18275
rect 1593 18173 1627 18207
rect 2145 18173 2179 18207
rect 2421 18173 2455 18207
rect 2881 18173 2915 18207
rect 3433 18173 3467 18207
rect 4261 18173 4295 18207
rect 7205 18173 7239 18207
rect 8033 18173 8067 18207
rect 4528 18105 4562 18139
rect 8300 18105 8334 18139
rect 9956 18105 9990 18139
rect 11805 18105 11839 18139
rect 14105 18241 14139 18275
rect 14565 18241 14599 18275
rect 18705 18241 18739 18275
rect 16313 18173 16347 18207
rect 16865 18173 16899 18207
rect 17417 18173 17451 18207
rect 18429 18173 18463 18207
rect 19441 18173 19475 18207
rect 19993 18173 20027 18207
rect 20729 18173 20763 18207
rect 12909 18105 12943 18139
rect 13461 18105 13495 18139
rect 13921 18105 13955 18139
rect 14832 18105 14866 18139
rect 20269 18105 20303 18139
rect 3617 18037 3651 18071
rect 9413 18037 9447 18071
rect 11345 18037 11379 18071
rect 11713 18037 11747 18071
rect 12173 18037 12207 18071
rect 13553 18037 13587 18071
rect 14013 18037 14047 18071
rect 18521 18037 18555 18071
rect 3065 17833 3099 17867
rect 7021 17833 7055 17867
rect 7481 17833 7515 17867
rect 11897 17833 11931 17867
rect 13829 17833 13863 17867
rect 14197 17833 14231 17867
rect 14657 17833 14691 17867
rect 15301 17833 15335 17867
rect 10508 17765 10542 17799
rect 16589 17765 16623 17799
rect 18236 17765 18270 17799
rect 20269 17765 20303 17799
rect 1593 17697 1627 17731
rect 2155 17697 2189 17731
rect 2881 17697 2915 17731
rect 4721 17697 4755 17731
rect 5632 17697 5666 17731
rect 7389 17697 7423 17731
rect 8953 17697 8987 17731
rect 10241 17697 10275 17731
rect 12449 17697 12483 17731
rect 12716 17697 12750 17731
rect 14565 17697 14599 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 16313 17697 16347 17731
rect 17417 17697 17451 17731
rect 19993 17697 20027 17731
rect 2329 17629 2363 17663
rect 4813 17629 4847 17663
rect 4997 17629 5031 17663
rect 5365 17629 5399 17663
rect 7573 17629 7607 17663
rect 9045 17629 9079 17663
rect 9229 17629 9263 17663
rect 14841 17629 14875 17663
rect 15853 17629 15887 17663
rect 17969 17629 18003 17663
rect 8585 17561 8619 17595
rect 1777 17493 1811 17527
rect 4353 17493 4387 17527
rect 6745 17493 6779 17527
rect 11621 17493 11655 17527
rect 17601 17493 17635 17527
rect 19349 17493 19383 17527
rect 2513 17289 2547 17323
rect 4629 17289 4663 17323
rect 5641 17289 5675 17323
rect 9321 17289 9355 17323
rect 10333 17289 10367 17323
rect 4353 17221 4387 17255
rect 12449 17221 12483 17255
rect 13645 17221 13679 17255
rect 19625 17221 19659 17255
rect 2973 17153 3007 17187
rect 5273 17153 5307 17187
rect 6101 17153 6135 17187
rect 6285 17153 6319 17187
rect 9965 17153 9999 17187
rect 10885 17153 10919 17187
rect 11989 17153 12023 17187
rect 13093 17153 13127 17187
rect 14473 17153 14507 17187
rect 14565 17153 14599 17187
rect 18245 17153 18279 17187
rect 20637 17153 20671 17187
rect 1777 17085 1811 17119
rect 2329 17085 2363 17119
rect 5089 17085 5123 17119
rect 6009 17085 6043 17119
rect 6837 17085 6871 17119
rect 7093 17085 7127 17119
rect 9781 17085 9815 17119
rect 10701 17085 10735 17119
rect 11713 17085 11747 17119
rect 13461 17085 13495 17119
rect 15025 17085 15059 17119
rect 15853 17085 15887 17119
rect 18512 17085 18546 17119
rect 3218 17017 3252 17051
rect 9689 17017 9723 17051
rect 10793 17017 10827 17051
rect 12817 17017 12851 17051
rect 15301 17017 15335 17051
rect 16120 17017 16154 17051
rect 20453 17017 20487 17051
rect 1961 16949 1995 16983
rect 4997 16949 5031 16983
rect 8217 16949 8251 16983
rect 11345 16949 11379 16983
rect 11805 16949 11839 16983
rect 12909 16949 12943 16983
rect 14013 16949 14047 16983
rect 14381 16949 14415 16983
rect 17233 16949 17267 16983
rect 17509 16949 17543 16983
rect 19901 16949 19935 16983
rect 20085 16949 20119 16983
rect 20545 16949 20579 16983
rect 4445 16745 4479 16779
rect 4813 16745 4847 16779
rect 5917 16745 5951 16779
rect 6469 16745 6503 16779
rect 8309 16745 8343 16779
rect 10517 16745 10551 16779
rect 10977 16745 11011 16779
rect 11529 16745 11563 16779
rect 14657 16745 14691 16779
rect 15669 16745 15703 16779
rect 17417 16745 17451 16779
rect 18245 16745 18279 16779
rect 18613 16745 18647 16779
rect 18981 16745 19015 16779
rect 19625 16745 19659 16779
rect 5825 16677 5859 16711
rect 8677 16677 8711 16711
rect 10885 16677 10919 16711
rect 11989 16677 12023 16711
rect 12817 16677 12851 16711
rect 19073 16677 19107 16711
rect 1409 16609 1443 16643
rect 2228 16609 2262 16643
rect 4905 16609 4939 16643
rect 6837 16609 6871 16643
rect 8769 16609 8803 16643
rect 11897 16609 11931 16643
rect 13544 16609 13578 16643
rect 15485 16609 15519 16643
rect 16293 16609 16327 16643
rect 18061 16609 18095 16643
rect 19993 16609 20027 16643
rect 20913 16609 20947 16643
rect 1961 16541 1995 16575
rect 4997 16541 5031 16575
rect 6009 16541 6043 16575
rect 6929 16541 6963 16575
rect 7021 16541 7055 16575
rect 8861 16541 8895 16575
rect 11161 16541 11195 16575
rect 12081 16541 12115 16575
rect 13277 16541 13311 16575
rect 16037 16541 16071 16575
rect 19257 16541 19291 16575
rect 20085 16541 20119 16575
rect 20177 16541 20211 16575
rect 1593 16473 1627 16507
rect 3341 16405 3375 16439
rect 5457 16405 5491 16439
rect 3893 16201 3927 16235
rect 13461 16201 13495 16235
rect 14473 16201 14507 16235
rect 16221 16201 16255 16235
rect 17601 16201 17635 16235
rect 18429 16201 18463 16235
rect 15853 16133 15887 16167
rect 4721 16065 4755 16099
rect 5825 16065 5859 16099
rect 7573 16065 7607 16099
rect 10057 16065 10091 16099
rect 13001 16065 13035 16099
rect 14013 16065 14047 16099
rect 15025 16065 15059 16099
rect 16773 16065 16807 16099
rect 1777 15997 1811 16031
rect 2513 15997 2547 16031
rect 4629 15997 4663 16031
rect 5549 15997 5583 16031
rect 8401 15997 8435 16031
rect 8668 15997 8702 16031
rect 10324 15997 10358 16031
rect 12909 15997 12943 16031
rect 14841 15997 14875 16031
rect 15669 15997 15703 16031
rect 17417 15997 17451 16031
rect 18245 15997 18279 16031
rect 18797 15997 18831 16031
rect 19064 15997 19098 16031
rect 20453 15997 20487 16031
rect 2053 15929 2087 15963
rect 2780 15929 2814 15963
rect 4537 15929 4571 15963
rect 5641 15929 5675 15963
rect 12817 15929 12851 15963
rect 13829 15929 13863 15963
rect 14933 15929 14967 15963
rect 20729 15929 20763 15963
rect 4169 15861 4203 15895
rect 5181 15861 5215 15895
rect 7021 15861 7055 15895
rect 7389 15861 7423 15895
rect 7481 15861 7515 15895
rect 9781 15861 9815 15895
rect 11437 15861 11471 15895
rect 11897 15861 11931 15895
rect 12449 15861 12483 15895
rect 13921 15861 13955 15895
rect 16589 15861 16623 15895
rect 16681 15861 16715 15895
rect 20177 15861 20211 15895
rect 1961 15657 1995 15691
rect 2329 15657 2363 15691
rect 2789 15657 2823 15691
rect 5733 15657 5767 15691
rect 7849 15657 7883 15691
rect 8217 15657 8251 15691
rect 8861 15657 8895 15691
rect 11805 15657 11839 15691
rect 12173 15657 12207 15691
rect 15945 15657 15979 15691
rect 16497 15657 16531 15691
rect 16865 15657 16899 15691
rect 18981 15657 19015 15691
rect 4620 15589 4654 15623
rect 8309 15589 8343 15623
rect 10416 15589 10450 15623
rect 15853 15589 15887 15623
rect 18061 15589 18095 15623
rect 1777 15521 1811 15555
rect 2697 15521 2731 15555
rect 3341 15521 3375 15555
rect 6193 15521 6227 15555
rect 6460 15521 6494 15555
rect 9045 15521 9079 15555
rect 10149 15521 10183 15555
rect 12265 15521 12299 15555
rect 13185 15521 13219 15555
rect 13544 15521 13578 15555
rect 18153 15521 18187 15555
rect 19349 15521 19383 15555
rect 19993 15521 20027 15555
rect 2973 15453 3007 15487
rect 4353 15453 4387 15487
rect 8401 15453 8435 15487
rect 12357 15453 12391 15487
rect 13277 15453 13311 15487
rect 16037 15453 16071 15487
rect 16405 15453 16439 15487
rect 16957 15453 16991 15487
rect 17049 15453 17083 15487
rect 18337 15453 18371 15487
rect 19441 15453 19475 15487
rect 19533 15453 19567 15487
rect 20177 15453 20211 15487
rect 20913 15453 20947 15487
rect 3525 15385 3559 15419
rect 7573 15385 7607 15419
rect 15485 15385 15519 15419
rect 11529 15317 11563 15351
rect 13001 15317 13035 15351
rect 14657 15317 14691 15351
rect 16405 15317 16439 15351
rect 17693 15317 17727 15351
rect 2421 15113 2455 15147
rect 6285 15113 6319 15147
rect 7849 15113 7883 15147
rect 8677 15113 8711 15147
rect 12817 15113 12851 15147
rect 14565 15113 14599 15147
rect 15761 15113 15795 15147
rect 1961 15045 1995 15079
rect 6837 15045 6871 15079
rect 3065 14977 3099 15011
rect 4077 14977 4111 15011
rect 5825 14977 5859 15011
rect 6101 14977 6135 15011
rect 7297 14977 7331 15011
rect 7481 14977 7515 15011
rect 8401 14977 8435 15011
rect 1777 14909 1811 14943
rect 5733 14909 5767 14943
rect 6469 14909 6503 14943
rect 7665 14909 7699 14943
rect 2789 14841 2823 14875
rect 3801 14841 3835 14875
rect 4445 14841 4479 14875
rect 5641 14841 5675 14875
rect 6101 14841 6135 14875
rect 11345 15045 11379 15079
rect 9321 14977 9355 15011
rect 9505 14977 9539 15011
rect 10517 14977 10551 15011
rect 11989 14977 12023 15011
rect 15393 14977 15427 15011
rect 15669 14977 15703 15011
rect 9229 14909 9263 14943
rect 10333 14909 10367 14943
rect 12633 14909 12667 14943
rect 13185 14909 13219 14943
rect 11805 14841 11839 14875
rect 13452 14841 13486 14875
rect 17233 15045 17267 15079
rect 18521 15045 18555 15079
rect 15853 14977 15887 15011
rect 20729 14977 20763 15011
rect 15761 14909 15795 14943
rect 18337 14909 18371 14943
rect 18889 14909 18923 14943
rect 20545 14909 20579 14943
rect 16120 14841 16154 14875
rect 19156 14841 19190 14875
rect 2881 14773 2915 14807
rect 3433 14773 3467 14807
rect 3893 14773 3927 14807
rect 5273 14773 5307 14807
rect 7205 14773 7239 14807
rect 7665 14773 7699 14807
rect 8217 14773 8251 14807
rect 8309 14773 8343 14807
rect 8677 14773 8711 14807
rect 8861 14773 8895 14807
rect 9965 14773 9999 14807
rect 10425 14773 10459 14807
rect 11713 14773 11747 14807
rect 14841 14773 14875 14807
rect 15209 14773 15243 14807
rect 15301 14773 15335 14807
rect 15669 14773 15703 14807
rect 17509 14773 17543 14807
rect 20269 14773 20303 14807
rect 2789 14569 2823 14603
rect 8585 14569 8619 14603
rect 8953 14569 8987 14603
rect 9873 14569 9907 14603
rect 10333 14569 10367 14603
rect 12265 14569 12299 14603
rect 14841 14569 14875 14603
rect 16773 14569 16807 14603
rect 19257 14569 19291 14603
rect 19625 14569 19659 14603
rect 19993 14569 20027 14603
rect 3249 14501 3283 14535
rect 6184 14501 6218 14535
rect 15660 14501 15694 14535
rect 17325 14501 17359 14535
rect 20085 14501 20119 14535
rect 1685 14433 1719 14467
rect 3157 14433 3191 14467
rect 4333 14433 4367 14467
rect 5917 14433 5951 14467
rect 10241 14433 10275 14467
rect 11152 14433 11186 14467
rect 12889 14433 12923 14467
rect 14657 14433 14691 14467
rect 15393 14433 15427 14467
rect 17049 14433 17083 14467
rect 17877 14433 17911 14467
rect 18144 14433 18178 14467
rect 1869 14365 1903 14399
rect 3341 14365 3375 14399
rect 4077 14365 4111 14399
rect 9045 14365 9079 14399
rect 9137 14365 9171 14399
rect 10425 14365 10459 14399
rect 10885 14365 10919 14399
rect 12633 14365 12667 14399
rect 20177 14365 20211 14399
rect 5457 14297 5491 14331
rect 14013 14297 14047 14331
rect 7297 14229 7331 14263
rect 1593 14025 1627 14059
rect 1961 14025 1995 14059
rect 6837 14025 6871 14059
rect 8309 14025 8343 14059
rect 11621 14025 11655 14059
rect 12449 14025 12483 14059
rect 13737 14025 13771 14059
rect 15761 14025 15795 14059
rect 16037 14025 16071 14059
rect 18981 14025 19015 14059
rect 2973 13957 3007 13991
rect 4169 13957 4203 13991
rect 5733 13957 5767 13991
rect 13461 13957 13495 13991
rect 19993 13957 20027 13991
rect 2421 13889 2455 13923
rect 2605 13889 2639 13923
rect 3433 13889 3467 13923
rect 3525 13889 3559 13923
rect 4721 13889 4755 13923
rect 6193 13889 6227 13923
rect 6377 13889 6411 13923
rect 7481 13889 7515 13923
rect 13001 13889 13035 13923
rect 14289 13889 14323 13923
rect 15301 13889 15335 13923
rect 16497 13889 16531 13923
rect 16681 13889 16715 13923
rect 17233 13889 17267 13923
rect 19441 13889 19475 13923
rect 19625 13889 19659 13923
rect 20545 13889 20579 13923
rect 1409 13821 1443 13855
rect 4629 13821 4663 13855
rect 7205 13821 7239 13855
rect 8493 13821 8527 13855
rect 8585 13821 8619 13855
rect 8852 13821 8886 13855
rect 10241 13821 10275 13855
rect 12909 13821 12943 13855
rect 13645 13821 13679 13855
rect 15945 13821 15979 13855
rect 16405 13821 16439 13855
rect 17049 13821 17083 13855
rect 18245 13821 18279 13855
rect 18521 13821 18555 13855
rect 20453 13821 20487 13855
rect 6101 13753 6135 13787
rect 7849 13753 7883 13787
rect 10508 13753 10542 13787
rect 11897 13753 11931 13787
rect 14105 13753 14139 13787
rect 2329 13685 2363 13719
rect 3341 13685 3375 13719
rect 4537 13685 4571 13719
rect 7297 13685 7331 13719
rect 9965 13685 9999 13719
rect 12817 13685 12851 13719
rect 14197 13685 14231 13719
rect 14749 13685 14783 13719
rect 15117 13685 15151 13719
rect 15209 13685 15243 13719
rect 19349 13685 19383 13719
rect 20361 13685 20395 13719
rect 3157 13481 3191 13515
rect 3617 13481 3651 13515
rect 4077 13481 4111 13515
rect 4537 13481 4571 13515
rect 5089 13481 5123 13515
rect 5457 13481 5491 13515
rect 6193 13481 6227 13515
rect 10241 13481 10275 13515
rect 10609 13481 10643 13515
rect 10701 13481 10735 13515
rect 11253 13481 11287 13515
rect 11621 13481 11655 13515
rect 16129 13481 16163 13515
rect 16497 13481 16531 13515
rect 18521 13481 18555 13515
rect 18797 13481 18831 13515
rect 20269 13481 20303 13515
rect 6561 13413 6595 13447
rect 11713 13413 11747 13447
rect 12817 13413 12851 13447
rect 13921 13413 13955 13447
rect 15577 13413 15611 13447
rect 1777 13345 1811 13379
rect 2044 13345 2078 13379
rect 3433 13345 3467 13379
rect 4445 13345 4479 13379
rect 7389 13345 7423 13379
rect 7656 13345 7690 13379
rect 12725 13345 12759 13379
rect 13829 13345 13863 13379
rect 14657 13345 14691 13379
rect 15301 13345 15335 13379
rect 17141 13345 17175 13379
rect 17408 13345 17442 13379
rect 19165 13345 19199 13379
rect 20177 13345 20211 13379
rect 4629 13277 4663 13311
rect 5549 13277 5583 13311
rect 5641 13277 5675 13311
rect 6653 13277 6687 13311
rect 6837 13277 6871 13311
rect 10793 13277 10827 13311
rect 11897 13277 11931 13311
rect 13001 13277 13035 13311
rect 14013 13277 14047 13311
rect 16589 13277 16623 13311
rect 16681 13277 16715 13311
rect 19257 13277 19291 13311
rect 19349 13277 19383 13311
rect 20361 13277 20395 13311
rect 8769 13141 8803 13175
rect 12357 13141 12391 13175
rect 13461 13141 13495 13175
rect 14841 13141 14875 13175
rect 19809 13141 19843 13175
rect 3893 12937 3927 12971
rect 4997 12937 5031 12971
rect 12265 12937 12299 12971
rect 1869 12869 1903 12903
rect 10057 12869 10091 12903
rect 11345 12869 11379 12903
rect 2513 12801 2547 12835
rect 3433 12801 3467 12835
rect 4537 12801 4571 12835
rect 5549 12801 5583 12835
rect 7941 12801 7975 12835
rect 8677 12801 8711 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 11805 12801 11839 12835
rect 11989 12801 12023 12835
rect 2329 12733 2363 12767
rect 4261 12733 4295 12767
rect 7757 12733 7791 12767
rect 3341 12665 3375 12699
rect 4353 12665 4387 12699
rect 5365 12665 5399 12699
rect 5457 12665 5491 12699
rect 8944 12665 8978 12699
rect 11713 12665 11747 12699
rect 13829 12937 13863 12971
rect 14013 12937 14047 12971
rect 15025 12937 15059 12971
rect 17693 12937 17727 12971
rect 18061 12937 18095 12971
rect 13001 12801 13035 12835
rect 13553 12801 13587 12835
rect 12817 12733 12851 12767
rect 12909 12733 12943 12767
rect 17785 12869 17819 12903
rect 14657 12801 14691 12835
rect 15577 12801 15611 12835
rect 16313 12801 16347 12835
rect 18613 12801 18647 12835
rect 14381 12733 14415 12767
rect 15485 12733 15519 12767
rect 16580 12733 16614 12767
rect 17785 12733 17819 12767
rect 18429 12733 18463 12767
rect 19349 12733 19383 12767
rect 14473 12665 14507 12699
rect 18521 12665 18555 12699
rect 19616 12665 19650 12699
rect 2237 12597 2271 12631
rect 2881 12597 2915 12631
rect 3249 12597 3283 12631
rect 7297 12597 7331 12631
rect 7665 12597 7699 12631
rect 10333 12597 10367 12631
rect 10701 12597 10735 12631
rect 12265 12597 12299 12631
rect 12449 12597 12483 12631
rect 13829 12597 13863 12631
rect 15393 12597 15427 12631
rect 20729 12597 20763 12631
rect 2973 12393 3007 12427
rect 4445 12393 4479 12427
rect 5641 12393 5675 12427
rect 8401 12393 8435 12427
rect 10057 12393 10091 12427
rect 12633 12393 12667 12427
rect 12909 12393 12943 12427
rect 13369 12393 13403 12427
rect 13921 12393 13955 12427
rect 17141 12393 17175 12427
rect 18797 12393 18831 12427
rect 19533 12393 19567 12427
rect 3525 12325 3559 12359
rect 6009 12325 6043 12359
rect 6460 12325 6494 12359
rect 8493 12325 8527 12359
rect 13277 12325 13311 12359
rect 17684 12325 17718 12359
rect 19073 12325 19107 12359
rect 1860 12257 1894 12291
rect 3249 12257 3283 12291
rect 5549 12257 5583 12291
rect 6193 12257 6227 12291
rect 9229 12257 9263 12291
rect 11253 12257 11287 12291
rect 11520 12257 11554 12291
rect 14289 12257 14323 12291
rect 15761 12257 15795 12291
rect 16028 12257 16062 12291
rect 17417 12257 17451 12291
rect 19901 12257 19935 12291
rect 1593 12189 1627 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 5825 12189 5859 12223
rect 6009 12189 6043 12223
rect 8677 12189 8711 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 13461 12189 13495 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 19993 12189 20027 12223
rect 20177 12189 20211 12223
rect 4077 12121 4111 12155
rect 8033 12121 8067 12155
rect 5181 12053 5215 12087
rect 7573 12053 7607 12087
rect 9045 12053 9079 12087
rect 9689 12053 9723 12087
rect 1777 11849 1811 11883
rect 3341 11849 3375 11883
rect 12449 11849 12483 11883
rect 16037 11849 16071 11883
rect 17601 11849 17635 11883
rect 18061 11849 18095 11883
rect 20545 11849 20579 11883
rect 21005 11849 21039 11883
rect 4261 11781 4295 11815
rect 5733 11781 5767 11815
rect 8861 11781 8895 11815
rect 11345 11781 11379 11815
rect 2329 11713 2363 11747
rect 3801 11713 3835 11747
rect 3893 11713 3927 11747
rect 6009 11713 6043 11747
rect 7389 11713 7423 11747
rect 8401 11713 8435 11747
rect 9413 11713 9447 11747
rect 9965 11713 9999 11747
rect 12909 11713 12943 11747
rect 13093 11713 13127 11747
rect 13461 11713 13495 11747
rect 16865 11713 16899 11747
rect 18613 11713 18647 11747
rect 4353 11645 4387 11679
rect 10232 11645 10266 11679
rect 12265 11645 12299 11679
rect 12817 11645 12851 11679
rect 14657 11645 14691 11679
rect 14924 11645 14958 11679
rect 17417 11645 17451 11679
rect 18521 11645 18555 11679
rect 19165 11645 19199 11679
rect 20821 11645 20855 11679
rect 2145 11577 2179 11611
rect 3709 11577 3743 11611
rect 4261 11577 4295 11611
rect 4598 11577 4632 11611
rect 7205 11577 7239 11611
rect 9321 11577 9355 11611
rect 16773 11577 16807 11611
rect 19432 11577 19466 11611
rect 2237 11509 2271 11543
rect 6837 11509 6871 11543
rect 7297 11509 7331 11543
rect 7849 11509 7883 11543
rect 8217 11509 8251 11543
rect 8309 11509 8343 11543
rect 9229 11509 9263 11543
rect 12081 11509 12115 11543
rect 16313 11509 16347 11543
rect 16681 11509 16715 11543
rect 18429 11509 18463 11543
rect 1961 11305 1995 11339
rect 2329 11305 2363 11339
rect 2973 11305 3007 11339
rect 3433 11305 3467 11339
rect 5457 11305 5491 11339
rect 8677 11305 8711 11339
rect 11805 11305 11839 11339
rect 14565 11305 14599 11339
rect 15301 11305 15335 11339
rect 15669 11305 15703 11339
rect 16313 11305 16347 11339
rect 16681 11305 16715 11339
rect 17785 11305 17819 11339
rect 19717 11305 19751 11339
rect 4344 11237 4378 11271
rect 8769 11237 8803 11271
rect 12624 11237 12658 11271
rect 14657 11237 14691 11271
rect 16773 11237 16807 11271
rect 17693 11237 17727 11271
rect 3341 11169 3375 11203
rect 3893 11169 3927 11203
rect 6561 11169 6595 11203
rect 6920 11169 6954 11203
rect 10517 11169 10551 11203
rect 12357 11169 12391 11203
rect 18705 11169 18739 11203
rect 20085 11169 20119 11203
rect 2421 11101 2455 11135
rect 2605 11101 2639 11135
rect 3617 11101 3651 11135
rect 4077 11101 4111 11135
rect 6653 11101 6687 11135
rect 8861 11101 8895 11135
rect 14841 11101 14875 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 16957 11101 16991 11135
rect 17877 11101 17911 11135
rect 18797 11101 18831 11135
rect 18889 11101 18923 11135
rect 20177 11101 20211 11135
rect 20269 11101 20303 11135
rect 6377 11033 6411 11067
rect 8033 11033 8067 11067
rect 14197 11033 14231 11067
rect 3893 10965 3927 10999
rect 8309 10965 8343 10999
rect 13737 10965 13771 10999
rect 17325 10965 17359 10999
rect 18337 10965 18371 10999
rect 3893 10761 3927 10795
rect 16221 10761 16255 10795
rect 16497 10761 16531 10795
rect 18337 10761 18371 10795
rect 19901 10761 19935 10795
rect 20361 10761 20395 10795
rect 4997 10693 5031 10727
rect 8033 10693 8067 10727
rect 11069 10693 11103 10727
rect 2145 10625 2179 10659
rect 4445 10625 4479 10659
rect 6285 10625 6319 10659
rect 7573 10625 7607 10659
rect 8677 10625 8711 10659
rect 9413 10625 9447 10659
rect 9689 10625 9723 10659
rect 11713 10625 11747 10659
rect 13001 10625 13035 10659
rect 14289 10625 14323 10659
rect 14473 10625 14507 10659
rect 14841 10625 14875 10659
rect 16957 10625 16991 10659
rect 17049 10625 17083 10659
rect 20913 10625 20947 10659
rect 4353 10557 4387 10591
rect 5181 10557 5215 10591
rect 8401 10557 8435 10591
rect 8493 10557 8527 10591
rect 9321 10557 9355 10591
rect 11529 10557 11563 10591
rect 12817 10557 12851 10591
rect 13737 10557 13771 10591
rect 15097 10557 15131 10591
rect 16865 10557 16899 10591
rect 18153 10557 18187 10591
rect 18521 10557 18555 10591
rect 2412 10489 2446 10523
rect 7389 10489 7423 10523
rect 9229 10489 9263 10523
rect 9956 10489 9990 10523
rect 11621 10489 11655 10523
rect 14197 10489 14231 10523
rect 17509 10489 17543 10523
rect 18788 10489 18822 10523
rect 20821 10489 20855 10523
rect 1685 10421 1719 10455
rect 3525 10421 3559 10455
rect 4261 10421 4295 10455
rect 5733 10421 5767 10455
rect 6101 10421 6135 10455
rect 6193 10421 6227 10455
rect 6929 10421 6963 10455
rect 7297 10421 7331 10455
rect 8861 10421 8895 10455
rect 11161 10421 11195 10455
rect 12449 10421 12483 10455
rect 12909 10421 12943 10455
rect 13553 10421 13587 10455
rect 13829 10421 13863 10455
rect 20177 10421 20211 10455
rect 20729 10421 20763 10455
rect 2329 10217 2363 10251
rect 2421 10217 2455 10251
rect 2973 10217 3007 10251
rect 6837 10217 6871 10251
rect 7205 10217 7239 10251
rect 7297 10217 7331 10251
rect 7849 10217 7883 10251
rect 8217 10217 8251 10251
rect 8861 10217 8895 10251
rect 11069 10217 11103 10251
rect 11805 10217 11839 10251
rect 12357 10217 12391 10251
rect 13001 10217 13035 10251
rect 13369 10217 13403 10251
rect 15761 10217 15795 10251
rect 17785 10217 17819 10251
rect 18429 10217 18463 10251
rect 19809 10217 19843 10251
rect 20913 10217 20947 10251
rect 4782 10149 4816 10183
rect 11529 10149 11563 10183
rect 15669 10149 15703 10183
rect 3341 10081 3375 10115
rect 3433 10081 3467 10115
rect 4537 10081 4571 10115
rect 7665 10081 7699 10115
rect 8309 10081 8343 10115
rect 9045 10081 9079 10115
rect 9689 10081 9723 10115
rect 9956 10081 9990 10115
rect 11805 10081 11839 10115
rect 12449 10081 12483 10115
rect 14381 10081 14415 10115
rect 16405 10081 16439 10115
rect 16672 10081 16706 10115
rect 18797 10081 18831 10115
rect 2605 10013 2639 10047
rect 3617 10013 3651 10047
rect 7481 10013 7515 10047
rect 1961 9945 1995 9979
rect 8401 10013 8435 10047
rect 12541 10013 12575 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 14473 10013 14507 10047
rect 14565 10013 14599 10047
rect 15853 10013 15887 10047
rect 18889 10013 18923 10047
rect 19073 10013 19107 10047
rect 19901 10013 19935 10047
rect 19993 10013 20027 10047
rect 19441 9945 19475 9979
rect 5917 9877 5951 9911
rect 7665 9877 7699 9911
rect 11989 9877 12023 9911
rect 14013 9877 14047 9911
rect 15301 9877 15335 9911
rect 8217 9673 8251 9707
rect 16865 9673 16899 9707
rect 1869 9605 1903 9639
rect 2237 9605 2271 9639
rect 13369 9605 13403 9639
rect 2881 9537 2915 9571
rect 4353 9537 4387 9571
rect 10241 9537 10275 9571
rect 10977 9537 11011 9571
rect 13001 9537 13035 9571
rect 1685 9469 1719 9503
rect 4721 9469 4755 9503
rect 4988 9469 5022 9503
rect 6837 9469 6871 9503
rect 8769 9469 8803 9503
rect 2605 9401 2639 9435
rect 4077 9401 4111 9435
rect 7082 9401 7116 9435
rect 9014 9401 9048 9435
rect 10793 9469 10827 9503
rect 14013 9537 14047 9571
rect 14933 9537 14967 9571
rect 15117 9537 15151 9571
rect 15669 9537 15703 9571
rect 19625 9605 19659 9639
rect 19993 9605 20027 9639
rect 17417 9537 17451 9571
rect 17601 9537 17635 9571
rect 20545 9537 20579 9571
rect 13829 9469 13863 9503
rect 14841 9469 14875 9503
rect 15485 9469 15519 9503
rect 16405 9469 16439 9503
rect 16865 9469 16899 9503
rect 17325 9469 17359 9503
rect 18245 9469 18279 9503
rect 10885 9401 10919 9435
rect 12817 9401 12851 9435
rect 13369 9401 13403 9435
rect 18512 9401 18546 9435
rect 20453 9401 20487 9435
rect 2697 9333 2731 9367
rect 3709 9333 3743 9367
rect 4169 9333 4203 9367
rect 6101 9333 6135 9367
rect 10149 9333 10183 9367
rect 10241 9333 10275 9367
rect 10425 9333 10459 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 13461 9333 13495 9367
rect 13921 9333 13955 9367
rect 14473 9333 14507 9367
rect 16221 9333 16255 9367
rect 16957 9333 16991 9367
rect 20361 9333 20395 9367
rect 3617 9129 3651 9163
rect 5917 9129 5951 9163
rect 6837 9129 6871 9163
rect 12265 9129 12299 9163
rect 13277 9129 13311 9163
rect 17509 9129 17543 9163
rect 17877 9129 17911 9163
rect 19257 9129 19291 9163
rect 1777 9061 1811 9095
rect 7564 9061 7598 9095
rect 9956 9061 9990 9095
rect 13645 9061 13679 9095
rect 14565 9061 14599 9095
rect 19349 9061 19383 9095
rect 1501 8993 1535 9027
rect 2237 8993 2271 9027
rect 2504 8993 2538 9027
rect 4905 8993 4939 9027
rect 7297 8993 7331 9027
rect 9689 8993 9723 9027
rect 12173 8993 12207 9027
rect 12633 8993 12667 9027
rect 12725 8993 12759 9027
rect 13737 8993 13771 9027
rect 14289 8993 14323 9027
rect 16129 8993 16163 9027
rect 16396 8993 16430 9027
rect 18245 8993 18279 9027
rect 18337 8993 18371 9027
rect 20085 8993 20119 9027
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 6009 8925 6043 8959
rect 6101 8925 6135 8959
rect 12909 8925 12943 8959
rect 13829 8925 13863 8959
rect 18521 8925 18555 8959
rect 19441 8925 19475 8959
rect 20269 8925 20303 8959
rect 4537 8857 4571 8891
rect 18889 8857 18923 8891
rect 5549 8789 5583 8823
rect 8677 8789 8711 8823
rect 11069 8789 11103 8823
rect 11989 8789 12023 8823
rect 3065 8585 3099 8619
rect 4905 8585 4939 8619
rect 9597 8585 9631 8619
rect 16313 8585 16347 8619
rect 20177 8585 20211 8619
rect 20729 8585 20763 8619
rect 4077 8517 4111 8551
rect 10609 8517 10643 8551
rect 14381 8517 14415 8551
rect 14565 8517 14599 8551
rect 4537 8449 4571 8483
rect 4721 8449 4755 8483
rect 4905 8449 4939 8483
rect 5641 8449 5675 8483
rect 10149 8449 10183 8483
rect 11069 8449 11103 8483
rect 11161 8449 11195 8483
rect 13001 8449 13035 8483
rect 1685 8381 1719 8415
rect 1952 8381 1986 8415
rect 5457 8381 5491 8415
rect 10057 8381 10091 8415
rect 13268 8381 13302 8415
rect 14657 8449 14691 8483
rect 16957 8449 16991 8483
rect 18797 8449 18831 8483
rect 20545 8381 20579 8415
rect 4445 8313 4479 8347
rect 9965 8313 9999 8347
rect 14565 8313 14599 8347
rect 14902 8313 14936 8347
rect 16681 8313 16715 8347
rect 19064 8313 19098 8347
rect 5089 8245 5123 8279
rect 5549 8245 5583 8279
rect 10977 8245 11011 8279
rect 16037 8245 16071 8279
rect 16773 8245 16807 8279
rect 2605 8041 2639 8075
rect 2973 8041 3007 8075
rect 5549 8041 5583 8075
rect 5825 8041 5859 8075
rect 10241 8041 10275 8075
rect 12541 8041 12575 8075
rect 13001 8041 13035 8075
rect 14105 8041 14139 8075
rect 14565 8041 14599 8075
rect 17693 8041 17727 8075
rect 3065 7973 3099 8007
rect 6285 7973 6319 8007
rect 10333 7973 10367 8007
rect 12909 7973 12943 8007
rect 16282 7973 16316 8007
rect 19248 7973 19282 8007
rect 4169 7905 4203 7939
rect 4436 7905 4470 7939
rect 6193 7905 6227 7939
rect 10885 7905 10919 7939
rect 11152 7905 11186 7939
rect 14473 7905 14507 7939
rect 18061 7905 18095 7939
rect 18153 7905 18187 7939
rect 18981 7905 19015 7939
rect 3157 7837 3191 7871
rect 6377 7837 6411 7871
rect 10517 7837 10551 7871
rect 13093 7837 13127 7871
rect 14657 7837 14691 7871
rect 16037 7837 16071 7871
rect 18245 7837 18279 7871
rect 20913 7837 20947 7871
rect 17417 7769 17451 7803
rect 9873 7701 9907 7735
rect 12265 7701 12299 7735
rect 20361 7701 20395 7735
rect 3985 7497 4019 7531
rect 11713 7497 11747 7531
rect 15485 7497 15519 7531
rect 16221 7497 16255 7531
rect 18061 7497 18095 7531
rect 20453 7497 20487 7531
rect 13829 7429 13863 7463
rect 4629 7361 4663 7395
rect 4997 7361 5031 7395
rect 10333 7361 10367 7395
rect 16865 7361 16899 7395
rect 18613 7361 18647 7395
rect 19073 7361 19107 7395
rect 12449 7293 12483 7327
rect 14105 7293 14139 7327
rect 14361 7293 14395 7327
rect 18521 7293 18555 7327
rect 10600 7225 10634 7259
rect 12694 7225 12728 7259
rect 19340 7225 19374 7259
rect 4353 7157 4387 7191
rect 4445 7157 4479 7191
rect 16589 7157 16623 7191
rect 16681 7157 16715 7191
rect 17509 7157 17543 7191
rect 18429 7157 18463 7191
rect 11621 6953 11655 6987
rect 12173 6953 12207 6987
rect 12633 6953 12667 6987
rect 13185 6953 13219 6987
rect 13645 6953 13679 6987
rect 14197 6953 14231 6987
rect 14565 6953 14599 6987
rect 15301 6953 15335 6987
rect 15761 6953 15795 6987
rect 18061 6953 18095 6987
rect 20177 6953 20211 6987
rect 13553 6885 13587 6919
rect 16773 6885 16807 6919
rect 11529 6817 11563 6851
rect 12541 6817 12575 6851
rect 15669 6817 15703 6851
rect 16681 6817 16715 6851
rect 11805 6749 11839 6783
rect 12725 6749 12759 6783
rect 13737 6749 13771 6783
rect 14657 6749 14691 6783
rect 14841 6749 14875 6783
rect 15945 6749 15979 6783
rect 16865 6749 16899 6783
rect 18153 6749 18187 6783
rect 18337 6749 18371 6783
rect 20269 6749 20303 6783
rect 20453 6749 20487 6783
rect 16313 6681 16347 6715
rect 17693 6681 17727 6715
rect 19809 6681 19843 6715
rect 11161 6613 11195 6647
rect 10977 6409 11011 6443
rect 12449 6409 12483 6443
rect 14841 6409 14875 6443
rect 16497 6409 16531 6443
rect 20085 6409 20119 6443
rect 11621 6273 11655 6307
rect 13093 6273 13127 6307
rect 14381 6273 14415 6307
rect 15301 6273 15335 6307
rect 15485 6273 15519 6307
rect 17049 6273 17083 6307
rect 20637 6273 20671 6307
rect 11345 6205 11379 6239
rect 12909 6205 12943 6239
rect 16865 6205 16899 6239
rect 12817 6137 12851 6171
rect 11437 6069 11471 6103
rect 15209 6069 15243 6103
rect 16957 6069 16991 6103
rect 19901 6069 19935 6103
rect 20453 6069 20487 6103
rect 20545 6069 20579 6103
rect 10333 5865 10367 5899
rect 11612 5797 11646 5831
rect 10701 5729 10735 5763
rect 10793 5661 10827 5695
rect 10977 5661 11011 5695
rect 11345 5661 11379 5695
rect 12725 5525 12759 5559
rect 11345 5321 11379 5355
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 11713 5049 11747 5083
rect 12449 5049 12483 5083
rect 12081 3689 12115 3723
rect 10968 3621 11002 3655
rect 10701 3553 10735 3587
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2774 20040 2780 20052
rect 1995 20012 2780 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 12161 20043 12219 20049
rect 12161 20009 12173 20043
rect 12207 20040 12219 20043
rect 13446 20040 13452 20052
rect 12207 20012 13452 20040
rect 12207 20009 12219 20012
rect 12161 20003 12219 20009
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13964 20012 14105 20040
rect 13964 20000 13970 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 14093 20003 14151 20009
rect 14458 20000 14464 20052
rect 14516 20040 14522 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 14516 20012 15025 20040
rect 14516 20000 14522 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15841 20043 15899 20049
rect 15841 20040 15853 20043
rect 15436 20012 15853 20040
rect 15436 20000 15442 20012
rect 15841 20009 15853 20012
rect 15887 20009 15899 20043
rect 15841 20003 15899 20009
rect 15930 20000 15936 20052
rect 15988 20040 15994 20052
rect 16393 20043 16451 20049
rect 16393 20040 16405 20043
rect 15988 20012 16405 20040
rect 15988 20000 15994 20012
rect 16393 20009 16405 20012
rect 16439 20009 16451 20043
rect 16393 20003 16451 20009
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 17770 20040 17776 20052
rect 17175 20012 17776 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 17865 20043 17923 20049
rect 17865 20009 17877 20043
rect 17911 20040 17923 20043
rect 18230 20040 18236 20052
rect 17911 20012 18236 20040
rect 17911 20009 17923 20012
rect 17865 20003 17923 20009
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 6638 19972 6644 19984
rect 1780 19944 6644 19972
rect 1780 19913 1808 19944
rect 6638 19932 6644 19944
rect 6696 19932 6702 19984
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 1765 19867 1823 19873
rect 2323 19907 2381 19913
rect 2323 19873 2335 19907
rect 2369 19873 2381 19907
rect 2323 19867 2381 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19873 2927 19907
rect 2869 19867 2927 19873
rect 2332 19768 2360 19867
rect 2884 19836 2912 19867
rect 3142 19864 3148 19916
rect 3200 19904 3206 19916
rect 3421 19907 3479 19913
rect 3421 19904 3433 19907
rect 3200 19876 3433 19904
rect 3200 19864 3206 19876
rect 3421 19873 3433 19876
rect 3467 19873 3479 19907
rect 11974 19904 11980 19916
rect 11935 19876 11980 19904
rect 3421 19867 3479 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12894 19864 12900 19916
rect 12952 19904 12958 19916
rect 13081 19907 13139 19913
rect 13081 19904 13093 19907
rect 12952 19876 13093 19904
rect 12952 19864 12958 19876
rect 13081 19873 13093 19876
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 13173 19907 13231 19913
rect 13173 19873 13185 19907
rect 13219 19904 13231 19907
rect 13538 19904 13544 19916
rect 13219 19876 13544 19904
rect 13219 19873 13231 19876
rect 13173 19867 13231 19873
rect 3234 19836 3240 19848
rect 2884 19808 3240 19836
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 12158 19796 12164 19848
rect 12216 19836 12222 19848
rect 13188 19836 13216 19867
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 13909 19907 13967 19913
rect 13909 19873 13921 19907
rect 13955 19904 13967 19907
rect 14090 19904 14096 19916
rect 13955 19876 14096 19904
rect 13955 19873 13967 19876
rect 13909 19867 13967 19873
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19904 14887 19907
rect 15470 19904 15476 19916
rect 14875 19876 15476 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19873 15715 19907
rect 15657 19867 15715 19873
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19873 16267 19907
rect 16209 19867 16267 19873
rect 13354 19836 13360 19848
rect 12216 19808 13216 19836
rect 13315 19808 13360 19836
rect 12216 19796 12222 19808
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 3326 19768 3332 19780
rect 2332 19740 3332 19768
rect 3326 19728 3332 19740
rect 3384 19728 3390 19780
rect 15672 19768 15700 19867
rect 16224 19836 16252 19867
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 16632 19876 16957 19904
rect 16632 19864 16638 19876
rect 16945 19873 16957 19876
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 17310 19836 17316 19848
rect 16224 19808 17316 19836
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 17696 19836 17724 19867
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18325 19907 18383 19913
rect 18325 19904 18337 19907
rect 18012 19876 18337 19904
rect 18012 19864 18018 19876
rect 18325 19873 18337 19876
rect 18371 19873 18383 19907
rect 18325 19867 18383 19873
rect 19429 19907 19487 19913
rect 19429 19873 19441 19907
rect 19475 19904 19487 19907
rect 19886 19904 19892 19916
rect 19475 19876 19892 19904
rect 19475 19873 19487 19876
rect 19429 19867 19487 19873
rect 19886 19864 19892 19876
rect 19944 19864 19950 19916
rect 19978 19864 19984 19916
rect 20036 19904 20042 19916
rect 20533 19907 20591 19913
rect 20036 19876 20081 19904
rect 20036 19864 20042 19876
rect 20533 19873 20545 19907
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 18509 19839 18567 19845
rect 18509 19836 18521 19839
rect 17696 19808 18521 19836
rect 18509 19805 18521 19808
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20548 19836 20576 19867
rect 19852 19808 20576 19836
rect 19852 19796 19858 19808
rect 17126 19768 17132 19780
rect 15672 19740 17132 19768
rect 17126 19728 17132 19740
rect 17184 19728 17190 19780
rect 19610 19768 19616 19780
rect 19571 19740 19616 19768
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 2498 19700 2504 19712
rect 2459 19672 2504 19700
rect 2498 19660 2504 19672
rect 2556 19660 2562 19712
rect 3053 19703 3111 19709
rect 3053 19669 3065 19703
rect 3099 19700 3111 19703
rect 3418 19700 3424 19712
rect 3099 19672 3424 19700
rect 3099 19669 3111 19672
rect 3053 19663 3111 19669
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 3602 19700 3608 19712
rect 3563 19672 3608 19700
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 12710 19700 12716 19712
rect 12671 19672 12716 19700
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 3694 19496 3700 19508
rect 3655 19468 3700 19496
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 3786 19456 3792 19508
rect 3844 19496 3850 19508
rect 4249 19499 4307 19505
rect 4249 19496 4261 19499
rect 3844 19468 4261 19496
rect 3844 19456 3850 19468
rect 4249 19465 4261 19468
rect 4295 19465 4307 19499
rect 4249 19459 4307 19465
rect 16945 19499 17003 19505
rect 16945 19465 16957 19499
rect 16991 19496 17003 19499
rect 17773 19499 17831 19505
rect 17773 19496 17785 19499
rect 16991 19468 17785 19496
rect 16991 19465 17003 19468
rect 16945 19459 17003 19465
rect 17773 19465 17785 19468
rect 17819 19465 17831 19499
rect 17773 19459 17831 19465
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18049 19499 18107 19505
rect 18049 19496 18061 19499
rect 18012 19468 18061 19496
rect 18012 19456 18018 19468
rect 18049 19465 18061 19468
rect 18095 19465 18107 19499
rect 18049 19459 18107 19465
rect 2774 19388 2780 19440
rect 2832 19428 2838 19440
rect 5810 19428 5816 19440
rect 2832 19400 4200 19428
rect 2832 19388 2838 19400
rect 3694 19360 3700 19372
rect 2792 19332 3700 19360
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19261 1823 19295
rect 2590 19292 2596 19304
rect 2551 19264 2596 19292
rect 1765 19255 1823 19261
rect 1780 19224 1808 19255
rect 2590 19252 2596 19264
rect 2648 19252 2654 19304
rect 2792 19224 2820 19332
rect 3694 19320 3700 19332
rect 3752 19320 3758 19372
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 3786 19292 3792 19304
rect 3559 19264 3792 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 3878 19252 3884 19304
rect 3936 19252 3942 19304
rect 4065 19295 4123 19301
rect 4065 19261 4077 19295
rect 4111 19261 4123 19295
rect 4172 19292 4200 19400
rect 4632 19400 5816 19428
rect 4522 19292 4528 19304
rect 4172 19264 4528 19292
rect 4065 19255 4123 19261
rect 1780 19196 2820 19224
rect 2777 19159 2835 19165
rect 2777 19125 2789 19159
rect 2823 19156 2835 19159
rect 2866 19156 2872 19168
rect 2823 19128 2872 19156
rect 2823 19125 2835 19128
rect 2777 19119 2835 19125
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 3050 19116 3056 19168
rect 3108 19156 3114 19168
rect 3602 19156 3608 19168
rect 3108 19128 3608 19156
rect 3108 19116 3114 19128
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3896 19156 3924 19252
rect 4080 19224 4108 19255
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 4632 19301 4660 19400
rect 5810 19388 5816 19400
rect 5868 19388 5874 19440
rect 19978 19428 19984 19440
rect 15120 19400 19984 19428
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 8938 19360 8944 19372
rect 4764 19332 8944 19360
rect 4764 19320 4770 19332
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 11701 19363 11759 19369
rect 9784 19332 11551 19360
rect 4617 19295 4675 19301
rect 4617 19261 4629 19295
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 4798 19252 4804 19304
rect 4856 19292 4862 19304
rect 9784 19292 9812 19332
rect 4856 19264 9812 19292
rect 4856 19252 4862 19264
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 10505 19295 10563 19301
rect 10505 19292 10517 19295
rect 9916 19264 10517 19292
rect 9916 19252 9922 19264
rect 10505 19261 10517 19264
rect 10551 19261 10563 19295
rect 11422 19292 11428 19304
rect 10505 19255 10563 19261
rect 10704 19264 11284 19292
rect 11383 19264 11428 19292
rect 10704 19224 10732 19264
rect 4080 19196 10732 19224
rect 10781 19227 10839 19233
rect 10781 19193 10793 19227
rect 10827 19193 10839 19227
rect 11256 19224 11284 19264
rect 11422 19252 11428 19264
rect 11480 19252 11486 19304
rect 11523 19292 11551 19332
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 11974 19360 11980 19372
rect 11747 19332 11980 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12158 19320 12164 19372
rect 12216 19320 12222 19372
rect 12894 19360 12900 19372
rect 12360 19332 12900 19360
rect 12176 19292 12204 19320
rect 12360 19292 12388 19332
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 11523 19264 12204 19292
rect 12268 19264 12388 19292
rect 12437 19295 12495 19301
rect 12268 19224 12296 19264
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 13170 19252 13176 19304
rect 13228 19292 13234 19304
rect 13228 19264 13273 19292
rect 13228 19252 13234 19264
rect 14182 19252 14188 19304
rect 14240 19292 14246 19304
rect 14826 19292 14832 19304
rect 14240 19264 14832 19292
rect 14240 19252 14246 19264
rect 14826 19252 14832 19264
rect 14884 19252 14890 19304
rect 14918 19252 14924 19304
rect 14976 19292 14982 19304
rect 15120 19292 15148 19400
rect 19978 19388 19984 19400
rect 20036 19388 20042 19440
rect 15746 19360 15752 19372
rect 15707 19332 15752 19360
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19360 17647 19363
rect 17862 19360 17868 19372
rect 17635 19332 17868 19360
rect 17635 19329 17647 19332
rect 17589 19323 17647 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19360 18659 19363
rect 18966 19360 18972 19372
rect 18647 19332 18972 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 16117 19295 16175 19301
rect 16117 19292 16129 19295
rect 14976 19264 15148 19292
rect 15212 19264 16129 19292
rect 14976 19252 14982 19264
rect 11256 19196 12296 19224
rect 12713 19227 12771 19233
rect 10781 19187 10839 19193
rect 12713 19193 12725 19227
rect 12759 19224 12771 19227
rect 13262 19224 13268 19236
rect 12759 19196 13268 19224
rect 12759 19193 12771 19196
rect 12713 19187 12771 19193
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 3896 19128 4813 19156
rect 4801 19125 4813 19128
rect 4847 19125 4859 19159
rect 4801 19119 4859 19125
rect 4982 19116 4988 19168
rect 5040 19156 5046 19168
rect 10502 19156 10508 19168
rect 5040 19128 10508 19156
rect 5040 19116 5046 19128
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 10796 19156 10824 19187
rect 13262 19184 13268 19196
rect 13320 19184 13326 19236
rect 13446 19233 13452 19236
rect 13440 19187 13452 19233
rect 13504 19224 13510 19236
rect 15212 19224 15240 19264
rect 16117 19261 16129 19264
rect 16163 19261 16175 19295
rect 16117 19255 16175 19261
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19292 16451 19295
rect 16574 19292 16580 19304
rect 16439 19264 16580 19292
rect 16439 19261 16451 19264
rect 16393 19255 16451 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 16675 19264 18644 19292
rect 16675 19224 16703 19264
rect 17405 19227 17463 19233
rect 17405 19224 17417 19227
rect 13504 19196 13540 19224
rect 13648 19196 15056 19224
rect 13446 19184 13452 19187
rect 13504 19184 13510 19196
rect 13648 19156 13676 19196
rect 15028 19168 15056 19196
rect 15120 19196 15240 19224
rect 15292 19196 16703 19224
rect 16776 19196 17417 19224
rect 10796 19128 13676 19156
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 14608 19128 14653 19156
rect 14608 19116 14614 19128
rect 15010 19116 15016 19168
rect 15068 19116 15074 19168
rect 15120 19165 15148 19196
rect 15105 19159 15163 19165
rect 15105 19125 15117 19159
rect 15151 19125 15163 19159
rect 15105 19119 15163 19125
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15292 19156 15320 19196
rect 15252 19128 15320 19156
rect 15252 19116 15258 19128
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 15473 19159 15531 19165
rect 15473 19156 15485 19159
rect 15436 19128 15485 19156
rect 15436 19116 15442 19128
rect 15473 19125 15485 19128
rect 15519 19125 15531 19159
rect 15473 19119 15531 19125
rect 15562 19116 15568 19168
rect 15620 19156 15626 19168
rect 15620 19128 15665 19156
rect 15620 19116 15626 19128
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16776 19156 16804 19196
rect 17405 19193 17417 19196
rect 17451 19193 17463 19227
rect 17405 19187 17463 19193
rect 17773 19227 17831 19233
rect 17773 19193 17785 19227
rect 17819 19224 17831 19227
rect 18509 19227 18567 19233
rect 18509 19224 18521 19227
rect 17819 19196 18521 19224
rect 17819 19193 17831 19196
rect 17773 19187 17831 19193
rect 18509 19193 18521 19196
rect 18555 19193 18567 19227
rect 18616 19224 18644 19264
rect 18690 19252 18696 19304
rect 18748 19292 18754 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 18748 19264 19073 19292
rect 18748 19252 18754 19264
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19061 19255 19119 19261
rect 19159 19264 19993 19292
rect 19159 19224 19187 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 20346 19252 20352 19304
rect 20404 19292 20410 19304
rect 20533 19295 20591 19301
rect 20533 19292 20545 19295
rect 20404 19264 20545 19292
rect 20404 19252 20410 19264
rect 20533 19261 20545 19264
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 19334 19224 19340 19236
rect 18616 19196 19187 19224
rect 19295 19196 19340 19224
rect 18509 19187 18567 19193
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 16172 19128 16804 19156
rect 17313 19159 17371 19165
rect 16172 19116 16178 19128
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17586 19156 17592 19168
rect 17359 19128 17592 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17586 19116 17592 19128
rect 17644 19116 17650 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18417 19159 18475 19165
rect 18417 19156 18429 19159
rect 18012 19128 18429 19156
rect 18012 19116 18018 19128
rect 18417 19125 18429 19128
rect 18463 19125 18475 19159
rect 18417 19119 18475 19125
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 19300 19128 20177 19156
rect 19300 19116 19306 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20165 19119 20223 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 2501 18955 2559 18961
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 2958 18952 2964 18964
rect 2547 18924 2964 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 2958 18912 2964 18924
rect 3016 18912 3022 18964
rect 3050 18912 3056 18964
rect 3108 18952 3114 18964
rect 5813 18955 5871 18961
rect 5813 18952 5825 18955
rect 3108 18924 5825 18952
rect 3108 18912 3114 18924
rect 5813 18921 5825 18924
rect 5859 18921 5871 18955
rect 5813 18915 5871 18921
rect 7374 18912 7380 18964
rect 7432 18912 7438 18964
rect 8294 18952 8300 18964
rect 8207 18924 8300 18952
rect 8294 18912 8300 18924
rect 8352 18952 8358 18964
rect 8754 18952 8760 18964
rect 8352 18924 8760 18952
rect 8352 18912 8358 18924
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 9493 18955 9551 18961
rect 9493 18921 9505 18955
rect 9539 18952 9551 18955
rect 10962 18952 10968 18964
rect 9539 18924 10968 18952
rect 9539 18921 9551 18924
rect 9493 18915 9551 18921
rect 10962 18912 10968 18924
rect 11020 18912 11026 18964
rect 13446 18952 13452 18964
rect 11992 18924 13308 18952
rect 13407 18924 13452 18952
rect 2590 18844 2596 18896
rect 2648 18884 2654 18896
rect 3237 18887 3295 18893
rect 3237 18884 3249 18887
rect 2648 18856 3249 18884
rect 2648 18844 2654 18856
rect 3237 18853 3249 18856
rect 3283 18853 3295 18887
rect 3237 18847 3295 18853
rect 3694 18844 3700 18896
rect 3752 18884 3758 18896
rect 4982 18884 4988 18896
rect 3752 18856 4988 18884
rect 3752 18844 3758 18856
rect 4982 18844 4988 18856
rect 5040 18844 5046 18896
rect 7392 18884 7420 18912
rect 11992 18884 12020 18924
rect 12434 18884 12440 18896
rect 7392 18856 12020 18884
rect 12084 18856 12440 18884
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18816 1823 18819
rect 2222 18816 2228 18828
rect 1811 18788 2228 18816
rect 1811 18785 1823 18788
rect 1765 18779 1823 18785
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 2314 18776 2320 18828
rect 2372 18816 2378 18828
rect 2961 18819 3019 18825
rect 2372 18788 2417 18816
rect 2372 18776 2378 18788
rect 2961 18785 2973 18819
rect 3007 18816 3019 18819
rect 6273 18819 6331 18825
rect 3007 18788 3648 18816
rect 3007 18785 3019 18788
rect 2961 18779 3019 18785
rect 3620 18760 3648 18788
rect 6273 18785 6285 18819
rect 6319 18816 6331 18819
rect 7006 18816 7012 18828
rect 6319 18788 7012 18816
rect 6319 18785 6331 18788
rect 6273 18779 6331 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 7156 18788 9505 18816
rect 7156 18776 7162 18788
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 10318 18816 10324 18828
rect 10279 18788 10324 18816
rect 9493 18779 9551 18785
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 12084 18825 12112 18856
rect 12434 18844 12440 18856
rect 12492 18884 12498 18896
rect 13170 18884 13176 18896
rect 12492 18856 13176 18884
rect 12492 18844 12498 18856
rect 13170 18844 13176 18856
rect 13228 18844 13234 18896
rect 13280 18884 13308 18924
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 15102 18912 15108 18964
rect 15160 18952 15166 18964
rect 15473 18955 15531 18961
rect 15473 18952 15485 18955
rect 15160 18924 15485 18952
rect 15160 18912 15166 18924
rect 15473 18921 15485 18924
rect 15519 18921 15531 18955
rect 15473 18915 15531 18921
rect 15654 18912 15660 18964
rect 15712 18952 15718 18964
rect 20438 18952 20444 18964
rect 15712 18924 20208 18952
rect 20399 18924 20444 18952
rect 15712 18912 15718 18924
rect 13280 18856 15516 18884
rect 11517 18819 11575 18825
rect 11517 18785 11529 18819
rect 11563 18816 11575 18819
rect 12069 18819 12127 18825
rect 11563 18788 12020 18816
rect 11563 18785 11575 18788
rect 11517 18779 11575 18785
rect 3418 18748 3424 18760
rect 2976 18720 3424 18748
rect 1118 18640 1124 18692
rect 1176 18680 1182 18692
rect 2976 18680 3004 18720
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 3602 18708 3608 18760
rect 3660 18708 3666 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18717 4859 18751
rect 6362 18748 6368 18760
rect 6323 18720 6368 18748
rect 4801 18711 4859 18717
rect 1176 18652 3004 18680
rect 1176 18640 1182 18652
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 4816 18612 4844 18711
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 6512 18720 6557 18748
rect 6512 18708 6518 18720
rect 7282 18708 7288 18760
rect 7340 18748 7346 18760
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 7340 18720 8401 18748
rect 7340 18708 7346 18720
rect 8389 18717 8401 18720
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18748 8631 18751
rect 9122 18748 9128 18760
rect 8619 18720 9128 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 9732 18720 10425 18748
rect 9732 18708 9738 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10594 18748 10600 18760
rect 10555 18720 10600 18748
rect 10413 18711 10471 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11606 18748 11612 18760
rect 11103 18720 11612 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 5813 18683 5871 18689
rect 5813 18649 5825 18683
rect 5859 18680 5871 18683
rect 9950 18680 9956 18692
rect 5859 18652 9812 18680
rect 9911 18652 9956 18680
rect 5859 18649 5871 18652
rect 5813 18643 5871 18649
rect 4764 18584 4844 18612
rect 4764 18572 4770 18584
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 5442 18612 5448 18624
rect 4948 18584 5448 18612
rect 4948 18572 4954 18584
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 5902 18612 5908 18624
rect 5863 18584 5908 18612
rect 5902 18572 5908 18584
rect 5960 18572 5966 18624
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 9030 18612 9036 18624
rect 7975 18584 9036 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9784 18612 9812 18652
rect 9950 18640 9956 18652
rect 10008 18640 10014 18692
rect 11698 18680 11704 18692
rect 11659 18652 11704 18680
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 11992 18680 12020 18788
rect 12069 18785 12081 18819
rect 12115 18785 12127 18819
rect 12069 18779 12127 18785
rect 12336 18819 12394 18825
rect 12336 18785 12348 18819
rect 12382 18816 12394 18819
rect 13354 18816 13360 18828
rect 12382 18788 13360 18816
rect 12382 18785 12394 18788
rect 12336 18779 12394 18785
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13725 18819 13783 18825
rect 13725 18785 13737 18819
rect 13771 18816 13783 18819
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 13771 18788 14565 18816
rect 13771 18785 13783 18788
rect 13725 18779 13783 18785
rect 14553 18785 14565 18788
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 15289 18819 15347 18825
rect 15289 18785 15301 18819
rect 15335 18816 15347 18819
rect 15378 18816 15384 18828
rect 15335 18788 15384 18816
rect 15335 18785 15347 18788
rect 15289 18779 15347 18785
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 15488 18816 15516 18856
rect 15746 18844 15752 18896
rect 15804 18884 15810 18896
rect 16178 18887 16236 18893
rect 16178 18884 16190 18887
rect 15804 18856 16190 18884
rect 15804 18844 15810 18856
rect 16178 18853 16190 18856
rect 16224 18853 16236 18887
rect 20070 18884 20076 18896
rect 16178 18847 16236 18853
rect 16296 18856 20076 18884
rect 16296 18816 16324 18856
rect 20070 18844 20076 18856
rect 20128 18844 20134 18896
rect 20180 18884 20208 18924
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 22462 18884 22468 18896
rect 20180 18856 22468 18884
rect 22462 18844 22468 18856
rect 22520 18844 22526 18896
rect 15488 18788 16324 18816
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 17862 18825 17868 18828
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 16632 18788 17601 18816
rect 16632 18776 16638 18788
rect 17589 18785 17601 18788
rect 17635 18785 17647 18819
rect 17856 18816 17868 18825
rect 17589 18779 17647 18785
rect 17696 18788 17868 18816
rect 13372 18748 13400 18776
rect 13998 18748 14004 18760
rect 13372 18720 14004 18748
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 14642 18748 14648 18760
rect 14603 18720 14648 18748
rect 14642 18708 14648 18720
rect 14700 18708 14706 18760
rect 14826 18748 14832 18760
rect 14787 18720 14832 18748
rect 14826 18708 14832 18720
rect 14884 18708 14890 18760
rect 15930 18748 15936 18760
rect 15891 18720 15936 18748
rect 15930 18708 15936 18720
rect 15988 18708 15994 18760
rect 17696 18748 17724 18788
rect 17856 18779 17868 18788
rect 17862 18776 17868 18779
rect 17920 18776 17926 18828
rect 18782 18776 18788 18828
rect 18840 18816 18846 18828
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 18840 18788 19073 18816
rect 18840 18776 18846 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19242 18816 19248 18828
rect 19203 18788 19248 18816
rect 19061 18779 19119 18785
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19352 18788 19656 18816
rect 19352 18748 19380 18788
rect 19518 18748 19524 18760
rect 17328 18720 17724 18748
rect 18616 18720 19380 18748
rect 19479 18720 19524 18748
rect 12066 18680 12072 18692
rect 11992 18652 12072 18680
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 14185 18683 14243 18689
rect 14185 18649 14197 18683
rect 14231 18680 14243 18683
rect 15286 18680 15292 18692
rect 14231 18652 15292 18680
rect 14231 18649 14243 18652
rect 14185 18643 14243 18649
rect 15286 18640 15292 18652
rect 15344 18640 15350 18692
rect 17328 18689 17356 18720
rect 17313 18683 17371 18689
rect 17313 18649 17325 18683
rect 17359 18649 17371 18683
rect 17313 18643 17371 18649
rect 15838 18612 15844 18624
rect 9784 18584 15844 18612
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 15930 18572 15936 18624
rect 15988 18612 15994 18624
rect 16574 18612 16580 18624
rect 15988 18584 16580 18612
rect 15988 18572 15994 18584
rect 16574 18572 16580 18584
rect 16632 18572 16638 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 18616 18612 18644 18720
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 19628 18748 19656 18788
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 20036 18788 20269 18816
rect 20036 18776 20042 18788
rect 20257 18785 20269 18788
rect 20303 18785 20315 18819
rect 21542 18816 21548 18828
rect 20257 18779 20315 18785
rect 20364 18788 21548 18816
rect 20364 18748 20392 18788
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 19628 18720 20392 18748
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 18969 18683 19027 18689
rect 18969 18680 18981 18683
rect 18932 18652 18981 18680
rect 18932 18640 18938 18652
rect 18969 18649 18981 18652
rect 19015 18649 19027 18683
rect 18969 18643 19027 18649
rect 19061 18683 19119 18689
rect 19061 18649 19073 18683
rect 19107 18680 19119 18683
rect 20916 18680 20944 18711
rect 19107 18652 20944 18680
rect 19107 18649 19119 18652
rect 19061 18643 19119 18649
rect 16724 18584 18644 18612
rect 16724 18572 16730 18584
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1762 18408 1768 18420
rect 1723 18380 1768 18408
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 2314 18368 2320 18420
rect 2372 18408 2378 18420
rect 3050 18408 3056 18420
rect 2372 18380 2912 18408
rect 3011 18380 3056 18408
rect 2372 18368 2378 18380
rect 2884 18340 2912 18380
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 6178 18408 6184 18420
rect 4264 18380 6184 18408
rect 4154 18340 4160 18352
rect 2884 18312 4160 18340
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 4264 18272 4292 18380
rect 6178 18368 6184 18380
rect 6236 18368 6242 18420
rect 6362 18368 6368 18420
rect 6420 18408 6426 18420
rect 6825 18411 6883 18417
rect 6825 18408 6837 18411
rect 6420 18380 6837 18408
rect 6420 18368 6426 18380
rect 6825 18377 6837 18380
rect 6871 18377 6883 18411
rect 8294 18408 8300 18420
rect 6825 18371 6883 18377
rect 7944 18380 8300 18408
rect 5626 18340 5632 18352
rect 5539 18312 5632 18340
rect 5626 18300 5632 18312
rect 5684 18340 5690 18352
rect 6454 18340 6460 18352
rect 5684 18312 6460 18340
rect 5684 18300 5690 18312
rect 6454 18300 6460 18312
rect 6512 18300 6518 18352
rect 2148 18244 4292 18272
rect 1578 18204 1584 18216
rect 1539 18176 1584 18204
rect 1578 18164 1584 18176
rect 1636 18164 1642 18216
rect 2148 18213 2176 18244
rect 5350 18232 5356 18284
rect 5408 18272 5414 18284
rect 7282 18272 7288 18284
rect 5408 18244 7288 18272
rect 5408 18232 5414 18244
rect 7282 18232 7288 18244
rect 7340 18272 7346 18284
rect 7469 18275 7527 18281
rect 7340 18244 7433 18272
rect 7340 18232 7346 18244
rect 7469 18241 7481 18275
rect 7515 18272 7527 18275
rect 7558 18272 7564 18284
rect 7515 18244 7564 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2409 18207 2467 18213
rect 2409 18204 2421 18207
rect 2280 18176 2421 18204
rect 2280 18164 2286 18176
rect 2409 18173 2421 18176
rect 2455 18173 2467 18207
rect 2409 18167 2467 18173
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18173 2927 18207
rect 2869 18167 2927 18173
rect 2884 18136 2912 18167
rect 2958 18164 2964 18216
rect 3016 18204 3022 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3016 18176 3433 18204
rect 3016 18164 3022 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 4212 18176 4261 18204
rect 4212 18164 4218 18176
rect 4249 18173 4261 18176
rect 4295 18204 4307 18207
rect 4295 18176 5396 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 5368 18148 5396 18176
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 7098 18204 7104 18216
rect 5500 18176 7104 18204
rect 5500 18164 5506 18176
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 7193 18207 7251 18213
rect 7193 18173 7205 18207
rect 7239 18204 7251 18207
rect 7944 18204 7972 18380
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 10042 18408 10048 18420
rect 8444 18380 9260 18408
rect 8444 18368 8450 18380
rect 9232 18272 9260 18380
rect 9692 18380 10048 18408
rect 9692 18281 9720 18380
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 10594 18368 10600 18420
rect 10652 18408 10658 18420
rect 11057 18411 11115 18417
rect 11057 18408 11069 18411
rect 10652 18380 11069 18408
rect 10652 18368 10658 18380
rect 11057 18377 11069 18380
rect 11103 18377 11115 18411
rect 12526 18408 12532 18420
rect 12487 18380 12532 18408
rect 11057 18371 11115 18377
rect 12526 18368 12532 18380
rect 12584 18368 12590 18420
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 13228 18380 14228 18408
rect 13228 18368 13234 18380
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 13449 18343 13507 18349
rect 13449 18340 13461 18343
rect 11664 18312 13461 18340
rect 11664 18300 11670 18312
rect 13449 18309 13461 18312
rect 13495 18309 13507 18343
rect 13449 18303 13507 18309
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9232 18244 9689 18272
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 11977 18275 12035 18281
rect 11977 18241 11989 18275
rect 12023 18272 12035 18275
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 12023 18244 12173 18272
rect 12023 18241 12035 18244
rect 11977 18235 12035 18241
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12768 18244 13001 18272
rect 12768 18232 12774 18244
rect 12989 18241 13001 18244
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13354 18272 13360 18284
rect 13219 18244 13360 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 13998 18232 14004 18284
rect 14056 18272 14062 18284
rect 14093 18275 14151 18281
rect 14093 18272 14105 18275
rect 14056 18244 14105 18272
rect 14056 18232 14062 18244
rect 14093 18241 14105 18244
rect 14139 18241 14151 18275
rect 14200 18272 14228 18380
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 15562 18408 15568 18420
rect 15344 18380 15568 18408
rect 15344 18368 15350 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 15933 18411 15991 18417
rect 15933 18408 15945 18411
rect 15804 18380 15945 18408
rect 15804 18368 15810 18380
rect 15933 18377 15945 18380
rect 15979 18377 15991 18411
rect 15933 18371 15991 18377
rect 16298 18368 16304 18420
rect 16356 18408 16362 18420
rect 16485 18411 16543 18417
rect 16485 18408 16497 18411
rect 16356 18380 16497 18408
rect 16356 18368 16362 18380
rect 16485 18377 16497 18380
rect 16531 18377 16543 18411
rect 16485 18371 16543 18377
rect 17037 18411 17095 18417
rect 17037 18377 17049 18411
rect 17083 18408 17095 18411
rect 17494 18408 17500 18420
rect 17083 18380 17500 18408
rect 17083 18377 17095 18380
rect 17037 18371 17095 18377
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 17770 18408 17776 18420
rect 17635 18380 17776 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 18012 18380 18061 18408
rect 18012 18368 18018 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18874 18408 18880 18420
rect 18049 18371 18107 18377
rect 18156 18380 18880 18408
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 16666 18340 16672 18352
rect 15896 18312 16672 18340
rect 15896 18300 15902 18312
rect 16666 18300 16672 18312
rect 16724 18300 16730 18352
rect 18156 18340 18184 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 19150 18368 19156 18420
rect 19208 18408 19214 18420
rect 19613 18411 19671 18417
rect 19613 18408 19625 18411
rect 19208 18380 19625 18408
rect 19208 18368 19214 18380
rect 19613 18377 19625 18380
rect 19659 18377 19671 18411
rect 19613 18371 19671 18377
rect 16776 18312 18184 18340
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14200 18244 14565 18272
rect 14093 18235 14151 18241
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 16776 18272 16804 18312
rect 18230 18300 18236 18352
rect 18288 18340 18294 18352
rect 20898 18340 20904 18352
rect 18288 18312 20024 18340
rect 20859 18312 20904 18340
rect 18288 18300 18294 18312
rect 14553 18235 14611 18241
rect 15580 18244 16804 18272
rect 7239 18176 7972 18204
rect 8021 18207 8079 18213
rect 7239 18173 7251 18176
rect 7193 18167 7251 18173
rect 8021 18173 8033 18207
rect 8067 18204 8079 18207
rect 8110 18204 8116 18216
rect 8067 18176 8116 18204
rect 8067 18173 8079 18176
rect 8021 18167 8079 18173
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 15580 18204 15608 18244
rect 17862 18232 17868 18284
rect 17920 18272 17926 18284
rect 18693 18275 18751 18281
rect 18693 18272 18705 18275
rect 17920 18244 18705 18272
rect 17920 18232 17926 18244
rect 18693 18241 18705 18244
rect 18739 18241 18751 18275
rect 18693 18235 18751 18241
rect 18874 18232 18880 18284
rect 18932 18272 18938 18284
rect 19794 18272 19800 18284
rect 18932 18244 19800 18272
rect 18932 18232 18938 18244
rect 19794 18232 19800 18244
rect 19852 18232 19858 18284
rect 8220 18176 15608 18204
rect 16301 18207 16359 18213
rect 3786 18136 3792 18148
rect 2884 18108 3792 18136
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 4516 18139 4574 18145
rect 4516 18105 4528 18139
rect 4562 18136 4574 18139
rect 4982 18136 4988 18148
rect 4562 18108 4988 18136
rect 4562 18105 4574 18108
rect 4516 18099 4574 18105
rect 4982 18096 4988 18108
rect 5040 18096 5046 18148
rect 5350 18096 5356 18148
rect 5408 18096 5414 18148
rect 8220 18136 8248 18176
rect 16301 18173 16313 18207
rect 16347 18204 16359 18207
rect 16574 18204 16580 18216
rect 16347 18176 16580 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 16850 18204 16856 18216
rect 16811 18176 16856 18204
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 16942 18164 16948 18216
rect 17000 18204 17006 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 17000 18176 17417 18204
rect 17000 18164 17006 18176
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 18417 18207 18475 18213
rect 18417 18173 18429 18207
rect 18463 18204 18475 18207
rect 18782 18204 18788 18216
rect 18463 18176 18788 18204
rect 18463 18173 18475 18176
rect 18417 18167 18475 18173
rect 18782 18164 18788 18176
rect 18840 18164 18846 18216
rect 19426 18204 19432 18216
rect 19387 18176 19432 18204
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 19996 18213 20024 18312
rect 20898 18300 20904 18312
rect 20956 18300 20962 18352
rect 19981 18207 20039 18213
rect 19981 18173 19993 18207
rect 20027 18173 20039 18207
rect 20714 18204 20720 18216
rect 20675 18176 20720 18204
rect 19981 18167 20039 18173
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 7668 18108 8248 18136
rect 8288 18139 8346 18145
rect 658 18028 664 18080
rect 716 18068 722 18080
rect 2590 18068 2596 18080
rect 716 18040 2596 18068
rect 716 18028 722 18040
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 7668 18068 7696 18108
rect 8288 18105 8300 18139
rect 8334 18136 8346 18139
rect 9122 18136 9128 18148
rect 8334 18108 9128 18136
rect 8334 18105 8346 18108
rect 8288 18099 8346 18105
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 9766 18136 9772 18148
rect 9416 18108 9772 18136
rect 3651 18040 7696 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 8386 18068 8392 18080
rect 7800 18040 8392 18068
rect 7800 18028 7806 18040
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 9416 18077 9444 18108
rect 9766 18096 9772 18108
rect 9824 18136 9830 18148
rect 9944 18139 10002 18145
rect 9944 18136 9956 18139
rect 9824 18108 9956 18136
rect 9824 18096 9830 18108
rect 9944 18105 9956 18108
rect 9990 18136 10002 18139
rect 10870 18136 10876 18148
rect 9990 18108 10876 18136
rect 9990 18105 10002 18108
rect 9944 18099 10002 18105
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 11606 18096 11612 18148
rect 11664 18136 11670 18148
rect 14826 18145 14832 18148
rect 11793 18139 11851 18145
rect 11793 18136 11805 18139
rect 11664 18108 11805 18136
rect 11664 18096 11670 18108
rect 11793 18105 11805 18108
rect 11839 18105 11851 18139
rect 11793 18099 11851 18105
rect 12897 18139 12955 18145
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 13449 18139 13507 18145
rect 12943 18108 13400 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18037 9459 18071
rect 9401 18031 9459 18037
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11333 18071 11391 18077
rect 11333 18068 11345 18071
rect 11112 18040 11345 18068
rect 11112 18028 11118 18040
rect 11333 18037 11345 18040
rect 11379 18037 11391 18071
rect 11698 18068 11704 18080
rect 11659 18040 11704 18068
rect 11333 18031 11391 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12158 18068 12164 18080
rect 12071 18040 12164 18068
rect 12158 18028 12164 18040
rect 12216 18068 12222 18080
rect 13078 18068 13084 18080
rect 12216 18040 13084 18068
rect 12216 18028 12222 18040
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13372 18068 13400 18108
rect 13449 18105 13461 18139
rect 13495 18136 13507 18139
rect 13909 18139 13967 18145
rect 13909 18136 13921 18139
rect 13495 18108 13921 18136
rect 13495 18105 13507 18108
rect 13449 18099 13507 18105
rect 13909 18105 13921 18108
rect 13955 18105 13967 18139
rect 14820 18136 14832 18145
rect 14739 18108 14832 18136
rect 13909 18099 13967 18105
rect 14820 18099 14832 18108
rect 14884 18136 14890 18148
rect 15838 18136 15844 18148
rect 14884 18108 15844 18136
rect 14826 18096 14832 18099
rect 14884 18096 14890 18108
rect 15838 18096 15844 18108
rect 15896 18096 15902 18148
rect 18046 18096 18052 18148
rect 18104 18136 18110 18148
rect 20257 18139 20315 18145
rect 20257 18136 20269 18139
rect 18104 18108 20269 18136
rect 18104 18096 18110 18108
rect 20257 18105 20269 18108
rect 20303 18105 20315 18139
rect 20257 18099 20315 18105
rect 13541 18071 13599 18077
rect 13541 18068 13553 18071
rect 13372 18040 13553 18068
rect 13541 18037 13553 18040
rect 13587 18037 13599 18071
rect 13541 18031 13599 18037
rect 14001 18071 14059 18077
rect 14001 18037 14013 18071
rect 14047 18068 14059 18071
rect 14182 18068 14188 18080
rect 14047 18040 14188 18068
rect 14047 18037 14059 18040
rect 14001 18031 14059 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 15194 18028 15200 18080
rect 15252 18068 15258 18080
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 15252 18040 18521 18068
rect 15252 18028 15258 18040
rect 18509 18037 18521 18040
rect 18555 18068 18567 18071
rect 18598 18068 18604 18080
rect 18555 18040 18604 18068
rect 18555 18037 18567 18040
rect 18509 18031 18567 18037
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 18782 18028 18788 18080
rect 18840 18068 18846 18080
rect 19702 18068 19708 18080
rect 18840 18040 19708 18068
rect 18840 18028 18846 18040
rect 19702 18028 19708 18040
rect 19760 18028 19766 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 3050 17864 3056 17876
rect 3011 17836 3056 17864
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 4246 17824 4252 17876
rect 4304 17864 4310 17876
rect 5074 17864 5080 17876
rect 4304 17836 5080 17864
rect 4304 17824 4310 17836
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 7006 17864 7012 17876
rect 6967 17836 7012 17864
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 7469 17867 7527 17873
rect 7469 17833 7481 17867
rect 7515 17864 7527 17867
rect 10410 17864 10416 17876
rect 7515 17836 10416 17864
rect 7515 17833 7527 17836
rect 7469 17827 7527 17833
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 11885 17867 11943 17873
rect 11885 17864 11897 17867
rect 11756 17836 11897 17864
rect 11756 17824 11762 17836
rect 11885 17833 11897 17836
rect 11931 17833 11943 17867
rect 13722 17864 13728 17876
rect 11885 17827 11943 17833
rect 11992 17836 13728 17864
rect 2682 17756 2688 17808
rect 2740 17796 2746 17808
rect 9950 17796 9956 17808
rect 2740 17768 9956 17796
rect 2740 17756 2746 17768
rect 9950 17756 9956 17768
rect 10008 17756 10014 17808
rect 10502 17805 10508 17808
rect 10496 17759 10508 17805
rect 10560 17796 10566 17808
rect 10560 17768 10596 17796
rect 10502 17756 10508 17759
rect 10560 17756 10566 17768
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17697 1639 17731
rect 2130 17728 2136 17740
rect 2188 17737 2194 17740
rect 2188 17731 2201 17737
rect 2101 17700 2136 17728
rect 1581 17691 1639 17697
rect 1596 17660 1624 17691
rect 2130 17688 2136 17700
rect 2189 17697 2201 17731
rect 2188 17691 2201 17697
rect 2869 17731 2927 17737
rect 2869 17697 2881 17731
rect 2915 17697 2927 17731
rect 2869 17691 2927 17697
rect 2188 17688 2194 17691
rect 2317 17663 2375 17669
rect 2317 17660 2329 17663
rect 1596 17632 2329 17660
rect 2317 17629 2329 17632
rect 2363 17629 2375 17663
rect 2884 17660 2912 17691
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 5626 17737 5632 17740
rect 4709 17731 4767 17737
rect 4709 17728 4721 17731
rect 4304 17700 4721 17728
rect 4304 17688 4310 17700
rect 4709 17697 4721 17700
rect 4755 17697 4767 17731
rect 5620 17728 5632 17737
rect 4709 17691 4767 17697
rect 5000 17700 5632 17728
rect 4614 17660 4620 17672
rect 2884 17632 4620 17660
rect 2317 17623 2375 17629
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 5000 17669 5028 17700
rect 5620 17691 5632 17700
rect 5626 17688 5632 17691
rect 5684 17688 5690 17740
rect 7006 17688 7012 17740
rect 7064 17728 7070 17740
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 7064 17700 7389 17728
rect 7064 17688 7070 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 8941 17731 8999 17737
rect 8941 17697 8953 17731
rect 8987 17728 8999 17731
rect 9306 17728 9312 17740
rect 8987 17700 9312 17728
rect 8987 17697 8999 17700
rect 8941 17691 8999 17697
rect 9306 17688 9312 17700
rect 9364 17688 9370 17740
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9456 17700 9996 17728
rect 9456 17688 9462 17700
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17629 5043 17663
rect 5350 17660 5356 17672
rect 5311 17632 5356 17660
rect 4985 17623 5043 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 7558 17660 7564 17672
rect 7519 17632 7564 17660
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 9030 17660 9036 17672
rect 8991 17632 9036 17660
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17660 9275 17663
rect 9766 17660 9772 17672
rect 9263 17632 9772 17660
rect 9263 17629 9275 17632
rect 9217 17623 9275 17629
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 9968 17660 9996 17700
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 10229 17731 10287 17737
rect 10229 17728 10241 17731
rect 10100 17700 10241 17728
rect 10100 17688 10106 17700
rect 10229 17697 10241 17700
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 10336 17700 11560 17728
rect 10336 17660 10364 17700
rect 9968 17632 10364 17660
rect 11532 17660 11560 17700
rect 11992 17660 12020 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 13817 17867 13875 17873
rect 13817 17833 13829 17867
rect 13863 17864 13875 17867
rect 13998 17864 14004 17876
rect 13863 17836 14004 17864
rect 13863 17833 13875 17836
rect 13817 17827 13875 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 14274 17864 14280 17876
rect 14231 17836 14280 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 14458 17824 14464 17876
rect 14516 17864 14522 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14516 17836 14657 17864
rect 14516 17824 14522 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 14645 17827 14703 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15396 17836 15792 17864
rect 15102 17756 15108 17808
rect 15160 17796 15166 17808
rect 15396 17796 15424 17836
rect 15160 17768 15424 17796
rect 15160 17756 15166 17768
rect 12437 17731 12495 17737
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 12526 17728 12532 17740
rect 12483 17700 12532 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 12704 17731 12762 17737
rect 12704 17697 12716 17731
rect 12750 17728 12762 17731
rect 14366 17728 14372 17740
rect 12750 17700 14372 17728
rect 12750 17697 12762 17700
rect 12704 17691 12762 17697
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 14550 17728 14556 17740
rect 14511 17700 14556 17728
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 15764 17737 15792 17836
rect 16206 17824 16212 17876
rect 16264 17864 16270 17876
rect 20438 17864 20444 17876
rect 16264 17836 20444 17864
rect 16264 17824 16270 17836
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 16574 17796 16580 17808
rect 16535 17768 16580 17796
rect 16574 17756 16580 17768
rect 16632 17756 16638 17808
rect 18224 17799 18282 17805
rect 18224 17765 18236 17799
rect 18270 17796 18282 17799
rect 18966 17796 18972 17808
rect 18270 17768 18972 17796
rect 18270 17765 18282 17768
rect 18224 17759 18282 17765
rect 18966 17756 18972 17768
rect 19024 17756 19030 17808
rect 19426 17756 19432 17808
rect 19484 17796 19490 17808
rect 20257 17799 20315 17805
rect 20257 17796 20269 17799
rect 19484 17768 20269 17796
rect 19484 17756 19490 17768
rect 20257 17765 20269 17768
rect 20303 17765 20315 17799
rect 20257 17759 20315 17765
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17728 15807 17731
rect 16022 17728 16028 17740
rect 15795 17700 16028 17728
rect 15795 17697 15807 17700
rect 15749 17691 15807 17697
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 16298 17728 16304 17740
rect 16259 17700 16304 17728
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 17405 17731 17463 17737
rect 17405 17697 17417 17731
rect 17451 17728 17463 17731
rect 18046 17728 18052 17740
rect 17451 17700 18052 17728
rect 17451 17697 17463 17700
rect 17405 17691 17463 17697
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 19978 17728 19984 17740
rect 19939 17700 19984 17728
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 11532 17632 12020 17660
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15010 17660 15016 17672
rect 14875 17632 15016 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 15930 17620 15936 17672
rect 15988 17660 15994 17672
rect 17954 17660 17960 17672
rect 15988 17632 17960 17660
rect 15988 17620 15994 17632
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 8573 17595 8631 17601
rect 8573 17561 8585 17595
rect 8619 17592 8631 17595
rect 9674 17592 9680 17604
rect 8619 17564 9680 17592
rect 8619 17561 8631 17564
rect 8573 17555 8631 17561
rect 9674 17552 9680 17564
rect 9732 17552 9738 17604
rect 12158 17592 12164 17604
rect 11155 17564 12164 17592
rect 1762 17524 1768 17536
rect 1723 17496 1768 17524
rect 1762 17484 1768 17496
rect 1820 17484 1826 17536
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 4154 17524 4160 17536
rect 2556 17496 4160 17524
rect 2556 17484 2562 17496
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 5994 17524 6000 17536
rect 4387 17496 6000 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 5994 17484 6000 17496
rect 6052 17484 6058 17536
rect 6730 17524 6736 17536
rect 6691 17496 6736 17524
rect 6730 17484 6736 17496
rect 6788 17484 6794 17536
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 8846 17524 8852 17536
rect 6880 17496 8852 17524
rect 6880 17484 6886 17496
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 9122 17484 9128 17536
rect 9180 17524 9186 17536
rect 9950 17524 9956 17536
rect 9180 17496 9956 17524
rect 9180 17484 9186 17496
rect 9950 17484 9956 17496
rect 10008 17524 10014 17536
rect 11155 17524 11183 17564
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 13630 17552 13636 17604
rect 13688 17592 13694 17604
rect 17218 17592 17224 17604
rect 13688 17564 17224 17592
rect 13688 17552 13694 17564
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 11606 17524 11612 17536
rect 10008 17496 11183 17524
rect 11567 17496 11612 17524
rect 10008 17484 10014 17496
rect 11606 17484 11612 17496
rect 11664 17484 11670 17536
rect 13722 17484 13728 17536
rect 13780 17524 13786 17536
rect 16574 17524 16580 17536
rect 13780 17496 16580 17524
rect 13780 17484 13786 17496
rect 16574 17484 16580 17496
rect 16632 17524 16638 17536
rect 17494 17524 17500 17536
rect 16632 17496 17500 17524
rect 16632 17484 16638 17496
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 17589 17527 17647 17533
rect 17589 17493 17601 17527
rect 17635 17524 17647 17527
rect 18598 17524 18604 17536
rect 17635 17496 18604 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 19334 17524 19340 17536
rect 19295 17496 19340 17524
rect 19334 17484 19340 17496
rect 19392 17484 19398 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 4617 17323 4675 17329
rect 2884 17292 4476 17320
rect 2884 17252 2912 17292
rect 2056 17224 2912 17252
rect 4341 17255 4399 17261
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 2056 17116 2084 17224
rect 4341 17221 4353 17255
rect 4387 17221 4399 17255
rect 4448 17252 4476 17292
rect 4617 17289 4629 17323
rect 4663 17320 4675 17323
rect 4798 17320 4804 17332
rect 4663 17292 4804 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5592 17292 5641 17320
rect 5592 17280 5598 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 7558 17320 7564 17332
rect 5629 17283 5687 17289
rect 5736 17292 7564 17320
rect 5442 17252 5448 17264
rect 4448 17224 5448 17252
rect 4341 17215 4399 17221
rect 2498 17144 2504 17196
rect 2556 17184 2562 17196
rect 2961 17187 3019 17193
rect 2961 17184 2973 17187
rect 2556 17156 2973 17184
rect 2556 17144 2562 17156
rect 2961 17153 2973 17156
rect 3007 17153 3019 17187
rect 4356 17184 4384 17215
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 4982 17184 4988 17196
rect 4356 17156 4988 17184
rect 2961 17147 3019 17153
rect 4982 17144 4988 17156
rect 5040 17184 5046 17196
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 5040 17156 5273 17184
rect 5040 17144 5046 17156
rect 5261 17153 5273 17156
rect 5307 17184 5319 17187
rect 5736 17184 5764 17292
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 9306 17320 9312 17332
rect 9267 17292 9312 17320
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 10318 17320 10324 17332
rect 10279 17292 10324 17320
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 19978 17320 19984 17332
rect 10560 17292 19984 17320
rect 10560 17280 10566 17292
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 6822 17252 6828 17264
rect 5307 17156 5764 17184
rect 5828 17224 6828 17252
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 1811 17088 2084 17116
rect 2317 17119 2375 17125
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2317 17085 2329 17119
rect 2363 17116 2375 17119
rect 4890 17116 4896 17128
rect 2363 17088 4896 17116
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 5074 17116 5080 17128
rect 4987 17088 5080 17116
rect 5074 17076 5080 17088
rect 5132 17116 5138 17128
rect 5828 17116 5856 17224
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 8202 17212 8208 17264
rect 8260 17252 8266 17264
rect 12342 17252 12348 17264
rect 8260 17224 12348 17252
rect 8260 17212 8266 17224
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 12437 17255 12495 17261
rect 12437 17221 12449 17255
rect 12483 17252 12495 17255
rect 13630 17252 13636 17264
rect 12483 17224 12572 17252
rect 13591 17224 13636 17252
rect 12483 17221 12495 17224
rect 12437 17215 12495 17221
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 5960 17156 6101 17184
rect 5960 17144 5966 17156
rect 6089 17153 6101 17156
rect 6135 17153 6147 17187
rect 6089 17147 6147 17153
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17184 6331 17187
rect 6730 17184 6736 17196
rect 6319 17156 6736 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 6730 17144 6736 17156
rect 6788 17184 6794 17196
rect 9950 17184 9956 17196
rect 6788 17156 6960 17184
rect 9911 17156 9956 17184
rect 6788 17144 6794 17156
rect 5994 17116 6000 17128
rect 5132 17088 5856 17116
rect 5955 17088 6000 17116
rect 5132 17076 5138 17088
rect 5994 17076 6000 17088
rect 6052 17076 6058 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6932 17116 6960 17156
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10870 17184 10876 17196
rect 10831 17156 10876 17184
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 11974 17184 11980 17196
rect 11935 17156 11980 17184
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 7081 17119 7139 17125
rect 7081 17116 7093 17119
rect 6932 17088 7093 17116
rect 6825 17079 6883 17085
rect 7081 17085 7093 17088
rect 7127 17085 7139 17119
rect 7081 17079 7139 17085
rect 9769 17119 9827 17125
rect 9769 17085 9781 17119
rect 9815 17116 9827 17119
rect 10594 17116 10600 17128
rect 9815 17088 10600 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 3206 17051 3264 17057
rect 3206 17048 3218 17051
rect 3016 17020 3218 17048
rect 3016 17008 3022 17020
rect 3206 17017 3218 17020
rect 3252 17017 3264 17051
rect 3206 17011 3264 17017
rect 3510 17008 3516 17060
rect 3568 17048 3574 17060
rect 3568 17020 5304 17048
rect 3568 17008 3574 17020
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 2590 16940 2596 16992
rect 2648 16980 2654 16992
rect 4154 16980 4160 16992
rect 2648 16952 4160 16980
rect 2648 16940 2654 16952
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 4856 16952 4997 16980
rect 4856 16940 4862 16952
rect 4985 16949 4997 16952
rect 5031 16949 5043 16983
rect 5276 16980 5304 17020
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 6840 17048 6868 17079
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 11054 17116 11060 17128
rect 10735 17088 11060 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17116 11759 17119
rect 12434 17116 12440 17128
rect 11747 17088 12440 17116
rect 11747 17085 11759 17088
rect 11701 17079 11759 17085
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 9398 17048 9404 17060
rect 5408 17020 6868 17048
rect 7668 17020 9404 17048
rect 5408 17008 5414 17020
rect 7668 16980 7696 17020
rect 9398 17008 9404 17020
rect 9456 17008 9462 17060
rect 9677 17051 9735 17057
rect 9677 17017 9689 17051
rect 9723 17048 9735 17051
rect 10781 17051 10839 17057
rect 9723 17020 10640 17048
rect 9723 17017 9735 17020
rect 9677 17011 9735 17017
rect 5276 16952 7696 16980
rect 4985 16943 5043 16949
rect 7742 16940 7748 16992
rect 7800 16980 7806 16992
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 7800 16952 8217 16980
rect 7800 16940 7806 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 10612 16980 10640 17020
rect 10781 17017 10793 17051
rect 10827 17048 10839 17051
rect 12544 17048 12572 17224
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 14366 17212 14372 17264
rect 14424 17252 14430 17264
rect 19610 17252 19616 17264
rect 14424 17224 14596 17252
rect 19571 17224 19616 17252
rect 14424 17212 14430 17224
rect 13078 17184 13084 17196
rect 13039 17156 13084 17184
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 14568 17193 14596 17224
rect 19610 17212 19616 17224
rect 19668 17212 19674 17264
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14332 17156 14473 17184
rect 14332 17144 14338 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 15212 17156 15976 17184
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13320 17088 13461 17116
rect 13320 17076 13326 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 13449 17079 13507 17085
rect 14016 17088 15025 17116
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 10827 17020 12572 17048
rect 12728 17020 12817 17048
rect 10827 17017 10839 17020
rect 10781 17011 10839 17017
rect 10686 16980 10692 16992
rect 10612 16952 10692 16980
rect 8205 16943 8263 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11333 16983 11391 16989
rect 11333 16980 11345 16983
rect 11020 16952 11345 16980
rect 11020 16940 11026 16952
rect 11333 16949 11345 16952
rect 11379 16949 11391 16983
rect 11333 16943 11391 16949
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11480 16952 11805 16980
rect 11480 16940 11486 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11793 16943 11851 16949
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 12728 16980 12756 17020
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 12805 17011 12863 17017
rect 12894 16980 12900 16992
rect 12400 16952 12756 16980
rect 12855 16952 12900 16980
rect 12400 16940 12406 16952
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 14016 16989 14044 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 14274 17008 14280 17060
rect 14332 17048 14338 17060
rect 15212 17048 15240 17156
rect 15838 17116 15844 17128
rect 15799 17088 15844 17116
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 15948 17116 15976 17156
rect 17954 17144 17960 17196
rect 18012 17184 18018 17196
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 18012 17156 18245 17184
rect 18012 17144 18018 17156
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 16850 17116 16856 17128
rect 15948 17088 16856 17116
rect 16850 17076 16856 17088
rect 16908 17116 16914 17128
rect 18500 17119 18558 17125
rect 16908 17088 18092 17116
rect 16908 17076 16914 17088
rect 14332 17020 15240 17048
rect 15289 17051 15347 17057
rect 14332 17008 14338 17020
rect 15289 17017 15301 17051
rect 15335 17048 15347 17051
rect 15470 17048 15476 17060
rect 15335 17020 15476 17048
rect 15335 17017 15347 17020
rect 15289 17011 15347 17017
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 16108 17051 16166 17057
rect 16108 17017 16120 17051
rect 16154 17048 16166 17051
rect 16758 17048 16764 17060
rect 16154 17020 16764 17048
rect 16154 17017 16166 17020
rect 16108 17011 16166 17017
rect 16758 17008 16764 17020
rect 16816 17048 16822 17060
rect 17402 17048 17408 17060
rect 16816 17020 17408 17048
rect 16816 17008 16822 17020
rect 17402 17008 17408 17020
rect 17460 17008 17466 17060
rect 18064 17048 18092 17088
rect 18500 17085 18512 17119
rect 18546 17116 18558 17119
rect 19334 17116 19340 17128
rect 18546 17088 19340 17116
rect 18546 17085 18558 17088
rect 18500 17079 18558 17085
rect 19334 17076 19340 17088
rect 19392 17116 19398 17128
rect 20162 17116 20168 17128
rect 19392 17088 20168 17116
rect 19392 17076 19398 17088
rect 20162 17076 20168 17088
rect 20220 17116 20226 17128
rect 20640 17116 20668 17147
rect 20220 17088 20668 17116
rect 20220 17076 20226 17088
rect 19794 17048 19800 17060
rect 18064 17020 19800 17048
rect 19794 17008 19800 17020
rect 19852 17008 19858 17060
rect 20438 17048 20444 17060
rect 19904 17020 20208 17048
rect 20399 17020 20444 17048
rect 14001 16983 14059 16989
rect 14001 16949 14013 16983
rect 14047 16949 14059 16983
rect 14366 16980 14372 16992
rect 14327 16952 14372 16980
rect 14001 16943 14059 16949
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 17221 16983 17279 16989
rect 17221 16980 17233 16983
rect 15068 16952 17233 16980
rect 15068 16940 15074 16952
rect 17221 16949 17233 16952
rect 17267 16949 17279 16983
rect 17494 16980 17500 16992
rect 17455 16952 17500 16980
rect 17221 16943 17279 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 17586 16940 17592 16992
rect 17644 16980 17650 16992
rect 19904 16989 19932 17020
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 17644 16952 19901 16980
rect 17644 16940 17650 16952
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 20070 16980 20076 16992
rect 20031 16952 20076 16980
rect 19889 16943 19947 16949
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20180 16980 20208 17020
rect 20438 17008 20444 17020
rect 20496 17008 20502 17060
rect 20533 16983 20591 16989
rect 20533 16980 20545 16983
rect 20180 16952 20545 16980
rect 20533 16949 20545 16952
rect 20579 16949 20591 16983
rect 20533 16943 20591 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 4304 16748 4445 16776
rect 4304 16736 4310 16748
rect 4433 16745 4445 16748
rect 4479 16745 4491 16779
rect 4433 16739 4491 16745
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 4801 16779 4859 16785
rect 4801 16776 4813 16779
rect 4764 16748 4813 16776
rect 4764 16736 4770 16748
rect 4801 16745 4813 16748
rect 4847 16745 4859 16779
rect 4801 16739 4859 16745
rect 4890 16736 4896 16788
rect 4948 16736 4954 16788
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16776 5963 16779
rect 6457 16779 6515 16785
rect 6457 16776 6469 16779
rect 5951 16748 6469 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 6457 16745 6469 16748
rect 6503 16745 6515 16779
rect 6457 16739 6515 16745
rect 6730 16736 6736 16788
rect 6788 16776 6794 16788
rect 7558 16776 7564 16788
rect 6788 16748 7564 16776
rect 6788 16736 6794 16748
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8297 16779 8355 16785
rect 8297 16745 8309 16779
rect 8343 16776 8355 16779
rect 10502 16776 10508 16788
rect 8343 16748 10088 16776
rect 10463 16748 10508 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 4908 16708 4936 16736
rect 1412 16680 4936 16708
rect 5813 16711 5871 16717
rect 1412 16649 1440 16680
rect 5813 16677 5825 16711
rect 5859 16708 5871 16711
rect 8202 16708 8208 16720
rect 5859 16680 8208 16708
rect 5859 16677 5871 16680
rect 5813 16671 5871 16677
rect 8202 16668 8208 16680
rect 8260 16668 8266 16720
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 8665 16711 8723 16717
rect 8665 16708 8677 16711
rect 8628 16680 8677 16708
rect 8628 16668 8634 16680
rect 8665 16677 8677 16680
rect 8711 16708 8723 16711
rect 9214 16708 9220 16720
rect 8711 16680 9220 16708
rect 8711 16677 8723 16680
rect 8665 16671 8723 16677
rect 9214 16668 9220 16680
rect 9272 16668 9278 16720
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16609 1455 16643
rect 1397 16603 1455 16609
rect 2216 16643 2274 16649
rect 2216 16609 2228 16643
rect 2262 16640 2274 16643
rect 3050 16640 3056 16652
rect 2262 16612 3056 16640
rect 2262 16609 2274 16612
rect 2216 16603 2274 16609
rect 3050 16600 3056 16612
rect 3108 16640 3114 16652
rect 3878 16640 3884 16652
rect 3108 16612 3884 16640
rect 3108 16600 3114 16612
rect 3878 16600 3884 16612
rect 3936 16600 3942 16652
rect 4893 16643 4951 16649
rect 4893 16609 4905 16643
rect 4939 16640 4951 16643
rect 5074 16640 5080 16652
rect 4939 16612 5080 16640
rect 4939 16609 4951 16612
rect 4893 16603 4951 16609
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 5902 16600 5908 16652
rect 5960 16640 5966 16652
rect 6730 16640 6736 16652
rect 5960 16612 6736 16640
rect 5960 16600 5966 16612
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16640 6883 16643
rect 7374 16640 7380 16652
rect 6871 16612 7380 16640
rect 6871 16609 6883 16612
rect 6825 16603 6883 16609
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 7558 16600 7564 16652
rect 7616 16640 7622 16652
rect 8757 16643 8815 16649
rect 8757 16640 8769 16643
rect 7616 16612 8769 16640
rect 7616 16600 7622 16612
rect 8757 16609 8769 16612
rect 8803 16609 8815 16643
rect 10060 16640 10088 16748
rect 10502 16736 10508 16748
rect 10560 16736 10566 16788
rect 10962 16776 10968 16788
rect 10923 16748 10968 16776
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 11517 16779 11575 16785
rect 11517 16745 11529 16779
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 10873 16711 10931 16717
rect 10873 16677 10885 16711
rect 10919 16708 10931 16711
rect 11532 16708 11560 16739
rect 11698 16736 11704 16788
rect 11756 16776 11762 16788
rect 12250 16776 12256 16788
rect 11756 16748 12256 16776
rect 11756 16736 11762 16748
rect 12250 16736 12256 16748
rect 12308 16776 12314 16788
rect 14274 16776 14280 16788
rect 12308 16748 14280 16776
rect 12308 16736 12314 16748
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 14516 16748 14657 16776
rect 14516 16736 14522 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 15657 16779 15715 16785
rect 15657 16745 15669 16779
rect 15703 16776 15715 16779
rect 16666 16776 16672 16788
rect 15703 16748 16672 16776
rect 15703 16745 15715 16748
rect 15657 16739 15715 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 17402 16776 17408 16788
rect 17363 16748 17408 16776
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16776 18291 16779
rect 18506 16776 18512 16788
rect 18279 16748 18512 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16776 18659 16779
rect 18690 16776 18696 16788
rect 18647 16748 18696 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 18969 16779 19027 16785
rect 18969 16745 18981 16779
rect 19015 16776 19027 16779
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 19015 16748 19625 16776
rect 19015 16745 19027 16748
rect 18969 16739 19027 16745
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 10919 16680 11560 16708
rect 11977 16711 12035 16717
rect 10919 16677 10931 16680
rect 10873 16671 10931 16677
rect 11977 16677 11989 16711
rect 12023 16708 12035 16711
rect 12710 16708 12716 16720
rect 12023 16680 12716 16708
rect 12023 16677 12035 16680
rect 11977 16671 12035 16677
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 12805 16711 12863 16717
rect 12805 16677 12817 16711
rect 12851 16708 12863 16711
rect 14826 16708 14832 16720
rect 12851 16680 14832 16708
rect 12851 16677 12863 16680
rect 12805 16671 12863 16677
rect 14826 16668 14832 16680
rect 14884 16668 14890 16720
rect 19061 16711 19119 16717
rect 19061 16677 19073 16711
rect 19107 16708 19119 16711
rect 20070 16708 20076 16720
rect 19107 16680 20076 16708
rect 19107 16677 19119 16680
rect 19061 16671 19119 16677
rect 20070 16668 20076 16680
rect 20128 16668 20134 16720
rect 11422 16640 11428 16652
rect 10060 16612 11428 16640
rect 8757 16603 8815 16609
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11756 16612 11897 16640
rect 11756 16600 11762 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 13532 16643 13590 16649
rect 13532 16609 13544 16643
rect 13578 16640 13590 16643
rect 15010 16640 15016 16652
rect 13578 16612 15016 16640
rect 13578 16609 13590 16612
rect 13532 16603 13590 16609
rect 15010 16600 15016 16612
rect 15068 16600 15074 16652
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15930 16600 15936 16652
rect 15988 16640 15994 16652
rect 16281 16643 16339 16649
rect 16281 16640 16293 16643
rect 15988 16612 16293 16640
rect 15988 16600 15994 16612
rect 16281 16609 16293 16612
rect 16327 16609 16339 16643
rect 16281 16603 16339 16609
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 17862 16640 17868 16652
rect 16724 16612 17868 16640
rect 16724 16600 16730 16612
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16640 18107 16643
rect 19426 16640 19432 16652
rect 18095 16612 19432 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 19426 16600 19432 16612
rect 19484 16600 19490 16652
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 19981 16643 20039 16649
rect 19852 16612 19932 16640
rect 19852 16600 19858 16612
rect 1946 16572 1952 16584
rect 1907 16544 1952 16572
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 4982 16572 4988 16584
rect 4943 16544 4988 16572
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 5810 16532 5816 16584
rect 5868 16572 5874 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5868 16544 6009 16572
rect 5868 16532 5874 16544
rect 5997 16541 6009 16544
rect 6043 16541 6055 16575
rect 6748 16572 6776 16600
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6748 16544 6929 16572
rect 5997 16535 6055 16541
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 8849 16575 8907 16581
rect 8849 16541 8861 16575
rect 8895 16541 8907 16575
rect 8849 16535 8907 16541
rect 8947 16544 10088 16572
rect 1578 16504 1584 16516
rect 1539 16476 1584 16504
rect 1578 16464 1584 16476
rect 1636 16464 1642 16516
rect 5166 16464 5172 16516
rect 5224 16504 5230 16516
rect 7024 16504 7052 16535
rect 5224 16476 7052 16504
rect 5224 16464 5230 16476
rect 7374 16464 7380 16516
rect 7432 16504 7438 16516
rect 8570 16504 8576 16516
rect 7432 16476 8576 16504
rect 7432 16464 7438 16476
rect 8570 16464 8576 16476
rect 8628 16464 8634 16516
rect 8662 16464 8668 16516
rect 8720 16504 8726 16516
rect 8864 16504 8892 16535
rect 8720 16476 8892 16504
rect 8720 16464 8726 16476
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3329 16439 3387 16445
rect 3329 16436 3341 16439
rect 3016 16408 3341 16436
rect 3016 16396 3022 16408
rect 3329 16405 3341 16408
rect 3375 16405 3387 16439
rect 3329 16399 3387 16405
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5445 16439 5503 16445
rect 5445 16436 5457 16439
rect 5040 16408 5457 16436
rect 5040 16396 5046 16408
rect 5445 16405 5457 16408
rect 5491 16405 5503 16439
rect 5445 16399 5503 16405
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 8947 16436 8975 16544
rect 10060 16504 10088 16544
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10962 16572 10968 16584
rect 10192 16544 10968 16572
rect 10192 16532 10198 16544
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11146 16572 11152 16584
rect 11107 16544 11152 16572
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 12032 16544 12081 16572
rect 12032 16532 12038 16544
rect 12069 16541 12081 16544
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 13262 16572 13268 16584
rect 12584 16544 13268 16572
rect 12584 16532 12590 16544
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16025 16575 16083 16581
rect 16025 16572 16037 16575
rect 15896 16544 16037 16572
rect 15896 16532 15902 16544
rect 16025 16541 16037 16544
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16572 19303 16575
rect 19610 16572 19616 16584
rect 19291 16544 19616 16572
rect 19291 16541 19303 16544
rect 19245 16535 19303 16541
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 19904 16572 19932 16612
rect 19981 16609 19993 16643
rect 20027 16640 20039 16643
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 20027 16612 20913 16640
rect 20027 16609 20039 16612
rect 19981 16603 20039 16609
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 20073 16575 20131 16581
rect 20073 16572 20085 16575
rect 19904 16544 20085 16572
rect 20073 16541 20085 16544
rect 20119 16541 20131 16575
rect 20073 16535 20131 16541
rect 20162 16532 20168 16584
rect 20220 16572 20226 16584
rect 20220 16544 20265 16572
rect 20220 16532 20226 16544
rect 20714 16504 20720 16516
rect 10060 16476 10640 16504
rect 5592 16408 8975 16436
rect 5592 16396 5598 16408
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 10410 16436 10416 16448
rect 9640 16408 10416 16436
rect 9640 16396 9646 16408
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 10612 16436 10640 16476
rect 16960 16476 20720 16504
rect 15746 16436 15752 16448
rect 10612 16408 15752 16436
rect 15746 16396 15752 16408
rect 15804 16396 15810 16448
rect 16390 16396 16396 16448
rect 16448 16436 16454 16448
rect 16960 16436 16988 16476
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 16448 16408 16988 16436
rect 16448 16396 16454 16408
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 19886 16436 19892 16448
rect 17276 16408 19892 16436
rect 17276 16396 17282 16408
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 3878 16232 3884 16244
rect 3839 16204 3884 16232
rect 3878 16192 3884 16204
rect 3936 16192 3942 16244
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 5350 16232 5356 16244
rect 4212 16204 5356 16232
rect 4212 16192 4218 16204
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 11606 16232 11612 16244
rect 8720 16204 11612 16232
rect 8720 16192 8726 16204
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 11698 16192 11704 16244
rect 11756 16192 11762 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 12768 16204 13461 16232
rect 12768 16192 12774 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 13449 16195 13507 16201
rect 14366 16192 14372 16244
rect 14424 16232 14430 16244
rect 14461 16235 14519 16241
rect 14461 16232 14473 16235
rect 14424 16204 14473 16232
rect 14424 16192 14430 16204
rect 14461 16201 14473 16204
rect 14507 16201 14519 16235
rect 14461 16195 14519 16201
rect 16209 16235 16267 16241
rect 16209 16201 16221 16235
rect 16255 16232 16267 16235
rect 16298 16232 16304 16244
rect 16255 16204 16304 16232
rect 16255 16201 16267 16204
rect 16209 16195 16267 16201
rect 16298 16192 16304 16204
rect 16356 16192 16362 16244
rect 16666 16192 16672 16244
rect 16724 16192 16730 16244
rect 16758 16192 16764 16244
rect 16816 16192 16822 16244
rect 17589 16235 17647 16241
rect 17589 16201 17601 16235
rect 17635 16232 17647 16235
rect 18417 16235 18475 16241
rect 17635 16204 18368 16232
rect 17635 16201 17647 16204
rect 17589 16195 17647 16201
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 3896 16096 3924 16192
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 7282 16164 7288 16176
rect 4120 16136 7288 16164
rect 4120 16124 4126 16136
rect 7282 16124 7288 16136
rect 7340 16124 7346 16176
rect 11514 16124 11520 16176
rect 11572 16164 11578 16176
rect 11716 16164 11744 16192
rect 11572 16136 11744 16164
rect 11572 16124 11578 16136
rect 12526 16124 12532 16176
rect 12584 16164 12590 16176
rect 13906 16164 13912 16176
rect 12584 16136 13912 16164
rect 12584 16124 12590 16136
rect 13906 16124 13912 16136
rect 13964 16164 13970 16176
rect 15841 16167 15899 16173
rect 13964 16136 15792 16164
rect 13964 16124 13970 16136
rect 4709 16099 4767 16105
rect 4709 16096 4721 16099
rect 2004 16068 2544 16096
rect 3896 16068 4721 16096
rect 2004 16056 2010 16068
rect 2516 16040 2544 16068
rect 4709 16065 4721 16068
rect 4755 16065 4767 16099
rect 5810 16096 5816 16108
rect 5771 16068 5816 16096
rect 4709 16059 4767 16065
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 10042 16096 10048 16108
rect 10003 16068 10048 16096
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 11882 16096 11888 16108
rect 11756 16068 11888 16096
rect 11756 16056 11762 16068
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 12986 16096 12992 16108
rect 12947 16068 12992 16096
rect 12986 16056 12992 16068
rect 13044 16096 13050 16108
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13044 16068 14013 16096
rect 13044 16056 13050 16068
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 15010 16096 15016 16108
rect 14971 16068 15016 16096
rect 14001 16059 14059 16065
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 2314 16028 2320 16040
rect 1811 16000 2320 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2498 16028 2504 16040
rect 2459 16000 2504 16028
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 4982 16028 4988 16040
rect 4663 16000 4988 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4982 15988 4988 16000
rect 5040 15988 5046 16040
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 16028 5595 16031
rect 5718 16028 5724 16040
rect 5583 16000 5724 16028
rect 5583 15997 5595 16000
rect 5537 15991 5595 15997
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 8662 16037 8668 16040
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 8656 15991 8668 16037
rect 8720 16028 8726 16040
rect 8720 16000 8756 16028
rect 2038 15960 2044 15972
rect 1999 15932 2044 15960
rect 2038 15920 2044 15932
rect 2096 15920 2102 15972
rect 2768 15963 2826 15969
rect 2768 15929 2780 15963
rect 2814 15960 2826 15963
rect 4062 15960 4068 15972
rect 2814 15932 4068 15960
rect 2814 15929 2826 15932
rect 2768 15923 2826 15929
rect 4062 15920 4068 15932
rect 4120 15920 4126 15972
rect 4525 15963 4583 15969
rect 4525 15929 4537 15963
rect 4571 15960 4583 15963
rect 4571 15932 5212 15960
rect 4571 15929 4583 15932
rect 4525 15923 4583 15929
rect 1486 15852 1492 15904
rect 1544 15892 1550 15904
rect 3326 15892 3332 15904
rect 1544 15864 3332 15892
rect 1544 15852 1550 15864
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4154 15892 4160 15904
rect 4115 15864 4160 15892
rect 4154 15852 4160 15864
rect 4212 15852 4218 15904
rect 5184 15901 5212 15932
rect 5442 15920 5448 15972
rect 5500 15960 5506 15972
rect 5629 15963 5687 15969
rect 5629 15960 5641 15963
rect 5500 15932 5641 15960
rect 5500 15920 5506 15932
rect 5629 15929 5641 15932
rect 5675 15960 5687 15963
rect 8404 15960 8432 15991
rect 8662 15988 8668 15991
rect 8720 15988 8726 16000
rect 8846 15960 8852 15972
rect 5675 15932 7687 15960
rect 8404 15932 8852 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15861 5227 15895
rect 7006 15892 7012 15904
rect 6967 15864 7012 15892
rect 5169 15855 5227 15861
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 7374 15892 7380 15904
rect 7335 15864 7380 15892
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 7659 15892 7687 15932
rect 8846 15920 8852 15932
rect 8904 15960 8910 15972
rect 10060 15960 10088 16056
rect 10312 16031 10370 16037
rect 10312 16028 10324 16031
rect 8904 15932 10088 15960
rect 10244 16000 10324 16028
rect 8904 15920 8910 15932
rect 9490 15892 9496 15904
rect 7524 15864 7569 15892
rect 7659 15864 9496 15892
rect 7524 15852 7530 15864
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 10244 15892 10272 16000
rect 10312 15997 10324 16000
rect 10358 16028 10370 16031
rect 11974 16028 11980 16040
rect 10358 16000 11980 16028
rect 10358 15997 10370 16000
rect 10312 15991 10370 15997
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12676 16000 12909 16028
rect 12676 15988 12682 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 14826 16028 14832 16040
rect 14787 16000 14832 16028
rect 12897 15991 12955 15997
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15654 16028 15660 16040
rect 15615 16000 15660 16028
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 15764 16028 15792 16136
rect 15841 16133 15853 16167
rect 15887 16164 15899 16167
rect 16684 16164 16712 16192
rect 15887 16136 16712 16164
rect 15887 16133 15899 16136
rect 15841 16127 15899 16133
rect 16776 16105 16804 16192
rect 18340 16164 18368 16204
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 19058 16232 19064 16244
rect 18463 16204 19064 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 18782 16164 18788 16176
rect 18340 16136 18788 16164
rect 18782 16124 18788 16136
rect 18840 16124 18846 16176
rect 16761 16099 16819 16105
rect 16761 16065 16773 16099
rect 16807 16065 16819 16099
rect 16761 16059 16819 16065
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18690 16096 18696 16108
rect 18012 16068 18696 16096
rect 18012 16056 18018 16068
rect 18690 16056 18696 16068
rect 18748 16096 18754 16108
rect 18748 16068 18828 16096
rect 18748 16056 18754 16068
rect 17405 16031 17463 16037
rect 17405 16028 17417 16031
rect 15764 16000 17417 16028
rect 17405 15997 17417 16000
rect 17451 16028 17463 16031
rect 17678 16028 17684 16040
rect 17451 16000 17684 16028
rect 17451 15997 17463 16000
rect 17405 15991 17463 15997
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 18800 16037 18828 16068
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 15997 18291 16031
rect 18233 15991 18291 15997
rect 18785 16031 18843 16037
rect 18785 15997 18797 16031
rect 18831 15997 18843 16031
rect 18785 15991 18843 15997
rect 19052 16031 19110 16037
rect 19052 15997 19064 16031
rect 19098 16028 19110 16031
rect 19610 16028 19616 16040
rect 19098 16000 19616 16028
rect 19098 15997 19110 16000
rect 19052 15991 19110 15997
rect 12805 15963 12863 15969
rect 12805 15929 12817 15963
rect 12851 15960 12863 15963
rect 12986 15960 12992 15972
rect 12851 15932 12992 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 12986 15920 12992 15932
rect 13044 15920 13050 15972
rect 13817 15963 13875 15969
rect 13817 15929 13829 15963
rect 13863 15960 13875 15963
rect 14921 15963 14979 15969
rect 13863 15932 14872 15960
rect 13863 15929 13875 15932
rect 13817 15923 13875 15929
rect 9815 15864 10272 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11422 15892 11428 15904
rect 11204 15864 11428 15892
rect 11204 15852 11210 15864
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 11885 15895 11943 15901
rect 11885 15861 11897 15895
rect 11931 15892 11943 15895
rect 12158 15892 12164 15904
rect 11931 15864 12164 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 13909 15895 13967 15901
rect 12492 15864 12537 15892
rect 12492 15852 12498 15864
rect 13909 15861 13921 15895
rect 13955 15892 13967 15895
rect 14458 15892 14464 15904
rect 13955 15864 14464 15892
rect 13955 15861 13967 15864
rect 13909 15855 13967 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 14844 15892 14872 15932
rect 14921 15929 14933 15963
rect 14967 15960 14979 15963
rect 15010 15960 15016 15972
rect 14967 15932 15016 15960
rect 14967 15929 14979 15932
rect 14921 15923 14979 15929
rect 15010 15920 15016 15932
rect 15068 15960 15074 15972
rect 17218 15960 17224 15972
rect 15068 15932 17224 15960
rect 15068 15920 15074 15932
rect 17218 15920 17224 15932
rect 17276 15920 17282 15972
rect 18248 15960 18276 15991
rect 19610 15988 19616 16000
rect 19668 15988 19674 16040
rect 20441 16031 20499 16037
rect 20441 16028 20453 16031
rect 19720 16000 20453 16028
rect 19518 15960 19524 15972
rect 18248 15932 19524 15960
rect 19518 15920 19524 15932
rect 19576 15920 19582 15972
rect 16114 15892 16120 15904
rect 14844 15864 16120 15892
rect 16114 15852 16120 15864
rect 16172 15892 16178 15904
rect 16390 15892 16396 15904
rect 16172 15864 16396 15892
rect 16172 15852 16178 15864
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 16482 15852 16488 15904
rect 16540 15892 16546 15904
rect 16577 15895 16635 15901
rect 16577 15892 16589 15895
rect 16540 15864 16589 15892
rect 16540 15852 16546 15864
rect 16577 15861 16589 15864
rect 16623 15861 16635 15895
rect 16577 15855 16635 15861
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 16724 15864 16769 15892
rect 16724 15852 16730 15864
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 19720 15892 19748 16000
rect 20441 15997 20453 16000
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 19794 15920 19800 15972
rect 19852 15960 19858 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 19852 15932 20729 15960
rect 19852 15920 19858 15932
rect 20717 15929 20729 15932
rect 20763 15929 20775 15963
rect 20717 15923 20775 15929
rect 20162 15892 20168 15904
rect 17092 15864 19748 15892
rect 20123 15864 20168 15892
rect 17092 15852 17098 15864
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 2777 15691 2835 15697
rect 2777 15657 2789 15691
rect 2823 15688 2835 15691
rect 4154 15688 4160 15700
rect 2823 15660 4160 15688
rect 2823 15657 2835 15660
rect 2777 15651 2835 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 5721 15691 5779 15697
rect 5721 15688 5733 15691
rect 4264 15660 5733 15688
rect 4062 15580 4068 15632
rect 4120 15620 4126 15632
rect 4264 15620 4292 15660
rect 5721 15657 5733 15660
rect 5767 15688 5779 15691
rect 5810 15688 5816 15700
rect 5767 15660 5816 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 5810 15648 5816 15660
rect 5868 15648 5874 15700
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7524 15660 7849 15688
rect 7524 15648 7530 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 8202 15688 8208 15700
rect 8163 15660 8208 15688
rect 7837 15651 7895 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8846 15688 8852 15700
rect 8807 15660 8852 15688
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 11793 15691 11851 15697
rect 11793 15688 11805 15691
rect 11572 15660 11805 15688
rect 11572 15648 11578 15660
rect 11793 15657 11805 15660
rect 11839 15657 11851 15691
rect 12158 15688 12164 15700
rect 12119 15660 12164 15688
rect 11793 15651 11851 15657
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 15933 15691 15991 15697
rect 15933 15688 15945 15691
rect 12268 15660 15945 15688
rect 4120 15592 4292 15620
rect 4608 15623 4666 15629
rect 4120 15580 4126 15592
rect 4608 15589 4620 15623
rect 4654 15620 4666 15623
rect 5166 15620 5172 15632
rect 4654 15592 5172 15620
rect 4654 15589 4666 15592
rect 4608 15583 4666 15589
rect 5166 15580 5172 15592
rect 5224 15580 5230 15632
rect 7098 15580 7104 15632
rect 7156 15620 7162 15632
rect 8297 15623 8355 15629
rect 8297 15620 8309 15623
rect 7156 15592 8309 15620
rect 7156 15580 7162 15592
rect 8297 15589 8309 15592
rect 8343 15620 8355 15623
rect 8570 15620 8576 15632
rect 8343 15592 8576 15620
rect 8343 15589 8355 15592
rect 8297 15583 8355 15589
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 8754 15580 8760 15632
rect 8812 15620 8818 15632
rect 9950 15620 9956 15632
rect 8812 15592 9956 15620
rect 8812 15580 8818 15592
rect 9950 15580 9956 15592
rect 10008 15580 10014 15632
rect 10404 15623 10462 15629
rect 10404 15589 10416 15623
rect 10450 15620 10462 15623
rect 11422 15620 11428 15632
rect 10450 15592 11428 15620
rect 10450 15589 10462 15592
rect 10404 15583 10462 15589
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 12268 15620 12296 15660
rect 15933 15657 15945 15660
rect 15979 15657 15991 15691
rect 16482 15688 16488 15700
rect 16443 15660 16488 15688
rect 15933 15651 15991 15657
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 16853 15691 16911 15697
rect 16853 15657 16865 15691
rect 16899 15688 16911 15691
rect 17494 15688 17500 15700
rect 16899 15660 17500 15688
rect 16899 15657 16911 15660
rect 16853 15651 16911 15657
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 18969 15691 19027 15697
rect 18969 15657 18981 15691
rect 19015 15688 19027 15691
rect 19242 15688 19248 15700
rect 19015 15660 19248 15688
rect 19015 15657 19027 15660
rect 18969 15651 19027 15657
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 11808 15592 12296 15620
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 2038 15552 2044 15564
rect 1811 15524 2044 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2682 15552 2688 15564
rect 2643 15524 2688 15552
rect 2682 15512 2688 15524
rect 2740 15512 2746 15564
rect 3329 15555 3387 15561
rect 3329 15521 3341 15555
rect 3375 15521 3387 15555
rect 6181 15555 6239 15561
rect 6181 15552 6193 15555
rect 3329 15515 3387 15521
rect 4356 15524 6193 15552
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3344 15348 3372 15515
rect 4246 15444 4252 15496
rect 4304 15484 4310 15496
rect 4356 15493 4384 15524
rect 6181 15521 6193 15524
rect 6227 15552 6239 15555
rect 6270 15552 6276 15564
rect 6227 15524 6276 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 6448 15555 6506 15561
rect 6448 15521 6460 15555
rect 6494 15552 6506 15555
rect 7742 15552 7748 15564
rect 6494 15524 7748 15552
rect 6494 15521 6506 15524
rect 6448 15515 6506 15521
rect 7742 15512 7748 15524
rect 7800 15552 7806 15564
rect 7800 15524 8432 15552
rect 7800 15512 7806 15524
rect 8404 15493 8432 15524
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8536 15524 9045 15552
rect 8536 15512 8542 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 10100 15524 10149 15552
rect 10100 15512 10106 15524
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 11808 15552 11836 15592
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 15841 15623 15899 15629
rect 15841 15620 15853 15623
rect 12492 15592 15853 15620
rect 12492 15580 12498 15592
rect 15841 15589 15853 15592
rect 15887 15620 15899 15623
rect 17586 15620 17592 15632
rect 15887 15592 17592 15620
rect 15887 15589 15899 15592
rect 15841 15583 15899 15589
rect 17586 15580 17592 15592
rect 17644 15580 17650 15632
rect 18049 15623 18107 15629
rect 18049 15589 18061 15623
rect 18095 15620 18107 15623
rect 19058 15620 19064 15632
rect 18095 15592 19064 15620
rect 18095 15589 18107 15592
rect 18049 15583 18107 15589
rect 19058 15580 19064 15592
rect 19116 15580 19122 15632
rect 10284 15524 11836 15552
rect 10284 15512 10290 15524
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 12253 15555 12311 15561
rect 12253 15552 12265 15555
rect 11940 15524 12265 15552
rect 11940 15512 11946 15524
rect 12253 15521 12265 15524
rect 12299 15552 12311 15555
rect 12618 15552 12624 15564
rect 12299 15524 12624 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 13170 15512 13176 15564
rect 13228 15552 13234 15564
rect 13532 15555 13590 15561
rect 13228 15524 13273 15552
rect 13228 15512 13234 15524
rect 13532 15521 13544 15555
rect 13578 15552 13590 15555
rect 14550 15552 14556 15564
rect 13578 15524 14556 15552
rect 13578 15521 13590 15524
rect 13532 15515 13590 15521
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 18141 15555 18199 15561
rect 16040 15524 17080 15552
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 4304 15456 4353 15484
rect 4304 15444 4310 15456
rect 4341 15453 4353 15456
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15453 8447 15487
rect 8389 15447 8447 15453
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 11664 15456 12357 15484
rect 11664 15444 11670 15456
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 13262 15484 13268 15496
rect 12345 15447 12403 15453
rect 13004 15456 13268 15484
rect 3510 15416 3516 15428
rect 3471 15388 3516 15416
rect 3510 15376 3516 15388
rect 3568 15376 3574 15428
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 7558 15416 7564 15428
rect 5408 15388 5764 15416
rect 7519 15388 7564 15416
rect 5408 15376 5414 15388
rect 5626 15348 5632 15360
rect 3344 15320 5632 15348
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 5736 15348 5764 15388
rect 7558 15376 7564 15388
rect 7616 15376 7622 15428
rect 12526 15416 12532 15428
rect 11440 15388 12532 15416
rect 11440 15348 11468 15388
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 5736 15320 11468 15348
rect 11517 15351 11575 15357
rect 11517 15317 11529 15351
rect 11563 15348 11575 15351
rect 11974 15348 11980 15360
rect 11563 15320 11980 15348
rect 11563 15317 11575 15320
rect 11517 15311 11575 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12250 15348 12256 15360
rect 12124 15320 12256 15348
rect 12124 15308 12130 15320
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 13004 15357 13032 15456
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 15930 15444 15936 15496
rect 15988 15484 15994 15496
rect 16040 15493 16068 15524
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 15988 15456 16037 15484
rect 15988 15444 15994 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 16439 15456 16804 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 14274 15376 14280 15428
rect 14332 15416 14338 15428
rect 15473 15419 15531 15425
rect 14332 15388 15424 15416
rect 14332 15376 14338 15388
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12676 15320 13001 15348
rect 12676 15308 12682 15320
rect 12989 15317 13001 15320
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 13078 15308 13084 15360
rect 13136 15348 13142 15360
rect 14645 15351 14703 15357
rect 14645 15348 14657 15351
rect 13136 15320 14657 15348
rect 13136 15308 13142 15320
rect 14645 15317 14657 15320
rect 14691 15317 14703 15351
rect 15396 15348 15424 15388
rect 15473 15385 15485 15419
rect 15519 15416 15531 15419
rect 16666 15416 16672 15428
rect 15519 15388 16672 15416
rect 15519 15385 15531 15388
rect 15473 15379 15531 15385
rect 16666 15376 16672 15388
rect 16724 15376 16730 15428
rect 16776 15416 16804 15456
rect 16850 15444 16856 15496
rect 16908 15484 16914 15496
rect 17052 15493 17080 15524
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18782 15552 18788 15564
rect 18187 15524 18788 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 19334 15552 19340 15564
rect 19295 15524 19340 15552
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19610 15512 19616 15564
rect 19668 15552 19674 15564
rect 19981 15555 20039 15561
rect 19981 15552 19993 15555
rect 19668 15524 19993 15552
rect 19668 15512 19674 15524
rect 19981 15521 19993 15524
rect 20027 15521 20039 15555
rect 19981 15515 20039 15521
rect 16945 15487 17003 15493
rect 16945 15484 16957 15487
rect 16908 15456 16957 15484
rect 16908 15444 16914 15456
rect 16945 15453 16957 15456
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 17037 15487 17095 15493
rect 17037 15453 17049 15487
rect 17083 15484 17095 15487
rect 17218 15484 17224 15496
rect 17083 15456 17224 15484
rect 17083 15453 17095 15456
rect 17037 15447 17095 15453
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15484 18383 15487
rect 19242 15484 19248 15496
rect 18371 15456 19248 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 19426 15484 19432 15496
rect 19387 15456 19432 15484
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 20165 15487 20223 15493
rect 19576 15456 19621 15484
rect 19576 15444 19582 15456
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 16776 15388 19104 15416
rect 16393 15351 16451 15357
rect 16393 15348 16405 15351
rect 15396 15320 16405 15348
rect 14645 15311 14703 15317
rect 16393 15317 16405 15320
rect 16439 15317 16451 15351
rect 16393 15311 16451 15317
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 16632 15320 17693 15348
rect 16632 15308 16638 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 19076 15348 19104 15388
rect 19150 15376 19156 15428
rect 19208 15416 19214 15428
rect 20180 15416 20208 15447
rect 20254 15444 20260 15496
rect 20312 15484 20318 15496
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 20312 15456 20913 15484
rect 20312 15444 20318 15456
rect 20901 15453 20913 15456
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 19208 15388 20208 15416
rect 19208 15376 19214 15388
rect 20070 15348 20076 15360
rect 19076 15320 20076 15348
rect 17681 15311 17739 15317
rect 20070 15308 20076 15320
rect 20128 15348 20134 15360
rect 20346 15348 20352 15360
rect 20128 15320 20352 15348
rect 20128 15308 20134 15320
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 2409 15147 2467 15153
rect 2409 15113 2421 15147
rect 2455 15144 2467 15147
rect 2682 15144 2688 15156
rect 2455 15116 2688 15144
rect 2455 15113 2467 15116
rect 2409 15107 2467 15113
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 7374 15104 7380 15156
rect 7432 15144 7438 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7432 15116 7849 15144
rect 7432 15104 7438 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 8665 15147 8723 15153
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 11698 15144 11704 15156
rect 8711 15116 11704 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12805 15147 12863 15153
rect 12805 15113 12817 15147
rect 12851 15144 12863 15147
rect 14550 15144 14556 15156
rect 12851 15116 14412 15144
rect 14511 15116 14556 15144
rect 12851 15113 12863 15116
rect 12805 15107 12863 15113
rect 1946 15076 1952 15088
rect 1907 15048 1952 15076
rect 1946 15036 1952 15048
rect 2004 15036 2010 15088
rect 6178 15036 6184 15088
rect 6236 15076 6242 15088
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 6236 15048 6837 15076
rect 6236 15036 6242 15048
rect 6825 15045 6837 15048
rect 6871 15045 6883 15079
rect 9214 15076 9220 15088
rect 6825 15039 6883 15045
rect 6923 15048 9220 15076
rect 3050 15008 3056 15020
rect 3011 14980 3056 15008
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 4062 15008 4068 15020
rect 4023 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 5408 14980 5825 15008
rect 5408 14968 5414 14980
rect 5813 14977 5825 14980
rect 5859 14977 5871 15011
rect 5813 14971 5871 14977
rect 6089 15011 6147 15017
rect 6089 14977 6101 15011
rect 6135 15008 6147 15011
rect 6923 15008 6951 15048
rect 9214 15036 9220 15048
rect 9272 15036 9278 15088
rect 11146 15076 11152 15088
rect 9508 15048 11152 15076
rect 6135 14980 6951 15008
rect 6135 14977 6147 14980
rect 6089 14971 6147 14977
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 7064 14980 7297 15008
rect 7064 14968 7070 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 7285 14971 7343 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 7742 14968 7748 15020
rect 7800 15008 7806 15020
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 7800 14980 8401 15008
rect 7800 14968 7806 14980
rect 8389 14977 8401 14980
rect 8435 14977 8447 15011
rect 8389 14971 8447 14977
rect 8570 14968 8576 15020
rect 8628 15008 8634 15020
rect 9508 15017 9536 15048
rect 11146 15036 11152 15048
rect 11204 15036 11210 15088
rect 11333 15079 11391 15085
rect 11333 15045 11345 15079
rect 11379 15076 11391 15079
rect 13078 15076 13084 15088
rect 11379 15048 13084 15076
rect 11379 15045 11391 15048
rect 11333 15039 11391 15045
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 14384 15076 14412 15116
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 15795 15116 20760 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 17218 15076 17224 15088
rect 14384 15048 15608 15076
rect 17179 15048 17224 15076
rect 9309 15011 9367 15017
rect 9309 15008 9321 15011
rect 8628 14980 9321 15008
rect 8628 14968 8634 14980
rect 9309 14977 9321 14980
rect 9355 14977 9367 15011
rect 9309 14971 9367 14977
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 14977 9551 15011
rect 10502 15008 10508 15020
rect 10463 14980 10508 15008
rect 9493 14971 9551 14977
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12250 15008 12256 15020
rect 12023 14980 12256 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 14608 14980 15393 15008
rect 14608 14968 14614 14980
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 15580 15008 15608 15048
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 18509 15079 18567 15085
rect 18509 15045 18521 15079
rect 18555 15076 18567 15079
rect 18874 15076 18880 15088
rect 18555 15048 18880 15076
rect 18555 15045 18567 15048
rect 18509 15039 18567 15045
rect 18874 15036 18880 15048
rect 18932 15036 18938 15088
rect 15657 15011 15715 15017
rect 15657 15008 15669 15011
rect 15580 14980 15669 15008
rect 15381 14971 15439 14977
rect 15657 14977 15669 14980
rect 15703 14977 15715 15011
rect 15838 15008 15844 15020
rect 15799 14980 15844 15008
rect 15657 14971 15715 14977
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 20732 15017 20760 15116
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 2406 14940 2412 14952
rect 1811 14912 2412 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 6362 14940 6368 14952
rect 5767 14912 6368 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 6457 14943 6515 14949
rect 6457 14909 6469 14943
rect 6503 14909 6515 14943
rect 6457 14903 6515 14909
rect 2777 14875 2835 14881
rect 2777 14841 2789 14875
rect 2823 14872 2835 14875
rect 3789 14875 3847 14881
rect 2823 14844 3464 14872
rect 2823 14841 2835 14844
rect 2777 14835 2835 14841
rect 2866 14804 2872 14816
rect 2827 14776 2872 14804
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 3436 14813 3464 14844
rect 3789 14841 3801 14875
rect 3835 14872 3847 14875
rect 4433 14875 4491 14881
rect 4433 14872 4445 14875
rect 3835 14844 4445 14872
rect 3835 14841 3847 14844
rect 3789 14835 3847 14841
rect 4433 14841 4445 14844
rect 4479 14841 4491 14875
rect 4433 14835 4491 14841
rect 5629 14875 5687 14881
rect 5629 14841 5641 14875
rect 5675 14872 5687 14875
rect 6089 14875 6147 14881
rect 6089 14872 6101 14875
rect 5675 14844 6101 14872
rect 5675 14841 5687 14844
rect 5629 14835 5687 14841
rect 6089 14841 6101 14844
rect 6135 14841 6147 14875
rect 6472 14872 6500 14903
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 7248 14912 7665 14940
rect 7248 14900 7254 14912
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 8260 14912 9229 14940
rect 8260 14900 8266 14912
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 12434 14940 12440 14952
rect 10367 14912 12440 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12621 14943 12679 14949
rect 12621 14909 12633 14943
rect 12667 14909 12679 14943
rect 12621 14903 12679 14909
rect 8478 14872 8484 14884
rect 6472 14844 8484 14872
rect 6089 14835 6147 14841
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 11793 14875 11851 14881
rect 11793 14872 11805 14875
rect 8864 14844 11805 14872
rect 3421 14807 3479 14813
rect 3421 14773 3433 14807
rect 3467 14773 3479 14807
rect 3421 14767 3479 14773
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 3881 14807 3939 14813
rect 3881 14804 3893 14807
rect 3752 14776 3893 14804
rect 3752 14764 3758 14776
rect 3881 14773 3893 14776
rect 3927 14773 3939 14807
rect 5258 14804 5264 14816
rect 5219 14776 5264 14804
rect 3881 14767 3939 14773
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 7190 14804 7196 14816
rect 7151 14776 7196 14804
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 8202 14804 8208 14816
rect 7699 14776 8208 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8864 14813 8892 14844
rect 11793 14841 11805 14844
rect 11839 14841 11851 14875
rect 12636 14872 12664 14903
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 13173 14943 13231 14949
rect 13173 14940 13185 14943
rect 12768 14912 13185 14940
rect 12768 14900 12774 14912
rect 13173 14909 13185 14912
rect 13219 14909 13231 14943
rect 15749 14943 15807 14949
rect 15749 14940 15761 14943
rect 13173 14903 13231 14909
rect 13280 14912 15761 14940
rect 13280 14872 13308 14912
rect 15749 14909 15761 14912
rect 15795 14909 15807 14943
rect 15749 14903 15807 14909
rect 16040 14912 18276 14940
rect 12636 14844 13308 14872
rect 13440 14875 13498 14881
rect 11793 14835 11851 14841
rect 13440 14841 13452 14875
rect 13486 14872 13498 14875
rect 13998 14872 14004 14884
rect 13486 14844 14004 14872
rect 13486 14841 13498 14844
rect 13440 14835 13498 14841
rect 13998 14832 14004 14844
rect 14056 14832 14062 14884
rect 16040 14872 16068 14912
rect 14844 14844 16068 14872
rect 16108 14875 16166 14881
rect 8297 14807 8355 14813
rect 8297 14773 8309 14807
rect 8343 14804 8355 14807
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8343 14776 8677 14804
rect 8343 14773 8355 14776
rect 8297 14767 8355 14773
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14773 8907 14807
rect 9950 14804 9956 14816
rect 9911 14776 9956 14804
rect 8849 14767 8907 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10410 14804 10416 14816
rect 10371 14776 10416 14804
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 14844 14813 14872 14844
rect 16108 14841 16120 14875
rect 16154 14872 16166 14875
rect 16758 14872 16764 14884
rect 16154 14844 16764 14872
rect 16154 14841 16166 14844
rect 16108 14835 16166 14841
rect 16758 14832 16764 14844
rect 16816 14832 16822 14884
rect 17862 14872 17868 14884
rect 17328 14844 17868 14872
rect 14829 14807 14887 14813
rect 14829 14773 14841 14807
rect 14875 14773 14887 14807
rect 15194 14804 15200 14816
rect 15155 14776 15200 14804
rect 14829 14767 14887 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15470 14804 15476 14816
rect 15335 14776 15476 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15657 14807 15715 14813
rect 15657 14773 15669 14807
rect 15703 14804 15715 14807
rect 17328 14804 17356 14844
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 18248 14872 18276 14912
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 18598 14940 18604 14952
rect 18380 14912 18604 14940
rect 18380 14900 18386 14912
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18690 14900 18696 14952
rect 18748 14940 18754 14952
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18748 14912 18889 14940
rect 18748 14900 18754 14912
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 20533 14943 20591 14949
rect 20533 14940 20545 14943
rect 18877 14903 18935 14909
rect 18984 14912 20545 14940
rect 18984 14872 19012 14912
rect 20533 14909 20545 14912
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 18248 14844 19012 14872
rect 19144 14875 19202 14881
rect 19144 14841 19156 14875
rect 19190 14872 19202 14875
rect 20162 14872 20168 14884
rect 19190 14844 20168 14872
rect 19190 14841 19202 14844
rect 19144 14835 19202 14841
rect 20162 14832 20168 14844
rect 20220 14832 20226 14884
rect 17494 14804 17500 14816
rect 15703 14776 17356 14804
rect 17455 14776 17500 14804
rect 15703 14773 15715 14776
rect 15657 14767 15715 14773
rect 17494 14764 17500 14776
rect 17552 14764 17558 14816
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 20257 14807 20315 14813
rect 20257 14804 20269 14807
rect 19576 14776 20269 14804
rect 19576 14764 19582 14776
rect 20257 14773 20269 14776
rect 20303 14773 20315 14807
rect 20257 14767 20315 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 2866 14600 2872 14612
rect 2823 14572 2872 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 6270 14600 6276 14612
rect 3160 14572 5856 14600
rect 198 14492 204 14544
rect 256 14532 262 14544
rect 3160 14532 3188 14572
rect 256 14504 3188 14532
rect 3237 14535 3295 14541
rect 256 14492 262 14504
rect 3237 14501 3249 14535
rect 3283 14532 3295 14535
rect 5166 14532 5172 14544
rect 3283 14504 5172 14532
rect 3283 14501 3295 14504
rect 3237 14495 3295 14501
rect 5166 14492 5172 14504
rect 5224 14492 5230 14544
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14464 1731 14467
rect 1946 14464 1952 14476
rect 1719 14436 1952 14464
rect 1719 14433 1731 14436
rect 1673 14427 1731 14433
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 3142 14464 3148 14476
rect 3103 14436 3148 14464
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3418 14424 3424 14476
rect 3476 14464 3482 14476
rect 4321 14467 4379 14473
rect 4321 14464 4333 14467
rect 3476 14436 4333 14464
rect 3476 14424 3482 14436
rect 4321 14433 4333 14436
rect 4367 14433 4379 14467
rect 4321 14427 4379 14433
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 1857 14399 1915 14405
rect 1857 14396 1869 14399
rect 1452 14368 1869 14396
rect 1452 14356 1458 14368
rect 1857 14365 1869 14368
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 3970 14396 3976 14408
rect 3375 14368 3976 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 1762 14288 1768 14340
rect 1820 14328 1826 14340
rect 2498 14328 2504 14340
rect 1820 14300 2504 14328
rect 1820 14288 1826 14300
rect 2498 14288 2504 14300
rect 2556 14328 2562 14340
rect 4080 14328 4108 14359
rect 5442 14328 5448 14340
rect 2556 14300 4108 14328
rect 5403 14300 5448 14328
rect 2556 14288 2562 14300
rect 4080 14260 4108 14300
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 4246 14260 4252 14272
rect 4080 14232 4252 14260
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 5828 14260 5856 14572
rect 5920 14572 6276 14600
rect 5920 14473 5948 14572
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 8573 14603 8631 14609
rect 8573 14569 8585 14603
rect 8619 14569 8631 14603
rect 8573 14563 8631 14569
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9306 14600 9312 14612
rect 8987 14572 9312 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 6172 14535 6230 14541
rect 6172 14501 6184 14535
rect 6218 14532 6230 14535
rect 7558 14532 7564 14544
rect 6218 14504 7564 14532
rect 6218 14501 6230 14504
rect 6172 14495 6230 14501
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 8588 14532 8616 14563
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9858 14600 9864 14612
rect 9819 14572 9864 14600
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10321 14603 10379 14609
rect 10321 14600 10333 14603
rect 10008 14572 10333 14600
rect 10008 14560 10014 14572
rect 10321 14569 10333 14572
rect 10367 14569 10379 14603
rect 12250 14600 12256 14612
rect 12211 14572 12256 14600
rect 10321 14563 10379 14569
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 14829 14603 14887 14609
rect 14829 14569 14841 14603
rect 14875 14600 14887 14603
rect 16298 14600 16304 14612
rect 14875 14572 16304 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 16758 14600 16764 14612
rect 16719 14572 16764 14600
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 19242 14600 19248 14612
rect 16868 14572 19248 14600
rect 10410 14532 10416 14544
rect 8588 14504 10416 14532
rect 10410 14492 10416 14504
rect 10468 14492 10474 14544
rect 11974 14532 11980 14544
rect 10704 14504 11980 14532
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14433 5963 14467
rect 5905 14427 5963 14433
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 10226 14464 10232 14476
rect 6512 14436 7052 14464
rect 10187 14436 10232 14464
rect 6512 14424 6518 14436
rect 7024 14396 7052 14436
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 9033 14399 9091 14405
rect 9033 14396 9045 14399
rect 7024 14368 9045 14396
rect 9033 14365 9045 14368
rect 9079 14365 9091 14399
rect 9033 14359 9091 14365
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 9180 14368 9225 14396
rect 9180 14356 9186 14368
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 9640 14368 10425 14396
rect 9640 14356 9646 14368
rect 10413 14365 10425 14368
rect 10459 14396 10471 14399
rect 10594 14396 10600 14408
rect 10459 14368 10600 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 8846 14328 8852 14340
rect 6840 14300 8852 14328
rect 6840 14260 6868 14300
rect 8846 14288 8852 14300
rect 8904 14288 8910 14340
rect 9140 14328 9168 14356
rect 10704 14328 10732 14504
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 13722 14492 13728 14544
rect 13780 14532 13786 14544
rect 15470 14532 15476 14544
rect 13780 14504 15476 14532
rect 13780 14492 13786 14504
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 15648 14535 15706 14541
rect 15648 14501 15660 14535
rect 15694 14532 15706 14535
rect 16482 14532 16488 14544
rect 15694 14504 16488 14532
rect 15694 14501 15706 14504
rect 15648 14495 15706 14501
rect 16482 14492 16488 14504
rect 16540 14532 16546 14544
rect 16868 14532 16896 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 19392 14572 19625 14600
rect 19392 14560 19398 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 19613 14563 19671 14569
rect 19981 14603 20039 14609
rect 19981 14569 19993 14603
rect 20027 14600 20039 14603
rect 20254 14600 20260 14612
rect 20027 14572 20260 14600
rect 20027 14569 20039 14572
rect 19981 14563 20039 14569
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 17310 14532 17316 14544
rect 16540 14504 16896 14532
rect 17271 14504 17316 14532
rect 16540 14492 16546 14504
rect 17310 14492 17316 14504
rect 17368 14492 17374 14544
rect 18690 14532 18696 14544
rect 17880 14504 18696 14532
rect 11146 14473 11152 14476
rect 11140 14464 11152 14473
rect 11059 14436 11152 14464
rect 11140 14427 11152 14436
rect 11204 14464 11210 14476
rect 11606 14464 11612 14476
rect 11204 14436 11612 14464
rect 11146 14424 11152 14427
rect 11204 14424 11210 14436
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12877 14467 12935 14473
rect 12877 14464 12889 14467
rect 12308 14436 12889 14464
rect 12308 14424 12314 14436
rect 12877 14433 12889 14436
rect 12923 14464 12935 14467
rect 14642 14464 14648 14476
rect 12923 14436 13860 14464
rect 14603 14436 14648 14464
rect 12923 14433 12935 14436
rect 12877 14427 12935 14433
rect 10873 14399 10931 14405
rect 10873 14365 10885 14399
rect 10919 14365 10931 14399
rect 12618 14396 12624 14408
rect 12531 14368 12624 14396
rect 10873 14359 10931 14365
rect 9140 14300 10732 14328
rect 5828 14232 6868 14260
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 7285 14263 7343 14269
rect 7285 14260 7297 14263
rect 6972 14232 7297 14260
rect 6972 14220 6978 14232
rect 7285 14229 7297 14232
rect 7331 14260 7343 14263
rect 7374 14260 7380 14272
rect 7331 14232 7380 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8202 14220 8208 14272
rect 8260 14260 8266 14272
rect 10318 14260 10324 14272
rect 8260 14232 10324 14260
rect 8260 14220 8266 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10888 14260 10916 14359
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 13832 14396 13860 14436
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14464 15439 14467
rect 15930 14464 15936 14476
rect 15427 14436 15936 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 15930 14424 15936 14436
rect 15988 14464 15994 14476
rect 15988 14436 16896 14464
rect 15988 14424 15994 14436
rect 15010 14396 15016 14408
rect 13832 14368 15016 14396
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 16868 14396 16896 14436
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 17880 14473 17908 14504
rect 18690 14492 18696 14504
rect 18748 14532 18754 14544
rect 18874 14532 18880 14544
rect 18748 14504 18880 14532
rect 18748 14492 18754 14504
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 20070 14532 20076 14544
rect 20031 14504 20076 14532
rect 20070 14492 20076 14504
rect 20128 14492 20134 14544
rect 17037 14467 17095 14473
rect 17037 14464 17049 14467
rect 17000 14436 17049 14464
rect 17000 14424 17006 14436
rect 17037 14433 17049 14436
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14433 17923 14467
rect 17865 14427 17923 14433
rect 18132 14467 18190 14473
rect 18132 14433 18144 14467
rect 18178 14464 18190 14467
rect 18506 14464 18512 14476
rect 18178 14436 18512 14464
rect 18178 14433 18190 14436
rect 18132 14427 18190 14433
rect 17218 14396 17224 14408
rect 16868 14368 17224 14396
rect 17218 14356 17224 14368
rect 17276 14396 17282 14408
rect 17880 14396 17908 14427
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 18598 14424 18604 14476
rect 18656 14464 18662 14476
rect 20254 14464 20260 14476
rect 18656 14436 20260 14464
rect 18656 14424 18662 14436
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 17276 14368 17908 14396
rect 17276 14356 17282 14368
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20220 14368 20265 14396
rect 20220 14356 20226 14368
rect 11146 14260 11152 14272
rect 10888 14232 11152 14260
rect 11146 14220 11152 14232
rect 11204 14260 11210 14272
rect 12627 14260 12655 14356
rect 13998 14328 14004 14340
rect 13959 14300 14004 14328
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 20530 14328 20536 14340
rect 18800 14300 20536 14328
rect 11204 14232 12655 14260
rect 11204 14220 11210 14232
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 18800 14260 18828 14300
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 17920 14232 18828 14260
rect 17920 14220 17926 14232
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 6825 14059 6883 14065
rect 5500 14028 6224 14056
rect 5500 14016 5506 14028
rect 2961 13991 3019 13997
rect 2961 13988 2973 13991
rect 2424 13960 2973 13988
rect 2424 13929 2452 13960
rect 2961 13957 2973 13960
rect 3007 13957 3019 13991
rect 4157 13991 4215 13997
rect 4157 13988 4169 13991
rect 2961 13951 3019 13957
rect 3436 13960 4169 13988
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13889 2467 13923
rect 2409 13883 2467 13889
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 3326 13920 3332 13932
rect 2639 13892 3332 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3436 13929 3464 13960
rect 4157 13957 4169 13960
rect 4203 13957 4215 13991
rect 4157 13951 4215 13957
rect 5721 13991 5779 13997
rect 5721 13957 5733 13991
rect 5767 13957 5779 13991
rect 5721 13951 5779 13957
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13889 3571 13923
rect 4706 13920 4712 13932
rect 4667 13892 4712 13920
rect 3513 13883 3571 13889
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 3528 13852 3556 13883
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 2096 13824 3556 13852
rect 4617 13855 4675 13861
rect 2096 13812 2102 13824
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5258 13852 5264 13864
rect 4663 13824 5264 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 5736 13852 5764 13951
rect 6196 13929 6224 14028
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7190 14056 7196 14068
rect 6871 14028 7196 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 8297 14059 8355 14065
rect 8297 14025 8309 14059
rect 8343 14056 8355 14059
rect 8478 14056 8484 14068
rect 8343 14028 8484 14056
rect 8343 14025 8355 14028
rect 8297 14019 8355 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 8846 14016 8852 14068
rect 8904 14056 8910 14068
rect 9858 14056 9864 14068
rect 8904 14028 9864 14056
rect 8904 14016 8910 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 10652 14028 11621 14056
rect 10652 14016 10658 14028
rect 11609 14025 11621 14028
rect 11655 14025 11667 14059
rect 11609 14019 11667 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 13725 14059 13783 14065
rect 12492 14028 12537 14056
rect 12492 14016 12498 14028
rect 13725 14025 13737 14059
rect 13771 14056 13783 14059
rect 15194 14056 15200 14068
rect 13771 14028 15200 14056
rect 13771 14025 13783 14028
rect 13725 14019 13783 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 15749 14059 15807 14065
rect 15749 14025 15761 14059
rect 15795 14056 15807 14059
rect 15930 14056 15936 14068
rect 15795 14028 15936 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 16942 14056 16948 14068
rect 16071 14028 16948 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 18969 14059 19027 14065
rect 18969 14025 18981 14059
rect 19015 14056 19027 14059
rect 19426 14056 19432 14068
rect 19015 14028 19432 14056
rect 19015 14025 19027 14028
rect 18969 14019 19027 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 7006 13988 7012 14000
rect 6380 13960 7012 13988
rect 6380 13929 6408 13960
rect 7006 13948 7012 13960
rect 7064 13988 7070 14000
rect 7742 13988 7748 14000
rect 7064 13960 7748 13988
rect 7064 13948 7070 13960
rect 7742 13948 7748 13960
rect 7800 13948 7806 14000
rect 11514 13948 11520 14000
rect 11572 13988 11578 14000
rect 11882 13988 11888 14000
rect 11572 13960 11888 13988
rect 11572 13948 11578 13960
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 12250 13948 12256 14000
rect 12308 13988 12314 14000
rect 12308 13960 13124 13988
rect 12308 13948 12314 13960
rect 6181 13923 6239 13929
rect 6181 13889 6193 13923
rect 6227 13889 6239 13923
rect 6181 13883 6239 13889
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7558 13920 7564 13932
rect 7515 13892 7564 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 9916 13892 10364 13920
rect 9916 13880 9922 13892
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 5736 13824 7205 13852
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 8478 13852 8484 13864
rect 8439 13824 8484 13852
rect 7193 13815 7251 13821
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 8840 13855 8898 13861
rect 8840 13821 8852 13855
rect 8886 13852 8898 13855
rect 9122 13852 9128 13864
rect 8886 13824 9128 13852
rect 8886 13821 8898 13824
rect 8840 13815 8898 13821
rect 3602 13744 3608 13796
rect 3660 13784 3666 13796
rect 6089 13787 6147 13793
rect 3660 13756 6040 13784
rect 3660 13744 3666 13756
rect 2314 13716 2320 13728
rect 2275 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 3329 13719 3387 13725
rect 3329 13685 3341 13719
rect 3375 13716 3387 13719
rect 4062 13716 4068 13728
rect 3375 13688 4068 13716
rect 3375 13685 3387 13688
rect 3329 13679 3387 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4525 13719 4583 13725
rect 4525 13685 4537 13719
rect 4571 13716 4583 13719
rect 4982 13716 4988 13728
rect 4571 13688 4988 13716
rect 4571 13685 4583 13688
rect 4525 13679 4583 13685
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 6012 13716 6040 13756
rect 6089 13753 6101 13787
rect 6135 13784 6147 13787
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 6135 13756 7849 13784
rect 6135 13753 6147 13756
rect 6089 13747 6147 13753
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 8588 13784 8616 13815
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13821 10287 13855
rect 10336 13852 10364 13892
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12032 13892 13001 13920
rect 12032 13880 12038 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 13096 13920 13124 13960
rect 13170 13948 13176 14000
rect 13228 13988 13234 14000
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 13228 13960 13461 13988
rect 13228 13948 13234 13960
rect 13449 13957 13461 13960
rect 13495 13988 13507 13991
rect 13495 13960 15976 13988
rect 13495 13957 13507 13960
rect 13449 13951 13507 13957
rect 13096 13892 13952 13920
rect 12989 13883 13047 13889
rect 12250 13852 12256 13864
rect 10336 13824 12256 13852
rect 10229 13815 10287 13821
rect 9674 13784 9680 13796
rect 8588 13756 9680 13784
rect 7837 13747 7895 13753
rect 9674 13744 9680 13756
rect 9732 13784 9738 13796
rect 10042 13784 10048 13796
rect 9732 13756 10048 13784
rect 9732 13744 9738 13756
rect 10042 13744 10048 13756
rect 10100 13784 10106 13796
rect 10244 13784 10272 13815
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12860 13824 12909 13852
rect 12860 13812 12866 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13170 13812 13176 13864
rect 13228 13852 13234 13864
rect 13633 13855 13691 13861
rect 13633 13852 13645 13855
rect 13228 13824 13645 13852
rect 13228 13812 13234 13824
rect 13633 13821 13645 13824
rect 13679 13821 13691 13855
rect 13924 13852 13952 13892
rect 13998 13880 14004 13932
rect 14056 13920 14062 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 14056 13892 14289 13920
rect 14056 13880 14062 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 15068 13892 15301 13920
rect 15068 13880 15074 13892
rect 15289 13889 15301 13892
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15948 13861 15976 13960
rect 16031 13960 18368 13988
rect 15933 13855 15991 13861
rect 13924 13824 15884 13852
rect 13633 13815 13691 13821
rect 10502 13793 10508 13796
rect 10496 13784 10508 13793
rect 10100 13756 10272 13784
rect 10428 13756 10508 13784
rect 10100 13744 10106 13756
rect 6730 13716 6736 13728
rect 6012 13688 6736 13716
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7285 13719 7343 13725
rect 7285 13716 7297 13719
rect 7248 13688 7297 13716
rect 7248 13676 7254 13688
rect 7285 13685 7297 13688
rect 7331 13685 7343 13719
rect 7285 13679 7343 13685
rect 9953 13719 10011 13725
rect 9953 13685 9965 13719
rect 9999 13716 10011 13719
rect 10428 13716 10456 13756
rect 10496 13747 10508 13756
rect 10502 13744 10508 13747
rect 10560 13744 10566 13796
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 11885 13787 11943 13793
rect 11885 13784 11897 13787
rect 10652 13756 11897 13784
rect 10652 13744 10658 13756
rect 11885 13753 11897 13756
rect 11931 13753 11943 13787
rect 11885 13747 11943 13753
rect 14093 13787 14151 13793
rect 14093 13753 14105 13787
rect 14139 13784 14151 13787
rect 15856 13784 15884 13824
rect 15933 13821 15945 13855
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 16031 13784 16059 13960
rect 16485 13923 16543 13929
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 16574 13920 16580 13932
rect 16531 13892 16580 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 16758 13920 16764 13932
rect 16715 13892 16764 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17221 13923 17279 13929
rect 17221 13920 17233 13923
rect 17184 13892 17233 13920
rect 17184 13880 17190 13892
rect 17221 13889 17233 13892
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 17402 13880 17408 13932
rect 17460 13920 17466 13932
rect 18340 13920 18368 13960
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 19981 13991 20039 13997
rect 19981 13988 19993 13991
rect 18748 13960 19993 13988
rect 18748 13948 18754 13960
rect 19981 13957 19993 13960
rect 20027 13957 20039 13991
rect 19981 13951 20039 13957
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 17460 13892 18276 13920
rect 18340 13892 19441 13920
rect 17460 13880 17466 13892
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 16356 13824 16405 13852
rect 16356 13812 16362 13824
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13852 17095 13855
rect 17954 13852 17960 13864
rect 17083 13824 17960 13852
rect 17083 13821 17095 13824
rect 17037 13815 17095 13821
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 18248 13861 18276 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 20162 13920 20168 13932
rect 19659 13892 20168 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18233 13815 18291 13821
rect 18509 13855 18567 13861
rect 18509 13821 18521 13855
rect 18555 13852 18567 13855
rect 19334 13852 19340 13864
rect 18555 13824 19340 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19444 13852 19472 13883
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20530 13920 20536 13932
rect 20491 13892 20536 13920
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 19444 13824 20453 13852
rect 20441 13821 20453 13824
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 14139 13756 14780 13784
rect 15856 13756 16059 13784
rect 14139 13753 14151 13756
rect 14093 13747 14151 13753
rect 9999 13688 10456 13716
rect 9999 13685 10011 13688
rect 9953 13679 10011 13685
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 11848 13688 12817 13716
rect 11848 13676 11854 13688
rect 12805 13685 12817 13688
rect 12851 13716 12863 13719
rect 13814 13716 13820 13728
rect 12851 13688 13820 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14182 13716 14188 13728
rect 14143 13688 14188 13716
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 14752 13725 14780 13756
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 19794 13784 19800 13796
rect 16264 13756 19800 13784
rect 16264 13744 16270 13756
rect 19794 13744 19800 13756
rect 19852 13744 19858 13796
rect 14737 13719 14795 13725
rect 14737 13685 14749 13719
rect 14783 13685 14795 13719
rect 15102 13716 15108 13728
rect 15063 13688 15108 13716
rect 14737 13679 14795 13685
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15252 13688 15297 13716
rect 15252 13676 15258 13688
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 19242 13716 19248 13728
rect 18104 13688 19248 13716
rect 18104 13676 18110 13688
rect 19242 13676 19248 13688
rect 19300 13716 19306 13728
rect 19337 13719 19395 13725
rect 19337 13716 19349 13719
rect 19300 13688 19349 13716
rect 19300 13676 19306 13688
rect 19337 13685 19349 13688
rect 19383 13685 19395 13719
rect 19337 13679 19395 13685
rect 19426 13676 19432 13728
rect 19484 13716 19490 13728
rect 20346 13716 20352 13728
rect 19484 13688 20352 13716
rect 19484 13676 19490 13688
rect 20346 13676 20352 13688
rect 20404 13676 20410 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 3145 13515 3203 13521
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 3418 13512 3424 13524
rect 3191 13484 3424 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 3602 13512 3608 13524
rect 3563 13484 3608 13512
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 4062 13512 4068 13524
rect 4023 13484 4068 13512
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 5077 13515 5135 13521
rect 5077 13512 5089 13515
rect 4571 13484 5089 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 5077 13481 5089 13484
rect 5123 13481 5135 13515
rect 5077 13475 5135 13481
rect 5258 13472 5264 13524
rect 5316 13512 5322 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 5316 13484 5457 13512
rect 5316 13472 5322 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5445 13475 5503 13481
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 7190 13512 7196 13524
rect 6227 13484 7196 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 10226 13512 10232 13524
rect 7300 13484 10088 13512
rect 10187 13484 10232 13512
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 4304 13416 6561 13444
rect 4304 13404 4310 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 6549 13407 6607 13413
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2038 13385 2044 13388
rect 2032 13376 2044 13385
rect 1999 13348 2044 13376
rect 2032 13339 2044 13348
rect 2038 13336 2044 13339
rect 2096 13336 2102 13388
rect 2590 13336 2596 13388
rect 2648 13376 2654 13388
rect 3421 13379 3479 13385
rect 2648 13348 3372 13376
rect 2648 13336 2654 13348
rect 3344 13308 3372 13348
rect 3421 13345 3433 13379
rect 3467 13376 3479 13379
rect 3510 13376 3516 13388
rect 3467 13348 3516 13376
rect 3467 13345 3479 13348
rect 3421 13339 3479 13345
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 3878 13336 3884 13388
rect 3936 13376 3942 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 3936 13348 4445 13376
rect 3936 13336 3942 13348
rect 4433 13345 4445 13348
rect 4479 13345 4491 13379
rect 7300 13376 7328 13484
rect 9950 13444 9956 13456
rect 7392 13416 9956 13444
rect 7392 13385 7420 13416
rect 9950 13404 9956 13416
rect 10008 13404 10014 13456
rect 10060 13444 10088 13484
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 10594 13512 10600 13524
rect 10555 13484 10600 13512
rect 10594 13472 10600 13484
rect 10652 13472 10658 13524
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 11241 13515 11299 13521
rect 11241 13512 11253 13515
rect 10735 13484 11253 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 11241 13481 11253 13484
rect 11287 13481 11299 13515
rect 11241 13475 11299 13481
rect 11609 13515 11667 13521
rect 11609 13481 11621 13515
rect 11655 13512 11667 13515
rect 11882 13512 11888 13524
rect 11655 13484 11888 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 16117 13515 16175 13521
rect 12492 13484 16068 13512
rect 12492 13472 12498 13484
rect 11514 13444 11520 13456
rect 10060 13416 11520 13444
rect 11514 13404 11520 13416
rect 11572 13404 11578 13456
rect 11701 13447 11759 13453
rect 11701 13413 11713 13447
rect 11747 13444 11759 13447
rect 12805 13447 12863 13453
rect 12805 13444 12817 13447
rect 11747 13416 12817 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 12805 13413 12817 13416
rect 12851 13413 12863 13447
rect 12805 13407 12863 13413
rect 4433 13339 4491 13345
rect 5276 13348 7328 13376
rect 7377 13379 7435 13385
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 3344 13280 4629 13308
rect 4617 13277 4629 13280
rect 4663 13308 4675 13311
rect 4706 13308 4712 13320
rect 4663 13280 4712 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 3786 13200 3792 13252
rect 3844 13240 3850 13252
rect 4062 13240 4068 13252
rect 3844 13212 4068 13240
rect 3844 13200 3850 13212
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 5276 13240 5304 13348
rect 7377 13345 7389 13379
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 7644 13379 7702 13385
rect 7644 13345 7656 13379
rect 7690 13376 7702 13379
rect 9582 13376 9588 13388
rect 7690 13348 9588 13376
rect 7690 13345 7702 13348
rect 7644 13339 7702 13345
rect 9582 13336 9588 13348
rect 9640 13336 9646 13388
rect 12434 13376 12440 13388
rect 10428 13348 12440 13376
rect 5534 13308 5540 13320
rect 5495 13280 5540 13308
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13277 5687 13311
rect 6638 13308 6644 13320
rect 6599 13280 6644 13308
rect 5629 13271 5687 13277
rect 4172 13212 5304 13240
rect 3602 13132 3608 13184
rect 3660 13172 3666 13184
rect 4172 13172 4200 13212
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 5644 13240 5672 13271
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 7006 13308 7012 13320
rect 6871 13280 7012 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 10428 13308 10456 13348
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 12710 13376 12716 13388
rect 12671 13348 12716 13376
rect 12710 13336 12716 13348
rect 12768 13336 12774 13388
rect 12820 13376 12848 13407
rect 13078 13404 13084 13456
rect 13136 13444 13142 13456
rect 13909 13447 13967 13453
rect 13909 13444 13921 13447
rect 13136 13416 13921 13444
rect 13136 13404 13142 13416
rect 13909 13413 13921 13416
rect 13955 13413 13967 13447
rect 13909 13407 13967 13413
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15565 13447 15623 13453
rect 15565 13444 15577 13447
rect 15436 13416 15577 13444
rect 15436 13404 15442 13416
rect 15565 13413 15577 13416
rect 15611 13413 15623 13447
rect 16040 13444 16068 13484
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16298 13512 16304 13524
rect 16163 13484 16304 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16485 13515 16543 13521
rect 16485 13481 16497 13515
rect 16531 13512 16543 13515
rect 17494 13512 17500 13524
rect 16531 13484 17500 13512
rect 16531 13481 16543 13484
rect 16485 13475 16543 13481
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 17678 13472 17684 13524
rect 17736 13512 17742 13524
rect 18506 13512 18512 13524
rect 17736 13484 18175 13512
rect 18467 13484 18512 13512
rect 17736 13472 17742 13484
rect 18046 13444 18052 13456
rect 16040 13416 18052 13444
rect 15565 13407 15623 13413
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 13262 13376 13268 13388
rect 12820 13348 13268 13376
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13376 13875 13379
rect 14274 13376 14280 13388
rect 13863 13348 14280 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 14274 13336 14280 13348
rect 14332 13336 14338 13388
rect 14645 13379 14703 13385
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 15286 13376 15292 13388
rect 15247 13348 15292 13376
rect 14645 13339 14703 13345
rect 8628 13280 10456 13308
rect 8628 13268 8634 13280
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 10781 13311 10839 13317
rect 10781 13308 10793 13311
rect 10560 13280 10793 13308
rect 10560 13268 10566 13280
rect 10781 13277 10793 13280
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 11974 13308 11980 13320
rect 11931 13280 11980 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12308 13280 13001 13308
rect 12308 13268 12314 13280
rect 12989 13277 13001 13280
rect 13035 13308 13047 13311
rect 13446 13308 13452 13320
rect 13035 13280 13452 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 13630 13308 13636 13320
rect 13556 13280 13636 13308
rect 5408 13212 5672 13240
rect 5408 13200 5414 13212
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 12802 13240 12808 13252
rect 12584 13212 12808 13240
rect 12584 13200 12590 13212
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 3660 13144 4200 13172
rect 3660 13132 3666 13144
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8757 13175 8815 13181
rect 8757 13172 8769 13175
rect 8076 13144 8769 13172
rect 8076 13132 8082 13144
rect 8757 13141 8769 13144
rect 8803 13141 8815 13175
rect 8757 13135 8815 13141
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 13354 13172 13360 13184
rect 12391 13144 13360 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13449 13175 13507 13181
rect 13449 13141 13461 13175
rect 13495 13172 13507 13175
rect 13556 13172 13584 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13998 13308 14004 13320
rect 13959 13280 14004 13308
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 14660 13308 14688 13339
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15930 13336 15936 13388
rect 15988 13376 15994 13388
rect 16114 13376 16120 13388
rect 15988 13348 16120 13376
rect 15988 13336 15994 13348
rect 16114 13336 16120 13348
rect 16172 13376 16178 13388
rect 16172 13348 16436 13376
rect 16172 13336 16178 13348
rect 16206 13308 16212 13320
rect 14660 13280 16212 13308
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16408 13308 16436 13348
rect 16482 13336 16488 13388
rect 16540 13376 16546 13388
rect 17129 13379 17187 13385
rect 16540 13348 16712 13376
rect 16540 13336 16546 13348
rect 16684 13317 16712 13348
rect 17129 13345 17141 13379
rect 17175 13376 17187 13379
rect 17218 13376 17224 13388
rect 17175 13348 17224 13376
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 17396 13379 17454 13385
rect 17396 13345 17408 13379
rect 17442 13376 17454 13379
rect 17678 13376 17684 13388
rect 17442 13348 17684 13376
rect 17442 13345 17454 13348
rect 17396 13339 17454 13345
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 16577 13311 16635 13317
rect 16577 13308 16589 13311
rect 16408 13280 16589 13308
rect 16577 13277 16589 13280
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 16669 13311 16727 13317
rect 16669 13277 16681 13311
rect 16715 13277 16727 13311
rect 18147 13308 18175 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 18782 13512 18788 13524
rect 18743 13484 18788 13512
rect 18782 13472 18788 13484
rect 18840 13472 18846 13524
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 20254 13512 20260 13524
rect 18932 13484 19472 13512
rect 20215 13484 20260 13512
rect 18932 13472 18938 13484
rect 18524 13444 18552 13472
rect 18524 13416 19288 13444
rect 18414 13336 18420 13388
rect 18472 13376 18478 13388
rect 19153 13379 19211 13385
rect 19153 13376 19165 13379
rect 18472 13348 19165 13376
rect 18472 13336 18478 13348
rect 19153 13345 19165 13348
rect 19199 13345 19211 13379
rect 19260 13376 19288 13416
rect 19260 13348 19380 13376
rect 19153 13339 19211 13345
rect 19352 13317 19380 13348
rect 19444 13320 19472 13484
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 20162 13376 20168 13388
rect 20123 13348 20168 13376
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 18147 13280 19257 13308
rect 16669 13271 16727 13277
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19337 13311 19395 13317
rect 19337 13277 19349 13311
rect 19383 13277 19395 13311
rect 19337 13271 19395 13277
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13277 20407 13311
rect 20349 13271 20407 13277
rect 17034 13240 17040 13252
rect 13648 13212 17040 13240
rect 13648 13184 13676 13212
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 18782 13200 18788 13252
rect 18840 13240 18846 13252
rect 20364 13240 20392 13271
rect 18840 13212 20392 13240
rect 18840 13200 18846 13212
rect 13495 13144 13584 13172
rect 13495 13141 13507 13144
rect 13449 13135 13507 13141
rect 13630 13132 13636 13184
rect 13688 13132 13694 13184
rect 14829 13175 14887 13181
rect 14829 13141 14841 13175
rect 14875 13172 14887 13175
rect 18598 13172 18604 13184
rect 14875 13144 18604 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19797 13175 19855 13181
rect 19797 13172 19809 13175
rect 18932 13144 19809 13172
rect 18932 13132 18938 13144
rect 19797 13141 19809 13144
rect 19843 13141 19855 13175
rect 19797 13135 19855 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 3878 12968 3884 12980
rect 3839 12940 3884 12968
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4798 12968 4804 12980
rect 4212 12940 4804 12968
rect 4212 12928 4218 12940
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 8570 12968 8576 12980
rect 6696 12940 8576 12968
rect 6696 12928 6702 12940
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 9674 12968 9680 12980
rect 8680 12940 9680 12968
rect 1857 12903 1915 12909
rect 1857 12869 1869 12903
rect 1903 12900 1915 12903
rect 4338 12900 4344 12912
rect 1903 12872 4344 12900
rect 1903 12869 1915 12872
rect 1857 12863 1915 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 3292 12804 3433 12832
rect 3292 12792 3298 12804
rect 3421 12801 3433 12804
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 4430 12792 4436 12844
rect 4488 12832 4494 12844
rect 4525 12835 4583 12841
rect 4525 12832 4537 12835
rect 4488 12804 4537 12832
rect 4488 12792 4494 12804
rect 4525 12801 4537 12804
rect 4571 12832 4583 12835
rect 5350 12832 5356 12844
rect 4571 12804 5356 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 5350 12792 5356 12804
rect 5408 12832 5414 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5408 12804 5549 12832
rect 5408 12792 5414 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7248 12804 7941 12832
rect 7248 12792 7254 12804
rect 7929 12801 7941 12804
rect 7975 12832 7987 12835
rect 8018 12832 8024 12844
rect 7975 12804 8024 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8680 12841 8708 12940
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 12299 12940 13829 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 13817 12931 13875 12937
rect 14001 12971 14059 12977
rect 14001 12937 14013 12971
rect 14047 12968 14059 12971
rect 14182 12968 14188 12980
rect 14047 12940 14188 12968
rect 14047 12937 14059 12940
rect 14001 12931 14059 12937
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14274 12928 14280 12980
rect 14332 12968 14338 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 14332 12940 15025 12968
rect 14332 12928 14338 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 15102 12928 15108 12980
rect 15160 12928 15166 12980
rect 17218 12968 17224 12980
rect 16316 12940 17224 12968
rect 10045 12903 10103 12909
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 11333 12903 11391 12909
rect 10091 12872 11284 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12801 8723 12835
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 8665 12795 8723 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12832 11023 12835
rect 11256 12832 11284 12872
rect 11333 12869 11345 12903
rect 11379 12900 11391 12903
rect 12710 12900 12716 12912
rect 11379 12872 12716 12900
rect 11379 12869 11391 12872
rect 11333 12863 11391 12869
rect 12710 12860 12716 12872
rect 12768 12860 12774 12912
rect 12894 12860 12900 12912
rect 12952 12900 12958 12912
rect 13078 12900 13084 12912
rect 12952 12872 13084 12900
rect 12952 12860 12958 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 15120 12900 15148 12928
rect 13556 12872 15148 12900
rect 11790 12832 11796 12844
rect 11011 12804 11100 12832
rect 11256 12804 11376 12832
rect 11751 12804 11796 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 2317 12767 2375 12773
rect 2317 12733 2329 12767
rect 2363 12764 2375 12767
rect 3878 12764 3884 12776
rect 2363 12736 3884 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 4246 12764 4252 12776
rect 4028 12736 4252 12764
rect 4028 12724 4034 12736
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 7742 12764 7748 12776
rect 7340 12736 7748 12764
rect 7340 12724 7346 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 10870 12764 10876 12776
rect 8404 12736 10876 12764
rect 3326 12696 3332 12708
rect 3239 12668 3332 12696
rect 3326 12656 3332 12668
rect 3384 12696 3390 12708
rect 3694 12696 3700 12708
rect 3384 12668 3700 12696
rect 3384 12656 3390 12668
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 4341 12699 4399 12705
rect 4341 12665 4353 12699
rect 4387 12696 4399 12699
rect 4798 12696 4804 12708
rect 4387 12668 4804 12696
rect 4387 12665 4399 12668
rect 4341 12659 4399 12665
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5350 12696 5356 12708
rect 4948 12668 5356 12696
rect 4948 12656 4954 12668
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 5445 12699 5503 12705
rect 5445 12665 5457 12699
rect 5491 12696 5503 12699
rect 8404 12696 8432 12736
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 5491 12668 8432 12696
rect 5491 12665 5503 12668
rect 5445 12659 5503 12665
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 8932 12699 8990 12705
rect 8932 12696 8944 12699
rect 8812 12668 8944 12696
rect 8812 12656 8818 12668
rect 8932 12665 8944 12668
rect 8978 12696 8990 12699
rect 11072 12696 11100 12804
rect 11348 12776 11376 12804
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12832 12035 12835
rect 12250 12832 12256 12844
rect 12023 12804 12256 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 11992 12764 12020 12795
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 13556 12841 13584 12872
rect 15378 12860 15384 12912
rect 15436 12900 15442 12912
rect 15654 12900 15660 12912
rect 15436 12872 15660 12900
rect 15436 12860 15442 12872
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12676 12804 13001 12832
rect 12676 12792 12682 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12832 14703 12835
rect 15010 12832 15016 12844
rect 14691 12804 15016 12832
rect 14691 12801 14703 12804
rect 14645 12795 14703 12801
rect 15010 12792 15016 12804
rect 15068 12832 15074 12844
rect 15565 12835 15623 12841
rect 15565 12832 15577 12835
rect 15068 12804 15577 12832
rect 15068 12792 15074 12804
rect 15565 12801 15577 12804
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 16316 12841 16344 12940
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 17678 12968 17684 12980
rect 17639 12940 17684 12968
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18049 12971 18107 12977
rect 18049 12968 18061 12971
rect 18012 12940 18061 12968
rect 18012 12928 18018 12940
rect 18049 12937 18061 12940
rect 18095 12937 18107 12971
rect 18049 12931 18107 12937
rect 18506 12928 18512 12980
rect 18564 12968 18570 12980
rect 19978 12968 19984 12980
rect 18564 12940 19984 12968
rect 18564 12928 18570 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 15896 12804 16313 12832
rect 15896 12792 15902 12804
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 17696 12832 17724 12928
rect 17773 12903 17831 12909
rect 17773 12869 17785 12903
rect 17819 12900 17831 12903
rect 18782 12900 18788 12912
rect 17819 12872 18788 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 18782 12860 18788 12872
rect 18840 12860 18846 12912
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 17696 12804 18613 12832
rect 16301 12795 16359 12801
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 12802 12764 12808 12776
rect 11388 12736 12020 12764
rect 12763 12736 12808 12764
rect 11388 12724 11394 12736
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 12894 12724 12900 12776
rect 12952 12764 12958 12776
rect 14369 12767 14427 12773
rect 12952 12736 12997 12764
rect 12952 12724 12958 12736
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 15194 12764 15200 12776
rect 14415 12736 15200 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 15194 12724 15200 12736
rect 15252 12764 15258 12776
rect 15378 12764 15384 12776
rect 15252 12736 15384 12764
rect 15252 12724 15258 12736
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12764 15531 12767
rect 16568 12767 16626 12773
rect 15519 12736 16344 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 16316 12708 16344 12736
rect 16568 12733 16580 12767
rect 16614 12764 16626 12767
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 16614 12736 17785 12764
rect 16614 12733 16626 12736
rect 16568 12727 16626 12733
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 17773 12727 17831 12733
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12764 18475 12767
rect 18874 12764 18880 12776
rect 18463 12736 18880 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 19426 12764 19432 12776
rect 19383 12736 19432 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 8978 12668 11100 12696
rect 8978 12665 8990 12668
rect 8932 12659 8990 12665
rect 2225 12631 2283 12637
rect 2225 12597 2237 12631
rect 2271 12628 2283 12631
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2271 12600 2881 12628
rect 2271 12597 2283 12600
rect 2225 12591 2283 12597
rect 2869 12597 2881 12600
rect 2915 12597 2927 12631
rect 2869 12591 2927 12597
rect 3237 12631 3295 12637
rect 3237 12597 3249 12631
rect 3283 12628 3295 12631
rect 5994 12628 6000 12640
rect 3283 12600 6000 12628
rect 3283 12597 3295 12600
rect 3237 12591 3295 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 7650 12628 7656 12640
rect 7611 12600 7656 12628
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 10318 12628 10324 12640
rect 10279 12600 10324 12628
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10686 12628 10692 12640
rect 10647 12600 10692 12628
rect 10686 12588 10692 12600
rect 10744 12628 10750 12640
rect 10870 12628 10876 12640
rect 10744 12600 10876 12628
rect 10744 12588 10750 12600
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 11072 12628 11100 12668
rect 11701 12699 11759 12705
rect 11701 12665 11713 12699
rect 11747 12696 11759 12699
rect 12342 12696 12348 12708
rect 11747 12668 12348 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 12342 12656 12348 12668
rect 12400 12656 12406 12708
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 14461 12699 14519 12705
rect 14461 12696 14473 12699
rect 13964 12668 14473 12696
rect 13964 12656 13970 12668
rect 14461 12665 14473 12668
rect 14507 12665 14519 12699
rect 14461 12659 14519 12665
rect 14568 12668 15700 12696
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11072 12600 12265 12628
rect 12253 12597 12265 12600
rect 12299 12597 12311 12631
rect 12253 12591 12311 12597
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 13630 12628 13636 12640
rect 12483 12600 13636 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 14568 12628 14596 12668
rect 15378 12628 15384 12640
rect 13863 12600 14596 12628
rect 15339 12600 15384 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 15672 12628 15700 12668
rect 16298 12656 16304 12708
rect 16356 12656 16362 12708
rect 17954 12656 17960 12708
rect 18012 12696 18018 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 18012 12668 18521 12696
rect 18012 12656 18018 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 19604 12699 19662 12705
rect 19604 12665 19616 12699
rect 19650 12696 19662 12699
rect 20070 12696 20076 12708
rect 19650 12668 20076 12696
rect 19650 12665 19662 12668
rect 19604 12659 19662 12665
rect 20070 12656 20076 12668
rect 20128 12656 20134 12708
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 15672 12600 20729 12628
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2961 12427 3019 12433
rect 2961 12424 2973 12427
rect 2096 12396 2973 12424
rect 2096 12384 2102 12396
rect 2961 12393 2973 12396
rect 3007 12393 3019 12427
rect 2961 12387 3019 12393
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4433 12427 4491 12433
rect 4433 12424 4445 12427
rect 4396 12396 4445 12424
rect 4396 12384 4402 12396
rect 4433 12393 4445 12396
rect 4479 12393 4491 12427
rect 4433 12387 4491 12393
rect 5350 12384 5356 12436
rect 5408 12424 5414 12436
rect 5534 12424 5540 12436
rect 5408 12396 5540 12424
rect 5408 12384 5414 12396
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 5629 12427 5687 12433
rect 5629 12393 5641 12427
rect 5675 12424 5687 12427
rect 5902 12424 5908 12436
rect 5675 12396 5908 12424
rect 5675 12393 5687 12396
rect 5629 12387 5687 12393
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 7708 12396 8401 12424
rect 7708 12384 7714 12396
rect 8389 12393 8401 12396
rect 8435 12393 8447 12427
rect 8389 12387 8447 12393
rect 10045 12427 10103 12433
rect 10045 12393 10057 12427
rect 10091 12424 10103 12427
rect 10318 12424 10324 12436
rect 10091 12396 10324 12424
rect 10091 12393 10103 12396
rect 10045 12387 10103 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10962 12424 10968 12436
rect 10744 12396 10968 12424
rect 10744 12384 10750 12396
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12860 12396 12909 12424
rect 12860 12384 12866 12396
rect 12897 12393 12909 12396
rect 12943 12393 12955 12427
rect 13354 12424 13360 12436
rect 13315 12396 13360 12424
rect 12897 12387 12955 12393
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12393 13967 12427
rect 13909 12387 13967 12393
rect 17129 12427 17187 12433
rect 17129 12393 17141 12427
rect 17175 12393 17187 12427
rect 18782 12424 18788 12436
rect 18743 12396 18788 12424
rect 17129 12387 17187 12393
rect 3510 12356 3516 12368
rect 3471 12328 3516 12356
rect 3510 12316 3516 12328
rect 3568 12316 3574 12368
rect 5997 12359 6055 12365
rect 5997 12325 6009 12359
rect 6043 12356 6055 12359
rect 6448 12359 6506 12365
rect 6448 12356 6460 12359
rect 6043 12328 6460 12356
rect 6043 12325 6055 12328
rect 5997 12319 6055 12325
rect 6448 12325 6460 12328
rect 6494 12356 6506 12359
rect 7190 12356 7196 12368
rect 6494 12328 7196 12356
rect 6494 12325 6506 12328
rect 6448 12319 6506 12325
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 7742 12316 7748 12368
rect 7800 12356 7806 12368
rect 8481 12359 8539 12365
rect 8481 12356 8493 12359
rect 7800 12328 8493 12356
rect 7800 12316 7806 12328
rect 8481 12325 8493 12328
rect 8527 12325 8539 12359
rect 8481 12319 8539 12325
rect 8662 12316 8668 12368
rect 8720 12356 8726 12368
rect 12066 12356 12072 12368
rect 8720 12328 12072 12356
rect 8720 12316 8726 12328
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 13265 12359 13323 12365
rect 13265 12325 13277 12359
rect 13311 12356 13323 12359
rect 13924 12356 13952 12387
rect 13311 12328 13952 12356
rect 17144 12356 17172 12387
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 19610 12424 19616 12436
rect 19567 12396 19616 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 20162 12384 20168 12436
rect 20220 12384 20226 12436
rect 17672 12359 17730 12365
rect 17672 12356 17684 12359
rect 17144 12328 17684 12356
rect 13311 12325 13323 12328
rect 13265 12319 13323 12325
rect 17672 12325 17684 12328
rect 17718 12356 17730 12359
rect 17862 12356 17868 12368
rect 17718 12328 17868 12356
rect 17718 12325 17730 12328
rect 17672 12319 17730 12325
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 19061 12359 19119 12365
rect 19061 12325 19073 12359
rect 19107 12356 19119 12359
rect 20180 12356 20208 12384
rect 19107 12328 20208 12356
rect 19107 12325 19119 12328
rect 19061 12319 19119 12325
rect 1848 12291 1906 12297
rect 1848 12257 1860 12291
rect 1894 12288 1906 12291
rect 2590 12288 2596 12300
rect 1894 12260 2596 12288
rect 1894 12257 1906 12260
rect 1848 12251 1906 12257
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12288 3295 12291
rect 3283 12260 3556 12288
rect 3283 12257 3295 12260
rect 3237 12251 3295 12257
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 3528 12152 3556 12260
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 5074 12288 5080 12300
rect 4304 12260 5080 12288
rect 4304 12248 4310 12260
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5258 12248 5264 12300
rect 5316 12288 5322 12300
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 5316 12260 5549 12288
rect 5316 12248 5322 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 6181 12291 6239 12297
rect 6181 12288 6193 12291
rect 5960 12260 6193 12288
rect 5960 12248 5966 12260
rect 6181 12257 6193 12260
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 10962 12288 10968 12300
rect 9263 12260 10968 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 11146 12248 11152 12300
rect 11204 12288 11210 12300
rect 11241 12291 11299 12297
rect 11241 12288 11253 12291
rect 11204 12260 11253 12288
rect 11204 12248 11210 12260
rect 11241 12257 11253 12260
rect 11287 12257 11299 12291
rect 11241 12251 11299 12257
rect 11330 12248 11336 12300
rect 11388 12248 11394 12300
rect 11508 12291 11566 12297
rect 11508 12257 11520 12291
rect 11554 12288 11566 12291
rect 11790 12288 11796 12300
rect 11554 12260 11796 12288
rect 11554 12257 11566 12260
rect 11508 12251 11566 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 14274 12288 14280 12300
rect 14235 12260 14280 12288
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 15838 12288 15844 12300
rect 15795 12260 15844 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 16022 12297 16028 12300
rect 16016 12251 16028 12297
rect 16080 12288 16086 12300
rect 16080 12260 16116 12288
rect 16022 12248 16028 12251
rect 16080 12248 16086 12260
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 17405 12291 17463 12297
rect 17405 12288 17417 12291
rect 17276 12260 17417 12288
rect 17276 12248 17282 12260
rect 17405 12257 17417 12260
rect 17451 12257 17463 12291
rect 17405 12251 17463 12257
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 19760 12260 19901 12288
rect 19760 12248 19766 12260
rect 19889 12257 19901 12260
rect 19935 12257 19947 12291
rect 19889 12251 19947 12257
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4430 12220 4436 12232
rect 3752 12192 4436 12220
rect 3752 12180 3758 12192
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4706 12220 4712 12232
rect 4667 12192 4712 12220
rect 4525 12183 4583 12189
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 3528 12124 4077 12152
rect 4065 12121 4077 12124
rect 4111 12121 4123 12155
rect 4540 12152 4568 12183
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12220 5871 12223
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5859 12192 6009 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12220 8723 12223
rect 8754 12220 8760 12232
rect 8711 12192 8760 12220
rect 8711 12189 8723 12192
rect 8665 12183 8723 12189
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10502 12220 10508 12232
rect 10367 12192 10508 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 6086 12152 6092 12164
rect 4540 12124 6092 12152
rect 4065 12115 4123 12121
rect 6086 12112 6092 12124
rect 6144 12112 6150 12164
rect 8021 12155 8079 12161
rect 8021 12121 8033 12155
rect 8067 12152 8079 12155
rect 10152 12152 10180 12183
rect 10502 12180 10508 12192
rect 10560 12220 10566 12232
rect 11348 12220 11376 12248
rect 10560 12192 11376 12220
rect 10560 12180 10566 12192
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13412 12192 13461 12220
rect 13412 12180 13418 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 14366 12220 14372 12232
rect 14279 12192 14372 12220
rect 13449 12183 13507 12189
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 8067 12124 10180 12152
rect 8067 12121 8079 12124
rect 8021 12115 8079 12121
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 14384 12152 14412 12180
rect 12584 12124 14412 12152
rect 12584 12112 12590 12124
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 3844 12056 5181 12084
rect 3844 12044 3850 12056
rect 5169 12053 5181 12056
rect 5215 12053 5227 12087
rect 7558 12084 7564 12096
rect 7519 12056 7564 12084
rect 5169 12047 5227 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8478 12084 8484 12096
rect 8352 12056 8484 12084
rect 8352 12044 8358 12056
rect 8478 12044 8484 12056
rect 8536 12084 8542 12096
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 8536 12056 9045 12084
rect 8536 12044 8542 12056
rect 9033 12053 9045 12056
rect 9079 12053 9091 12087
rect 9033 12047 9091 12053
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 12894 12084 12900 12096
rect 9723 12056 12900 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 14476 12084 14504 12183
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19981 12223 20039 12229
rect 19981 12220 19993 12223
rect 19484 12192 19993 12220
rect 19484 12180 19490 12192
rect 19981 12189 19993 12192
rect 20027 12189 20039 12223
rect 20162 12220 20168 12232
rect 20123 12192 20168 12220
rect 19981 12183 20039 12189
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 19886 12152 19892 12164
rect 19024 12124 19892 12152
rect 19024 12112 19030 12124
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 13504 12056 14504 12084
rect 13504 12044 13510 12056
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11880 1823 11883
rect 2314 11880 2320 11892
rect 1811 11852 2320 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11880 3387 11883
rect 12437 11883 12495 11889
rect 3375 11852 9168 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 3234 11772 3240 11824
rect 3292 11812 3298 11824
rect 4249 11815 4307 11821
rect 4249 11812 4261 11815
rect 3292 11784 4261 11812
rect 3292 11772 3298 11784
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2317 11747 2375 11753
rect 2317 11744 2329 11747
rect 2096 11716 2329 11744
rect 2096 11704 2102 11716
rect 2317 11713 2329 11716
rect 2363 11713 2375 11747
rect 3786 11744 3792 11756
rect 3747 11716 3792 11744
rect 2317 11707 2375 11713
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 3896 11753 3924 11784
rect 4249 11781 4261 11784
rect 4295 11781 4307 11815
rect 5718 11812 5724 11824
rect 5679 11784 5724 11812
rect 4249 11775 4307 11781
rect 5718 11772 5724 11784
rect 5776 11772 5782 11824
rect 6086 11772 6092 11824
rect 6144 11812 6150 11824
rect 8849 11815 8907 11821
rect 8849 11812 8861 11815
rect 6144 11784 8861 11812
rect 6144 11772 6150 11784
rect 8849 11781 8861 11784
rect 8895 11781 8907 11815
rect 8849 11775 8907 11781
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11713 3939 11747
rect 5994 11744 6000 11756
rect 5955 11716 6000 11744
rect 3881 11707 3939 11713
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 6104 11716 7389 11744
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 4080 11648 4353 11676
rect 1946 11568 1952 11620
rect 2004 11608 2010 11620
rect 2133 11611 2191 11617
rect 2133 11608 2145 11611
rect 2004 11580 2145 11608
rect 2004 11568 2010 11580
rect 2133 11577 2145 11580
rect 2179 11577 2191 11611
rect 2133 11571 2191 11577
rect 3602 11568 3608 11620
rect 3660 11608 3666 11620
rect 3697 11611 3755 11617
rect 3697 11608 3709 11611
rect 3660 11580 3709 11608
rect 3660 11568 3666 11580
rect 3697 11577 3709 11580
rect 3743 11608 3755 11611
rect 3970 11608 3976 11620
rect 3743 11580 3976 11608
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 3970 11568 3976 11580
rect 4028 11568 4034 11620
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 3786 11500 3792 11552
rect 3844 11540 3850 11552
rect 4080 11540 4108 11648
rect 4341 11645 4353 11648
rect 4387 11676 4399 11679
rect 5902 11676 5908 11688
rect 4387 11648 5908 11676
rect 4387 11645 4399 11648
rect 4341 11639 4399 11645
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 4249 11611 4307 11617
rect 4249 11577 4261 11611
rect 4295 11608 4307 11611
rect 4586 11611 4644 11617
rect 4586 11608 4598 11611
rect 4295 11580 4598 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 4586 11577 4598 11580
rect 4632 11608 4644 11611
rect 6104 11608 6132 11716
rect 7377 11713 7389 11716
rect 7423 11744 7435 11747
rect 7558 11744 7564 11756
rect 7423 11716 7564 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 8389 11747 8447 11753
rect 8389 11744 8401 11747
rect 8260 11716 8401 11744
rect 8260 11704 8266 11716
rect 8389 11713 8401 11716
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 4632 11580 6132 11608
rect 7193 11611 7251 11617
rect 4632 11577 4644 11580
rect 4586 11571 4644 11577
rect 7193 11577 7205 11611
rect 7239 11608 7251 11611
rect 7239 11580 7420 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 6822 11540 6828 11552
rect 3844 11512 4108 11540
rect 6783 11512 6828 11540
rect 3844 11500 3850 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7285 11543 7343 11549
rect 7285 11540 7297 11543
rect 7156 11512 7297 11540
rect 7156 11500 7162 11512
rect 7285 11509 7297 11512
rect 7331 11509 7343 11543
rect 7392 11540 7420 11580
rect 7837 11543 7895 11549
rect 7837 11540 7849 11543
rect 7392 11512 7849 11540
rect 7285 11503 7343 11509
rect 7837 11509 7849 11512
rect 7883 11509 7895 11543
rect 8202 11540 8208 11552
rect 8163 11512 8208 11540
rect 7837 11503 7895 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8297 11543 8355 11549
rect 8297 11509 8309 11543
rect 8343 11540 8355 11543
rect 9030 11540 9036 11552
rect 8343 11512 9036 11540
rect 8343 11509 8355 11512
rect 8297 11503 8355 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9140 11540 9168 11852
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12802 11880 12808 11892
rect 12483 11852 12808 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 16022 11880 16028 11892
rect 15983 11852 16028 11880
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 17589 11883 17647 11889
rect 17589 11849 17601 11883
rect 17635 11880 17647 11883
rect 17770 11880 17776 11892
rect 17635 11852 17776 11880
rect 17635 11849 17647 11852
rect 17589 11843 17647 11849
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18049 11883 18107 11889
rect 18049 11880 18061 11883
rect 18012 11852 18061 11880
rect 18012 11840 18018 11852
rect 18049 11849 18061 11852
rect 18095 11849 18107 11883
rect 18049 11843 18107 11849
rect 20162 11840 20168 11892
rect 20220 11880 20226 11892
rect 20533 11883 20591 11889
rect 20533 11880 20545 11883
rect 20220 11852 20545 11880
rect 20220 11840 20226 11852
rect 20533 11849 20545 11852
rect 20579 11849 20591 11883
rect 20990 11880 20996 11892
rect 20951 11852 20996 11880
rect 20533 11843 20591 11849
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 11333 11815 11391 11821
rect 11333 11781 11345 11815
rect 11379 11812 11391 11815
rect 11790 11812 11796 11824
rect 11379 11784 11796 11812
rect 11379 11781 11391 11784
rect 11333 11775 11391 11781
rect 11790 11772 11796 11784
rect 11848 11812 11854 11824
rect 11848 11784 13124 11812
rect 11848 11772 11854 11784
rect 9398 11744 9404 11756
rect 9359 11716 9404 11744
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9950 11744 9956 11756
rect 9732 11716 9956 11744
rect 9732 11704 9738 11716
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 12894 11744 12900 11756
rect 12855 11716 12900 11744
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 13096 11753 13124 11784
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13354 11744 13360 11756
rect 13127 11716 13360 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 14274 11744 14280 11756
rect 13495 11716 14280 11744
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 16040 11744 16068 11840
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16040 11716 16865 11744
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11744 18659 11747
rect 18782 11744 18788 11756
rect 18647 11716 18788 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 10220 11679 10278 11685
rect 10220 11645 10232 11679
rect 10266 11676 10278 11679
rect 10502 11676 10508 11688
rect 10266 11648 10508 11676
rect 10266 11645 10278 11648
rect 10220 11639 10278 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 11020 11648 12265 11676
rect 11020 11636 11026 11648
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12768 11648 12817 11676
rect 12768 11636 12774 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14608 11648 14657 11676
rect 14608 11636 14614 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 14912 11679 14970 11685
rect 14912 11645 14924 11679
rect 14958 11676 14970 11679
rect 15654 11676 15660 11688
rect 14958 11648 15660 11676
rect 14958 11645 14970 11648
rect 14912 11639 14970 11645
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 17126 11636 17132 11688
rect 17184 11676 17190 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 17184 11648 17417 11676
rect 17184 11636 17190 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11676 18567 11679
rect 18690 11676 18696 11688
rect 18555 11648 18696 11676
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 19116 11648 19165 11676
rect 19116 11636 19122 11648
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 20806 11676 20812 11688
rect 20767 11648 20812 11676
rect 19153 11639 19211 11645
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 9306 11608 9312 11620
rect 9267 11580 9312 11608
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 9490 11568 9496 11620
rect 9548 11608 9554 11620
rect 15102 11608 15108 11620
rect 9548 11580 15108 11608
rect 9548 11568 9554 11580
rect 15102 11568 15108 11580
rect 15160 11568 15166 11620
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 16761 11611 16819 11617
rect 16761 11608 16773 11611
rect 15344 11580 16773 11608
rect 15344 11568 15350 11580
rect 16761 11577 16773 11580
rect 16807 11577 16819 11611
rect 16761 11571 16819 11577
rect 19420 11611 19478 11617
rect 19420 11577 19432 11611
rect 19466 11608 19478 11611
rect 19886 11608 19892 11620
rect 19466 11580 19892 11608
rect 19466 11577 19478 11580
rect 19420 11571 19478 11577
rect 19886 11568 19892 11580
rect 19944 11568 19950 11620
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 9140 11512 9229 11540
rect 9217 11509 9229 11512
rect 9263 11509 9275 11543
rect 9217 11503 9275 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10778 11540 10784 11552
rect 9456 11512 10784 11540
rect 9456 11500 9462 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 12069 11543 12127 11549
rect 12069 11509 12081 11543
rect 12115 11540 12127 11543
rect 13170 11540 13176 11552
rect 12115 11512 13176 11540
rect 12115 11509 12127 11512
rect 12069 11503 12127 11509
rect 13170 11500 13176 11512
rect 13228 11540 13234 11552
rect 13722 11540 13728 11552
rect 13228 11512 13728 11540
rect 13228 11500 13234 11512
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 15436 11512 16313 11540
rect 15436 11500 15442 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16666 11540 16672 11552
rect 16627 11512 16672 11540
rect 16301 11503 16359 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 18414 11540 18420 11552
rect 18375 11512 18420 11540
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2222 11336 2228 11348
rect 1995 11308 2228 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2363 11308 2973 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 2961 11299 3019 11305
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 4246 11336 4252 11348
rect 3467 11308 4252 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4764 11308 5457 11336
rect 4764 11296 4770 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5445 11299 5503 11305
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 8662 11336 8668 11348
rect 6604 11308 8524 11336
rect 8623 11308 8668 11336
rect 6604 11296 6610 11308
rect 2498 11228 2504 11280
rect 2556 11268 2562 11280
rect 4332 11271 4390 11277
rect 4332 11268 4344 11271
rect 2556 11240 4344 11268
rect 2556 11228 2562 11240
rect 4332 11237 4344 11240
rect 4378 11268 4390 11271
rect 5718 11268 5724 11280
rect 4378 11240 5724 11268
rect 4378 11237 4390 11240
rect 4332 11231 4390 11237
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 8294 11268 8300 11280
rect 6564 11240 8300 11268
rect 6564 11209 6592 11240
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 6914 11209 6920 11212
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3375 11172 3893 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 6908 11163 6920 11209
rect 6972 11200 6978 11212
rect 8496 11200 8524 11308
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 10594 11336 10600 11348
rect 8904 11308 10600 11336
rect 8904 11296 8910 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 11020 11308 11805 11336
rect 11020 11296 11026 11308
rect 11793 11305 11805 11308
rect 11839 11305 11851 11339
rect 11793 11299 11851 11305
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 14366 11336 14372 11348
rect 13688 11308 14372 11336
rect 13688 11296 13694 11308
rect 14366 11296 14372 11308
rect 14424 11336 14430 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 14424 11308 14565 11336
rect 14424 11296 14430 11308
rect 14553 11305 14565 11308
rect 14599 11305 14611 11339
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 14553 11299 14611 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 15703 11308 16313 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16632 11308 16681 11336
rect 16632 11296 16638 11308
rect 16669 11305 16681 11308
rect 16715 11336 16727 11339
rect 16942 11336 16948 11348
rect 16715 11308 16948 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17770 11336 17776 11348
rect 17731 11308 17776 11336
rect 17770 11296 17776 11308
rect 17828 11336 17834 11348
rect 19242 11336 19248 11348
rect 17828 11308 19248 11336
rect 17828 11296 17834 11308
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19702 11336 19708 11348
rect 19663 11308 19708 11336
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 11698 11268 11704 11280
rect 8803 11240 11704 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 12618 11277 12624 11280
rect 12612 11268 12624 11277
rect 12579 11240 12624 11268
rect 12612 11231 12624 11240
rect 12618 11228 12624 11231
rect 12676 11228 12682 11280
rect 14090 11228 14096 11280
rect 14148 11268 14154 11280
rect 14645 11271 14703 11277
rect 14645 11268 14657 11271
rect 14148 11240 14657 11268
rect 14148 11228 14154 11240
rect 14645 11237 14657 11240
rect 14691 11237 14703 11271
rect 14645 11231 14703 11237
rect 16114 11228 16120 11280
rect 16172 11268 16178 11280
rect 16761 11271 16819 11277
rect 16761 11268 16773 11271
rect 16172 11240 16773 11268
rect 16172 11228 16178 11240
rect 16761 11237 16773 11240
rect 16807 11237 16819 11271
rect 16761 11231 16819 11237
rect 17681 11271 17739 11277
rect 17681 11237 17693 11271
rect 17727 11268 17739 11271
rect 20162 11268 20168 11280
rect 17727 11240 20168 11268
rect 17727 11237 17739 11240
rect 17681 11231 17739 11237
rect 20162 11228 20168 11240
rect 20220 11228 20226 11280
rect 6972 11172 7008 11200
rect 8496 11172 9076 11200
rect 6914 11160 6920 11163
rect 6972 11160 6978 11172
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2280 11104 2421 11132
rect 2280 11092 2286 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2590 11132 2596 11144
rect 2551 11104 2596 11132
rect 2409 11095 2467 11101
rect 2590 11092 2596 11104
rect 2648 11092 2654 11144
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11132 3663 11135
rect 3694 11132 3700 11144
rect 3651 11104 3700 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 3694 11092 3700 11104
rect 3752 11092 3758 11144
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 3510 11064 3516 11076
rect 2188 11036 3516 11064
rect 2188 11024 2194 11036
rect 3510 11024 3516 11036
rect 3568 11064 3574 11076
rect 3786 11064 3792 11076
rect 3568 11036 3792 11064
rect 3568 11024 3574 11036
rect 3786 11024 3792 11036
rect 3844 11064 3850 11076
rect 4080 11064 4108 11095
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 5960 11104 6653 11132
rect 5960 11092 5966 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11101 8907 11135
rect 9048 11132 9076 11172
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 9180 11172 10517 11200
rect 9180 11160 9186 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11200 12403 11203
rect 12434 11200 12440 11212
rect 12391 11172 12440 11200
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 15252 11172 18000 11200
rect 15252 11160 15258 11172
rect 9048 11104 9536 11132
rect 8849 11095 8907 11101
rect 6362 11064 6368 11076
rect 3844 11036 4108 11064
rect 6323 11036 6368 11064
rect 3844 11024 3850 11036
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8478 11064 8484 11076
rect 8067 11036 8484 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 8478 11024 8484 11036
rect 8536 11064 8542 11076
rect 8864 11064 8892 11095
rect 9398 11064 9404 11076
rect 8536 11036 9404 11064
rect 8536 11024 8542 11036
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 3881 10999 3939 11005
rect 3881 10965 3893 10999
rect 3927 10996 3939 10999
rect 4798 10996 4804 11008
rect 3927 10968 4804 10996
rect 3927 10965 3939 10968
rect 3881 10959 3939 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 8294 10996 8300 11008
rect 8255 10968 8300 10996
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 9508 10996 9536 11104
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 12250 11132 12256 11144
rect 9640 11104 12256 11132
rect 9640 11092 9646 11104
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11132 14887 11135
rect 14918 11132 14924 11144
rect 14875 11104 14924 11132
rect 14875 11101 14887 11104
rect 14829 11095 14887 11101
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15028 11104 15761 11132
rect 14185 11067 14243 11073
rect 14185 11033 14197 11067
rect 14231 11064 14243 11067
rect 15028 11064 15056 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11132 17003 11135
rect 17770 11132 17776 11144
rect 16991 11104 17776 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 14231 11036 15056 11064
rect 14231 11033 14243 11036
rect 14185 11027 14243 11033
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 15856 11064 15884 11095
rect 16206 11064 16212 11076
rect 15712 11036 16212 11064
rect 15712 11024 15718 11036
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 16758 11024 16764 11076
rect 16816 11064 16822 11076
rect 16960 11064 16988 11095
rect 17770 11092 17776 11104
rect 17828 11132 17834 11144
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 17828 11104 17877 11132
rect 17828 11092 17834 11104
rect 17865 11101 17877 11104
rect 17911 11101 17923 11135
rect 17972 11132 18000 11172
rect 18598 11160 18604 11212
rect 18656 11200 18662 11212
rect 18693 11203 18751 11209
rect 18693 11200 18705 11203
rect 18656 11172 18705 11200
rect 18656 11160 18662 11172
rect 18693 11169 18705 11172
rect 18739 11169 18751 11203
rect 20070 11200 20076 11212
rect 20031 11172 20076 11200
rect 18693 11163 18751 11169
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 17972 11104 18797 11132
rect 17865 11095 17923 11101
rect 18785 11101 18797 11104
rect 18831 11101 18843 11135
rect 18785 11095 18843 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 16816 11036 16988 11064
rect 17880 11064 17908 11095
rect 18892 11064 18920 11095
rect 19978 11092 19984 11144
rect 20036 11132 20042 11144
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 20036 11104 20177 11132
rect 20036 11092 20042 11104
rect 20165 11101 20177 11104
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 20257 11135 20315 11141
rect 20257 11101 20269 11135
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 17880 11036 18920 11064
rect 16816 11024 16822 11036
rect 19886 11024 19892 11076
rect 19944 11064 19950 11076
rect 20272 11064 20300 11095
rect 19944 11036 20300 11064
rect 19944 11024 19950 11036
rect 11146 10996 11152 11008
rect 9508 10968 11152 10996
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 13725 10999 13783 11005
rect 13725 10996 13737 10999
rect 13596 10968 13737 10996
rect 13596 10956 13602 10968
rect 13725 10965 13737 10968
rect 13771 10965 13783 10999
rect 16224 10996 16252 11024
rect 16850 10996 16856 11008
rect 16224 10968 16856 10996
rect 13725 10959 13783 10965
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17313 10999 17371 11005
rect 17313 10996 17325 10999
rect 17000 10968 17325 10996
rect 17000 10956 17006 10968
rect 17313 10965 17325 10968
rect 17359 10965 17371 10999
rect 17313 10959 17371 10965
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18325 10999 18383 11005
rect 18325 10996 18337 10999
rect 18012 10968 18337 10996
rect 18012 10956 18018 10968
rect 18325 10965 18337 10968
rect 18371 10965 18383 10999
rect 18325 10959 18383 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 3878 10792 3884 10804
rect 3839 10764 3884 10792
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 10962 10792 10968 10804
rect 4120 10764 10968 10792
rect 4120 10752 4126 10764
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 15746 10792 15752 10804
rect 14844 10764 15752 10792
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 4985 10727 5043 10733
rect 4985 10724 4997 10727
rect 4672 10696 4997 10724
rect 4672 10684 4678 10696
rect 4985 10693 4997 10696
rect 5031 10693 5043 10727
rect 4985 10687 5043 10693
rect 8021 10727 8079 10733
rect 8021 10693 8033 10727
rect 8067 10724 8079 10727
rect 9582 10724 9588 10736
rect 8067 10696 9588 10724
rect 8067 10693 8079 10696
rect 8021 10687 8079 10693
rect 9582 10684 9588 10696
rect 9640 10684 9646 10736
rect 11057 10727 11115 10733
rect 11057 10693 11069 10727
rect 11103 10724 11115 10727
rect 11606 10724 11612 10736
rect 11103 10696 11612 10724
rect 11103 10693 11115 10696
rect 11057 10687 11115 10693
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 2130 10656 2136 10668
rect 1636 10628 2136 10656
rect 1636 10616 1642 10628
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 3292 10628 4445 10656
rect 3292 10616 3298 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5960 10628 6285 10656
rect 5960 10616 5966 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 7558 10656 7564 10668
rect 7519 10628 7564 10656
rect 6273 10619 6331 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8846 10656 8852 10668
rect 8711 10628 8852 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9398 10656 9404 10668
rect 9359 10628 9404 10656
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11072 10628 11713 10656
rect 2866 10548 2872 10600
rect 2924 10588 2930 10600
rect 3142 10588 3148 10600
rect 2924 10560 3148 10588
rect 2924 10548 2930 10560
rect 3142 10548 3148 10560
rect 3200 10588 3206 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 3200 10560 4353 10588
rect 3200 10548 3206 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 5169 10591 5227 10597
rect 5169 10557 5181 10591
rect 5215 10588 5227 10591
rect 6362 10588 6368 10600
rect 5215 10560 6368 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 8386 10588 8392 10600
rect 8347 10560 8392 10588
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8956 10588 8984 10616
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8527 10560 9321 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 2400 10523 2458 10529
rect 2400 10489 2412 10523
rect 2446 10520 2458 10523
rect 3694 10520 3700 10532
rect 2446 10492 3700 10520
rect 2446 10489 2458 10492
rect 2400 10483 2458 10489
rect 3694 10480 3700 10492
rect 3752 10480 3758 10532
rect 5810 10480 5816 10532
rect 5868 10520 5874 10532
rect 7377 10523 7435 10529
rect 7377 10520 7389 10523
rect 5868 10492 7389 10520
rect 5868 10480 5874 10492
rect 7377 10489 7389 10492
rect 7423 10489 7435 10523
rect 8404 10520 8432 10548
rect 9217 10523 9275 10529
rect 9217 10520 9229 10523
rect 8404 10492 9229 10520
rect 7377 10483 7435 10489
rect 9217 10489 9229 10492
rect 9263 10489 9275 10523
rect 9217 10483 9275 10489
rect 9944 10523 10002 10529
rect 9944 10489 9956 10523
rect 9990 10520 10002 10523
rect 10962 10520 10968 10532
rect 9990 10492 10968 10520
rect 9990 10489 10002 10492
rect 9944 10483 10002 10489
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 2590 10412 2596 10464
rect 2648 10452 2654 10464
rect 3513 10455 3571 10461
rect 3513 10452 3525 10455
rect 2648 10424 3525 10452
rect 2648 10412 2654 10424
rect 3513 10421 3525 10424
rect 3559 10421 3571 10455
rect 3513 10415 3571 10421
rect 4249 10455 4307 10461
rect 4249 10421 4261 10455
rect 4295 10452 4307 10455
rect 4798 10452 4804 10464
rect 4295 10424 4804 10452
rect 4295 10421 4307 10424
rect 4249 10415 4307 10421
rect 4798 10412 4804 10424
rect 4856 10452 4862 10464
rect 5350 10452 5356 10464
rect 4856 10424 5356 10452
rect 4856 10412 4862 10424
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 6086 10452 6092 10464
rect 6047 10424 6092 10452
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6546 10452 6552 10464
rect 6227 10424 6552 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6917 10455 6975 10461
rect 6917 10421 6929 10455
rect 6963 10452 6975 10455
rect 7190 10452 7196 10464
rect 6963 10424 7196 10452
rect 6963 10421 6975 10424
rect 6917 10415 6975 10421
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 8846 10452 8852 10464
rect 7340 10424 7385 10452
rect 8807 10424 8852 10452
rect 7340 10412 7346 10424
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 8938 10412 8944 10464
rect 8996 10452 9002 10464
rect 11072 10452 11100 10628
rect 11701 10625 11713 10628
rect 11747 10656 11759 10659
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 11747 10628 13001 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12989 10625 13001 10628
rect 13035 10656 13047 10659
rect 13538 10656 13544 10668
rect 13035 10628 13544 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 14148 10628 14289 10656
rect 14148 10616 14154 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 14550 10656 14556 10668
rect 14507 10628 14556 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 14844 10665 14872 10764
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16206 10792 16212 10804
rect 16167 10764 16212 10792
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 16485 10795 16543 10801
rect 16485 10761 16497 10795
rect 16531 10792 16543 10795
rect 16666 10792 16672 10804
rect 16531 10764 16672 10792
rect 16531 10761 16543 10764
rect 16485 10755 16543 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18874 10792 18880 10804
rect 18371 10764 18880 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 19886 10792 19892 10804
rect 19208 10764 19564 10792
rect 19847 10764 19892 10792
rect 19208 10752 19214 10764
rect 16850 10684 16856 10736
rect 16908 10724 16914 10736
rect 16908 10696 17080 10724
rect 16908 10684 16914 10696
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14700 10628 14841 10656
rect 14700 10616 14706 10628
rect 14829 10625 14841 10628
rect 14875 10625 14887 10659
rect 16942 10656 16948 10668
rect 16903 10628 16948 10656
rect 14829 10619 14887 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17052 10665 17080 10696
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 18156 10628 18644 10656
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11514 10588 11520 10600
rect 11204 10560 11376 10588
rect 11475 10560 11520 10588
rect 11204 10548 11210 10560
rect 8996 10424 11100 10452
rect 8996 10412 9002 10424
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 11348 10452 11376 10560
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 12802 10588 12808 10600
rect 12763 10560 12808 10588
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 13722 10588 13728 10600
rect 13683 10560 13728 10588
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 14108 10560 14596 10588
rect 11609 10523 11667 10529
rect 11609 10489 11621 10523
rect 11655 10520 11667 10523
rect 11698 10520 11704 10532
rect 11655 10492 11704 10520
rect 11655 10489 11667 10492
rect 11609 10483 11667 10489
rect 11698 10480 11704 10492
rect 11756 10480 11762 10532
rect 14108 10520 14136 10560
rect 11808 10492 14136 10520
rect 14185 10523 14243 10529
rect 11808 10452 11836 10492
rect 14185 10489 14197 10523
rect 14231 10520 14243 10523
rect 14366 10520 14372 10532
rect 14231 10492 14372 10520
rect 14231 10489 14243 10492
rect 14185 10483 14243 10489
rect 14366 10480 14372 10492
rect 14424 10480 14430 10532
rect 14568 10520 14596 10560
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15085 10591 15143 10597
rect 15085 10588 15097 10591
rect 14976 10560 15097 10588
rect 14976 10548 14982 10560
rect 15085 10557 15097 10560
rect 15131 10588 15143 10591
rect 16758 10588 16764 10600
rect 15131 10560 16764 10588
rect 15131 10557 15143 10560
rect 15085 10551 15143 10557
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 16853 10591 16911 10597
rect 16853 10557 16865 10591
rect 16899 10588 16911 10591
rect 17954 10588 17960 10600
rect 16899 10560 17960 10588
rect 16899 10557 16911 10560
rect 16853 10551 16911 10557
rect 17954 10548 17960 10560
rect 18012 10548 18018 10600
rect 18156 10597 18184 10628
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 18472 10560 18521 10588
rect 18472 10548 18478 10560
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18616 10588 18644 10628
rect 19536 10588 19564 10764
rect 19886 10752 19892 10764
rect 19944 10752 19950 10804
rect 20070 10752 20076 10804
rect 20128 10792 20134 10804
rect 20349 10795 20407 10801
rect 20349 10792 20361 10795
rect 20128 10764 20361 10792
rect 20128 10752 20134 10764
rect 20349 10761 20361 10764
rect 20395 10761 20407 10795
rect 20349 10755 20407 10761
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 20901 10659 20959 10665
rect 20901 10656 20913 10659
rect 20588 10628 20913 10656
rect 20588 10616 20594 10628
rect 20901 10625 20913 10628
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 18616 10560 19564 10588
rect 18509 10551 18567 10557
rect 17402 10520 17408 10532
rect 14568 10492 17408 10520
rect 17402 10480 17408 10492
rect 17460 10480 17466 10532
rect 17497 10523 17555 10529
rect 17497 10489 17509 10523
rect 17543 10520 17555 10523
rect 18598 10520 18604 10532
rect 17543 10492 18604 10520
rect 17543 10489 17555 10492
rect 17497 10483 17555 10489
rect 18598 10480 18604 10492
rect 18656 10480 18662 10532
rect 18776 10523 18834 10529
rect 18776 10489 18788 10523
rect 18822 10520 18834 10523
rect 20809 10523 20867 10529
rect 20809 10520 20821 10523
rect 18822 10492 19288 10520
rect 18822 10489 18834 10492
rect 18776 10483 18834 10489
rect 19260 10464 19288 10492
rect 20180 10492 20821 10520
rect 11204 10424 11249 10452
rect 11348 10424 11836 10452
rect 12437 10455 12495 10461
rect 11204 10412 11210 10424
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12710 10452 12716 10464
rect 12483 10424 12716 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13170 10452 13176 10464
rect 12943 10424 13176 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 13541 10455 13599 10461
rect 13541 10421 13553 10455
rect 13587 10452 13599 10455
rect 13722 10452 13728 10464
rect 13587 10424 13728 10452
rect 13587 10421 13599 10424
rect 13541 10415 13599 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 13817 10455 13875 10461
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 14090 10452 14096 10464
rect 13863 10424 14096 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 18322 10452 18328 10464
rect 16356 10424 18328 10452
rect 16356 10412 16362 10424
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 18414 10412 18420 10464
rect 18472 10452 18478 10464
rect 19058 10452 19064 10464
rect 18472 10424 19064 10452
rect 18472 10412 18478 10424
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 19242 10412 19248 10464
rect 19300 10412 19306 10464
rect 19702 10412 19708 10464
rect 19760 10452 19766 10464
rect 20180 10461 20208 10492
rect 20809 10489 20821 10492
rect 20855 10489 20867 10523
rect 20809 10483 20867 10489
rect 20165 10455 20223 10461
rect 20165 10452 20177 10455
rect 19760 10424 20177 10452
rect 19760 10412 19766 10424
rect 20165 10421 20177 10424
rect 20211 10421 20223 10455
rect 20714 10452 20720 10464
rect 20675 10424 20720 10452
rect 20165 10415 20223 10421
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 2317 10251 2375 10257
rect 2317 10248 2329 10251
rect 1728 10220 2329 10248
rect 1728 10208 1734 10220
rect 2317 10217 2329 10220
rect 2363 10217 2375 10251
rect 2317 10211 2375 10217
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2455 10220 2973 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2961 10217 2973 10220
rect 3007 10217 3019 10251
rect 2961 10211 3019 10217
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6788 10220 6837 10248
rect 6788 10208 6794 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 7190 10248 7196 10260
rect 7151 10220 7196 10248
rect 6825 10211 6883 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7331 10220 7849 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 8205 10251 8263 10257
rect 8205 10217 8217 10251
rect 8251 10248 8263 10251
rect 8294 10248 8300 10260
rect 8251 10220 8300 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8849 10251 8907 10257
rect 8849 10217 8861 10251
rect 8895 10248 8907 10251
rect 9674 10248 9680 10260
rect 8895 10220 9680 10248
rect 8895 10217 8907 10220
rect 8849 10211 8907 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 11020 10220 11069 10248
rect 11020 10208 11026 10220
rect 11057 10217 11069 10220
rect 11103 10248 11115 10251
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11103 10220 11805 10248
rect 11103 10217 11115 10220
rect 11057 10211 11115 10217
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10248 12403 10251
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 12391 10220 13001 10248
rect 12391 10217 12403 10220
rect 12345 10211 12403 10217
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 12989 10211 13047 10217
rect 13262 10208 13268 10260
rect 13320 10208 13326 10260
rect 13357 10251 13415 10257
rect 13357 10217 13369 10251
rect 13403 10248 13415 10251
rect 13906 10248 13912 10260
rect 13403 10220 13912 10248
rect 13403 10217 13415 10220
rect 13357 10211 13415 10217
rect 13906 10208 13912 10220
rect 13964 10248 13970 10260
rect 15010 10248 15016 10260
rect 13964 10220 15016 10248
rect 13964 10208 13970 10220
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 15749 10251 15807 10257
rect 15749 10217 15761 10251
rect 15795 10248 15807 10251
rect 16114 10248 16120 10260
rect 15795 10220 16120 10248
rect 15795 10217 15807 10220
rect 15749 10211 15807 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 17770 10248 17776 10260
rect 17731 10220 17776 10248
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 18417 10251 18475 10257
rect 18417 10217 18429 10251
rect 18463 10248 18475 10251
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 18463 10220 19809 10248
rect 18463 10217 18475 10220
rect 18417 10211 18475 10217
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 19797 10211 19855 10217
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20772 10220 20913 10248
rect 20772 10208 20778 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 3568 10152 4568 10180
rect 3568 10140 3574 10152
rect 3326 10112 3332 10124
rect 3287 10084 3332 10112
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3878 10112 3884 10124
rect 3467 10084 3884 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 4540 10121 4568 10152
rect 4706 10140 4712 10192
rect 4764 10189 4770 10192
rect 4764 10183 4828 10189
rect 4764 10149 4782 10183
rect 4816 10149 4828 10183
rect 4764 10143 4828 10149
rect 4764 10140 4770 10143
rect 6362 10140 6368 10192
rect 6420 10180 6426 10192
rect 10686 10180 10692 10192
rect 6420 10152 9076 10180
rect 6420 10140 6426 10152
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 4614 10112 4620 10124
rect 4571 10084 4620 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 7653 10115 7711 10121
rect 7653 10112 7665 10115
rect 7484 10084 7665 10112
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10044 3663 10047
rect 3694 10044 3700 10056
rect 3651 10016 3700 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 7484 10053 7512 10084
rect 7653 10081 7665 10084
rect 7699 10081 7711 10115
rect 7653 10075 7711 10081
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 8846 10112 8852 10124
rect 8343 10084 8852 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 9048 10121 9076 10152
rect 9784 10152 10692 10180
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10081 9091 10115
rect 9674 10112 9680 10124
rect 9635 10084 9680 10112
rect 9033 10075 9091 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 8202 10044 8208 10056
rect 7616 10016 8208 10044
rect 7616 10004 7622 10016
rect 8202 10004 8208 10016
rect 8260 10044 8266 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8260 10016 8401 10044
rect 8260 10004 8266 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9784 10044 9812 10152
rect 10686 10140 10692 10152
rect 10744 10180 10750 10192
rect 11517 10183 11575 10189
rect 10744 10152 11468 10180
rect 10744 10140 10750 10152
rect 9950 10121 9956 10124
rect 9944 10075 9956 10121
rect 10008 10112 10014 10124
rect 10008 10084 10044 10112
rect 9950 10072 9956 10075
rect 10008 10072 10014 10084
rect 8628 10016 9812 10044
rect 11440 10044 11468 10152
rect 11517 10149 11529 10183
rect 11563 10180 11575 10183
rect 12618 10180 12624 10192
rect 11563 10152 12624 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 13280 10180 13308 10208
rect 13280 10152 13400 10180
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10112 11851 10115
rect 12437 10115 12495 10121
rect 11839 10084 12204 10112
rect 11839 10081 11851 10084
rect 11793 10075 11851 10081
rect 11440 10016 12112 10044
rect 8628 10004 8634 10016
rect 1946 9976 1952 9988
rect 1907 9948 1952 9976
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 5460 9948 8975 9976
rect 3970 9868 3976 9920
rect 4028 9908 4034 9920
rect 5460 9908 5488 9948
rect 5902 9908 5908 9920
rect 4028 9880 5488 9908
rect 5863 9880 5908 9908
rect 4028 9868 4034 9880
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 7653 9911 7711 9917
rect 7653 9877 7665 9911
rect 7699 9908 7711 9911
rect 8662 9908 8668 9920
rect 7699 9880 8668 9908
rect 7699 9877 7711 9880
rect 7653 9871 7711 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 8947 9908 8975 9948
rect 11790 9908 11796 9920
rect 8947 9880 11796 9908
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 11974 9908 11980 9920
rect 11935 9880 11980 9908
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 12084 9908 12112 10016
rect 12176 9976 12204 10084
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 13262 10112 13268 10124
rect 12483 10084 12664 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 12342 10004 12348 10056
rect 12400 10044 12406 10056
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 12400 10016 12541 10044
rect 12400 10004 12406 10016
rect 12529 10013 12541 10016
rect 12575 10013 12587 10047
rect 12636 10044 12664 10084
rect 12728 10084 13268 10112
rect 12728 10044 12756 10084
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 12636 10016 12756 10044
rect 12529 10007 12587 10013
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 13372 10044 13400 10152
rect 14458 10140 14464 10192
rect 14516 10180 14522 10192
rect 14918 10180 14924 10192
rect 14516 10152 14924 10180
rect 14516 10140 14522 10152
rect 14918 10140 14924 10152
rect 14976 10140 14982 10192
rect 15657 10183 15715 10189
rect 15657 10149 15669 10183
rect 15703 10180 15715 10183
rect 16574 10180 16580 10192
rect 15703 10152 16580 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 18046 10140 18052 10192
rect 18104 10180 18110 10192
rect 19702 10180 19708 10192
rect 18104 10152 19708 10180
rect 18104 10140 18110 10152
rect 19702 10140 19708 10152
rect 19760 10140 19766 10192
rect 19886 10140 19892 10192
rect 19944 10140 19950 10192
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 13688 10084 14381 10112
rect 13688 10072 13694 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 15746 10072 15752 10124
rect 15804 10112 15810 10124
rect 16206 10112 16212 10124
rect 15804 10084 16212 10112
rect 15804 10072 15810 10084
rect 16206 10072 16212 10084
rect 16264 10112 16270 10124
rect 16393 10115 16451 10121
rect 16393 10112 16405 10115
rect 16264 10084 16405 10112
rect 16264 10072 16270 10084
rect 16393 10081 16405 10084
rect 16439 10081 16451 10115
rect 16393 10075 16451 10081
rect 16660 10115 16718 10121
rect 16660 10081 16672 10115
rect 16706 10112 16718 10115
rect 17494 10112 17500 10124
rect 16706 10084 17500 10112
rect 16706 10081 16718 10084
rect 16660 10075 16718 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 18322 10072 18328 10124
rect 18380 10112 18386 10124
rect 18690 10112 18696 10124
rect 18380 10084 18696 10112
rect 18380 10072 18386 10084
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 19904 10112 19932 10140
rect 18831 10084 19012 10112
rect 19904 10084 20024 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 12860 10016 13461 10044
rect 12860 10004 12866 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13596 10016 13641 10044
rect 13596 10004 13602 10016
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 14056 10016 14473 10044
rect 14056 10004 14062 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 14568 9976 14596 10007
rect 14642 10004 14648 10056
rect 14700 10044 14706 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 14700 10016 15853 10044
rect 14700 10004 14706 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 18874 10044 18880 10056
rect 18835 10016 18880 10044
rect 15841 10007 15899 10013
rect 18874 10004 18880 10016
rect 18932 10004 18938 10056
rect 12176 9948 14596 9976
rect 15120 9948 15700 9976
rect 13906 9908 13912 9920
rect 12084 9880 13912 9908
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14001 9911 14059 9917
rect 14001 9877 14013 9911
rect 14047 9908 14059 9911
rect 15120 9908 15148 9948
rect 15286 9908 15292 9920
rect 14047 9880 15148 9908
rect 15247 9880 15292 9908
rect 14047 9877 14059 9880
rect 14001 9871 14059 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15672 9908 15700 9948
rect 17310 9908 17316 9920
rect 15672 9880 17316 9908
rect 17310 9868 17316 9880
rect 17368 9868 17374 9920
rect 18984 9908 19012 10084
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10044 19119 10047
rect 19242 10044 19248 10056
rect 19107 10016 19248 10044
rect 19107 10013 19119 10016
rect 19061 10007 19119 10013
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19886 10044 19892 10056
rect 19847 10016 19892 10044
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 19996 10053 20024 10084
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 19426 9976 19432 9988
rect 19387 9948 19432 9976
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 19058 9908 19064 9920
rect 18984 9880 19064 9908
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 8202 9704 8208 9716
rect 4120 9676 8064 9704
rect 8163 9676 8208 9704
rect 4120 9664 4126 9676
rect 1854 9636 1860 9648
rect 1815 9608 1860 9636
rect 1854 9596 1860 9608
rect 1912 9596 1918 9648
rect 2222 9636 2228 9648
rect 2183 9608 2228 9636
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 8036 9636 8064 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 12526 9704 12532 9716
rect 8312 9676 12532 9704
rect 8312 9636 8340 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 16853 9707 16911 9713
rect 16853 9704 16865 9707
rect 13964 9676 16865 9704
rect 13964 9664 13970 9676
rect 16853 9673 16865 9676
rect 16899 9673 16911 9707
rect 18874 9704 18880 9716
rect 16853 9667 16911 9673
rect 17420 9676 18880 9704
rect 8036 9608 8340 9636
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 13357 9639 13415 9645
rect 13357 9636 13369 9639
rect 11388 9608 13369 9636
rect 11388 9596 11394 9608
rect 13357 9605 13369 9608
rect 13403 9605 13415 9639
rect 13630 9636 13636 9648
rect 13357 9599 13415 9605
rect 13464 9608 13636 9636
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 3510 9568 3516 9580
rect 2915 9540 3516 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3510 9528 3516 9540
rect 3568 9568 3574 9580
rect 3694 9568 3700 9580
rect 3568 9540 3700 9568
rect 3568 9528 3574 9540
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10275 9540 10977 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 10965 9537 10977 9540
rect 11011 9568 11023 9571
rect 12342 9568 12348 9580
rect 11011 9540 12348 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 1670 9500 1676 9512
rect 1631 9472 1676 9500
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2774 9432 2780 9444
rect 2639 9404 2780 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 2774 9392 2780 9404
rect 2832 9392 2838 9444
rect 4065 9435 4123 9441
rect 4065 9401 4077 9435
rect 4111 9432 4123 9435
rect 4172 9432 4200 9460
rect 4356 9432 4384 9531
rect 12342 9528 12348 9540
rect 12400 9568 12406 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12400 9540 13001 9568
rect 12400 9528 12406 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 13464 9568 13492 9608
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 13780 9608 16436 9636
rect 13780 9596 13786 9608
rect 12989 9531 13047 9537
rect 13280 9540 13492 9568
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 4709 9503 4767 9509
rect 4709 9500 4721 9503
rect 4672 9472 4721 9500
rect 4672 9460 4678 9472
rect 4709 9469 4721 9472
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4976 9503 5034 9509
rect 4976 9469 4988 9503
rect 5022 9500 5034 9503
rect 5902 9500 5908 9512
rect 5022 9472 5908 9500
rect 5022 9469 5034 9472
rect 4976 9463 5034 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 6871 9472 8769 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 8757 9469 8769 9472
rect 8803 9500 8815 9503
rect 9766 9500 9772 9512
rect 8803 9472 9772 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9500 10839 9503
rect 11146 9500 11152 9512
rect 10827 9472 11152 9500
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 13280 9500 13308 9540
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13596 9540 14013 9568
rect 13596 9528 13602 9540
rect 14001 9537 14013 9540
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14148 9540 14933 9568
rect 14148 9528 14154 9540
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 15102 9568 15108 9580
rect 15063 9540 15108 9568
rect 14921 9531 14979 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15562 9528 15568 9580
rect 15620 9568 15626 9580
rect 15657 9571 15715 9577
rect 15657 9568 15669 9571
rect 15620 9540 15669 9568
rect 15620 9528 15626 9540
rect 15657 9537 15669 9540
rect 15703 9537 15715 9571
rect 15657 9531 15715 9537
rect 11296 9472 13308 9500
rect 13817 9503 13875 9509
rect 11296 9460 11302 9472
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 14734 9500 14740 9512
rect 13863 9472 14740 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 15286 9500 15292 9512
rect 14875 9472 15292 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 15473 9503 15531 9509
rect 15473 9469 15485 9503
rect 15519 9500 15531 9503
rect 16298 9500 16304 9512
rect 15519 9472 16304 9500
rect 15519 9469 15531 9472
rect 15473 9463 15531 9469
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 16408 9509 16436 9608
rect 16482 9596 16488 9648
rect 16540 9636 16546 9648
rect 17420 9636 17448 9676
rect 18874 9664 18880 9676
rect 18932 9664 18938 9716
rect 16540 9608 17448 9636
rect 16540 9596 16546 9608
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 19613 9639 19671 9645
rect 19613 9636 19625 9639
rect 19300 9608 19625 9636
rect 19300 9596 19306 9608
rect 19613 9605 19625 9608
rect 19659 9605 19671 9639
rect 19978 9636 19984 9648
rect 19939 9608 19984 9636
rect 19613 9599 19671 9605
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 17589 9571 17647 9577
rect 17460 9540 17505 9568
rect 17460 9528 17466 9540
rect 17589 9537 17601 9571
rect 17635 9568 17647 9571
rect 19628 9568 19656 9599
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 20530 9568 20536 9580
rect 17635 9540 18368 9568
rect 19628 9540 20536 9568
rect 17635 9537 17647 9540
rect 17589 9531 17647 9537
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9500 16911 9503
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 16899 9472 17325 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 5534 9432 5540 9444
rect 4111 9404 4292 9432
rect 4356 9404 5540 9432
rect 4111 9401 4123 9404
rect 4065 9395 4123 9401
rect 2685 9367 2743 9373
rect 2685 9333 2697 9367
rect 2731 9364 2743 9367
rect 3234 9364 3240 9376
rect 2731 9336 3240 9364
rect 2731 9333 2743 9336
rect 2685 9327 2743 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3694 9364 3700 9376
rect 3655 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4154 9364 4160 9376
rect 4115 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 4264 9364 4292 9404
rect 5534 9392 5540 9404
rect 5592 9432 5598 9444
rect 5592 9404 6132 9432
rect 5592 9392 5598 9404
rect 4890 9364 4896 9376
rect 4264 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 6104 9373 6132 9404
rect 7006 9392 7012 9444
rect 7064 9441 7070 9444
rect 7064 9435 7128 9441
rect 7064 9401 7082 9435
rect 7116 9432 7128 9435
rect 8478 9432 8484 9444
rect 7116 9404 8484 9432
rect 7116 9401 7128 9404
rect 7064 9395 7128 9401
rect 7064 9392 7070 9395
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 8938 9392 8944 9444
rect 8996 9441 9002 9444
rect 8996 9435 9060 9441
rect 8996 9401 9014 9435
rect 9048 9401 9060 9435
rect 8996 9395 9060 9401
rect 8996 9392 9002 9395
rect 9582 9392 9588 9444
rect 9640 9432 9646 9444
rect 10873 9435 10931 9441
rect 10873 9432 10885 9435
rect 9640 9404 10885 9432
rect 9640 9392 9646 9404
rect 10873 9401 10885 9404
rect 10919 9401 10931 9435
rect 10873 9395 10931 9401
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 13357 9435 13415 9441
rect 12851 9404 13216 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 6089 9367 6147 9373
rect 6089 9333 6101 9367
rect 6135 9333 6147 9367
rect 10134 9364 10140 9376
rect 10047 9336 10140 9364
rect 6089 9327 6147 9333
rect 10134 9324 10140 9336
rect 10192 9364 10198 9376
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 10192 9336 10241 9364
rect 10192 9324 10198 9336
rect 10229 9333 10241 9336
rect 10275 9333 10287 9367
rect 10229 9327 10287 9333
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10778 9364 10784 9376
rect 10459 9336 10784 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 11664 9336 12449 9364
rect 11664 9324 11670 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12437 9327 12495 9333
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13188 9364 13216 9404
rect 13357 9401 13369 9435
rect 13403 9432 13415 9435
rect 15930 9432 15936 9444
rect 13403 9404 14596 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 13188 9336 13461 9364
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14090 9364 14096 9376
rect 13964 9336 14096 9364
rect 13964 9324 13970 9336
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14458 9364 14464 9376
rect 14419 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14568 9364 14596 9404
rect 14844 9404 15936 9432
rect 14844 9364 14872 9404
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 18248 9432 18276 9463
rect 16500 9404 18276 9432
rect 18340 9432 18368 9540
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 18506 9441 18512 9444
rect 18500 9432 18512 9441
rect 18340 9404 18512 9432
rect 16206 9364 16212 9376
rect 14568 9336 14872 9364
rect 16167 9336 16212 9364
rect 16206 9324 16212 9336
rect 16264 9364 16270 9376
rect 16500 9364 16528 9404
rect 16942 9364 16948 9376
rect 16264 9336 16528 9364
rect 16903 9336 16948 9364
rect 16264 9324 16270 9336
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 18248 9364 18276 9404
rect 18500 9395 18512 9404
rect 18506 9392 18512 9395
rect 18564 9392 18570 9444
rect 19426 9392 19432 9444
rect 19484 9432 19490 9444
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 19484 9404 20453 9432
rect 19484 9392 19490 9404
rect 20441 9401 20453 9404
rect 20487 9401 20499 9435
rect 20441 9395 20499 9401
rect 18414 9364 18420 9376
rect 18248 9336 18420 9364
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 18690 9324 18696 9376
rect 18748 9364 18754 9376
rect 20349 9367 20407 9373
rect 20349 9364 20361 9367
rect 18748 9336 20361 9364
rect 18748 9324 18754 9336
rect 20349 9333 20361 9336
rect 20395 9333 20407 9367
rect 20349 9327 20407 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 3605 9163 3663 9169
rect 3605 9160 3617 9163
rect 3568 9132 3617 9160
rect 3568 9120 3574 9132
rect 3605 9129 3617 9132
rect 3651 9129 3663 9163
rect 3605 9123 3663 9129
rect 3694 9120 3700 9172
rect 3752 9160 3758 9172
rect 5905 9163 5963 9169
rect 5905 9160 5917 9163
rect 3752 9132 5917 9160
rect 3752 9120 3758 9132
rect 5905 9129 5917 9132
rect 5951 9129 5963 9163
rect 5905 9123 5963 9129
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 7282 9160 7288 9172
rect 6871 9132 7288 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 11330 9160 11336 9172
rect 7392 9132 11336 9160
rect 1670 9052 1676 9104
rect 1728 9092 1734 9104
rect 1765 9095 1823 9101
rect 1765 9092 1777 9095
rect 1728 9064 1777 9092
rect 1728 9052 1734 9064
rect 1765 9061 1777 9064
rect 1811 9061 1823 9095
rect 1765 9055 1823 9061
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 7392 9092 7420 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12253 9163 12311 9169
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 12894 9160 12900 9172
rect 12299 9132 12900 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13262 9160 13268 9172
rect 13223 9132 13268 9160
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 13814 9160 13820 9172
rect 13740 9132 13820 9160
rect 7558 9101 7564 9104
rect 7552 9092 7564 9101
rect 4120 9064 7420 9092
rect 7519 9064 7564 9092
rect 4120 9052 4126 9064
rect 7552 9055 7564 9064
rect 7558 9052 7564 9055
rect 7616 9052 7622 9104
rect 9944 9095 10002 9101
rect 9944 9061 9956 9095
rect 9990 9092 10002 9095
rect 10134 9092 10140 9104
rect 9990 9064 10140 9092
rect 9990 9061 10002 9064
rect 9944 9055 10002 9061
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10318 9052 10324 9104
rect 10376 9092 10382 9104
rect 11238 9092 11244 9104
rect 10376 9064 11244 9092
rect 10376 9052 10382 9064
rect 11238 9052 11244 9064
rect 11296 9052 11302 9104
rect 13633 9095 13691 9101
rect 13633 9061 13645 9095
rect 13679 9092 13691 9095
rect 13740 9092 13768 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 15470 9160 15476 9172
rect 14332 9132 15476 9160
rect 14332 9120 14338 9132
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 17494 9160 17500 9172
rect 17455 9132 17500 9160
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 17865 9163 17923 9169
rect 17865 9129 17877 9163
rect 17911 9160 17923 9163
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 17911 9132 19257 9160
rect 17911 9129 17923 9132
rect 17865 9123 17923 9129
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 13679 9064 13768 9092
rect 13679 9061 13691 9064
rect 13633 9055 13691 9061
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 14553 9095 14611 9101
rect 14553 9092 14565 9095
rect 14240 9064 14565 9092
rect 14240 9052 14246 9064
rect 14553 9061 14565 9064
rect 14599 9061 14611 9095
rect 14553 9055 14611 9061
rect 16942 9052 16948 9104
rect 17000 9092 17006 9104
rect 19337 9095 19395 9101
rect 19337 9092 19349 9095
rect 17000 9064 19349 9092
rect 17000 9052 17006 9064
rect 19337 9061 19349 9064
rect 19383 9061 19395 9095
rect 19337 9055 19395 9061
rect 1486 9024 1492 9036
rect 1447 8996 1492 9024
rect 1486 8984 1492 8996
rect 1544 8984 1550 9036
rect 2130 8984 2136 9036
rect 2188 9024 2194 9036
rect 2225 9027 2283 9033
rect 2225 9024 2237 9027
rect 2188 8996 2237 9024
rect 2188 8984 2194 8996
rect 2225 8993 2237 8996
rect 2271 8993 2283 9027
rect 2225 8987 2283 8993
rect 2492 9027 2550 9033
rect 2492 8993 2504 9027
rect 2538 9024 2550 9027
rect 3050 9024 3056 9036
rect 2538 8996 3056 9024
rect 2538 8993 2550 8996
rect 2492 8987 2550 8993
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 3878 8984 3884 9036
rect 3936 9024 3942 9036
rect 4893 9027 4951 9033
rect 4893 9024 4905 9027
rect 3936 8996 4905 9024
rect 3936 8984 3942 8996
rect 4893 8993 4905 8996
rect 4939 8993 4951 9027
rect 7006 9024 7012 9036
rect 4893 8987 4951 8993
rect 5184 8996 7012 9024
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 4798 8956 4804 8968
rect 3292 8928 4804 8956
rect 3292 8916 3298 8928
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 5184 8965 5212 8996
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 9674 9024 9680 9036
rect 7331 8996 9680 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 12066 9024 12072 9036
rect 9784 8996 12072 9024
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4856 8928 4997 8956
rect 4856 8916 4862 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8925 5227 8959
rect 5810 8956 5816 8968
rect 5169 8919 5227 8925
rect 5552 8928 5816 8956
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 5552 8888 5580 8928
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8925 6147 8959
rect 9784 8956 9812 8996
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 12161 9027 12219 9033
rect 12161 8993 12173 9027
rect 12207 9024 12219 9027
rect 12250 9024 12256 9036
rect 12207 8996 12256 9024
rect 12207 8993 12219 8996
rect 12161 8987 12219 8993
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 12621 9027 12679 9033
rect 12621 9024 12633 9027
rect 12584 8996 12633 9024
rect 12584 8984 12590 8996
rect 12621 8993 12633 8996
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 9024 12771 9027
rect 13262 9024 13268 9036
rect 12759 8996 13268 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 6089 8919 6147 8925
rect 8312 8928 9812 8956
rect 4571 8860 5580 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 6104 8888 6132 8919
rect 5684 8860 6132 8888
rect 5684 8848 5690 8860
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 4764 8792 5549 8820
rect 4764 8780 4770 8792
rect 5537 8789 5549 8792
rect 5583 8789 5595 8823
rect 5537 8783 5595 8789
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 8312 8820 8340 8928
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 12728 8956 12756 8987
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 9024 13783 9027
rect 13771 8996 14044 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 10928 8928 12756 8956
rect 12897 8959 12955 8965
rect 10928 8916 10934 8928
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 13446 8956 13452 8968
rect 12943 8928 13452 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 13814 8956 13820 8968
rect 13775 8928 13820 8956
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 14016 8956 14044 8996
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 14332 8996 14377 9024
rect 14332 8984 14338 8996
rect 15930 8984 15936 9036
rect 15988 9024 15994 9036
rect 16117 9027 16175 9033
rect 16117 9024 16129 9027
rect 15988 8996 16129 9024
rect 15988 8984 15994 8996
rect 16117 8993 16129 8996
rect 16163 9024 16175 9027
rect 16206 9024 16212 9036
rect 16163 8996 16212 9024
rect 16163 8993 16175 8996
rect 16117 8987 16175 8993
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 16384 9027 16442 9033
rect 16384 8993 16396 9027
rect 16430 9024 16442 9027
rect 17402 9024 17408 9036
rect 16430 8996 17408 9024
rect 16430 8993 16442 8996
rect 16384 8987 16442 8993
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 17920 8996 18245 9024
rect 17920 8984 17926 8996
rect 18233 8993 18245 8996
rect 18279 8993 18291 9027
rect 18233 8987 18291 8993
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 9024 18383 9027
rect 18782 9024 18788 9036
rect 18371 8996 18788 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 19794 8984 19800 9036
rect 19852 9024 19858 9036
rect 20073 9027 20131 9033
rect 20073 9024 20085 9027
rect 19852 8996 20085 9024
rect 19852 8984 19858 8996
rect 20073 8993 20085 8996
rect 20119 8993 20131 9027
rect 20073 8987 20131 8993
rect 14182 8956 14188 8968
rect 14016 8928 14188 8956
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 18506 8956 18512 8968
rect 18467 8928 18512 8956
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19300 8928 19441 8956
rect 19300 8916 19306 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 13906 8848 13912 8900
rect 13964 8888 13970 8900
rect 14550 8888 14556 8900
rect 13964 8860 14556 8888
rect 13964 8848 13970 8860
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 17218 8848 17224 8900
rect 17276 8888 17282 8900
rect 18690 8888 18696 8900
rect 17276 8860 18696 8888
rect 17276 8848 17282 8860
rect 18690 8848 18696 8860
rect 18748 8848 18754 8900
rect 18877 8891 18935 8897
rect 18877 8857 18889 8891
rect 18923 8888 18935 8891
rect 19886 8888 19892 8900
rect 18923 8860 19892 8888
rect 18923 8857 18935 8860
rect 18877 8851 18935 8857
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 8662 8820 8668 8832
rect 5960 8792 8340 8820
rect 8623 8792 8668 8820
rect 5960 8780 5966 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10962 8820 10968 8832
rect 10008 8792 10968 8820
rect 10008 8780 10014 8792
rect 10962 8780 10968 8792
rect 11020 8820 11026 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 11020 8792 11069 8820
rect 11020 8780 11026 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 11977 8823 12035 8829
rect 11977 8789 11989 8823
rect 12023 8820 12035 8823
rect 12066 8820 12072 8832
rect 12023 8792 12072 8820
rect 12023 8789 12035 8792
rect 11977 8783 12035 8789
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 20272 8820 20300 8919
rect 12492 8792 20300 8820
rect 12492 8780 12498 8792
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 5534 8616 5540 8628
rect 4939 8588 5540 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 9585 8619 9643 8625
rect 9585 8585 9597 8619
rect 9631 8616 9643 8619
rect 10318 8616 10324 8628
rect 9631 8588 10324 8616
rect 9631 8585 9643 8588
rect 9585 8579 9643 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 11974 8616 11980 8628
rect 10520 8588 11980 8616
rect 4065 8551 4123 8557
rect 4065 8517 4077 8551
rect 4111 8548 4123 8551
rect 4111 8520 5488 8548
rect 4111 8517 4123 8520
rect 4065 8511 4123 8517
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 3936 8452 4537 8480
rect 3936 8440 3942 8452
rect 4525 8449 4537 8452
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4755 8452 4905 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5460 8421 5488 8520
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 1940 8415 1998 8421
rect 1940 8381 1952 8415
rect 1986 8412 1998 8415
rect 5445 8415 5503 8421
rect 1986 8384 5304 8412
rect 1986 8381 1998 8384
rect 1940 8375 1998 8381
rect 1688 8344 1716 8375
rect 2130 8344 2136 8356
rect 1688 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8344 2194 8356
rect 4154 8344 4160 8356
rect 2188 8316 4160 8344
rect 2188 8304 2194 8316
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4433 8347 4491 8353
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 4982 8344 4988 8356
rect 4479 8316 4988 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 4982 8304 4988 8316
rect 5040 8304 5046 8356
rect 5276 8344 5304 8384
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 5644 8356 5672 8443
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 10008 8452 10149 8480
rect 10008 8440 10014 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 10520 8412 10548 8588
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 13004 8588 14688 8616
rect 10597 8551 10655 8557
rect 10597 8517 10609 8551
rect 10643 8517 10655 8551
rect 10597 8511 10655 8517
rect 10091 8384 10548 8412
rect 10612 8412 10640 8511
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 11020 8520 11192 8548
rect 11020 8508 11026 8520
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11164 8489 11192 8520
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10836 8452 11069 8480
rect 10836 8440 10842 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12526 8480 12532 8492
rect 12216 8452 12532 8480
rect 12216 8440 12222 8452
rect 12526 8440 12532 8452
rect 12584 8480 12590 8492
rect 13004 8489 13032 8588
rect 14369 8551 14427 8557
rect 14369 8517 14381 8551
rect 14415 8548 14427 8551
rect 14553 8551 14611 8557
rect 14553 8548 14565 8551
rect 14415 8520 14565 8548
rect 14415 8517 14427 8520
rect 14369 8511 14427 8517
rect 14553 8517 14565 8520
rect 14599 8517 14611 8551
rect 14553 8511 14611 8517
rect 14660 8489 14688 8588
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 16298 8616 16304 8628
rect 15068 8588 15700 8616
rect 16259 8588 16304 8616
rect 15068 8576 15074 8588
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12584 8452 13001 8480
rect 12584 8440 12590 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 13256 8415 13314 8421
rect 10612 8384 12940 8412
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 5626 8344 5632 8356
rect 5276 8316 5632 8344
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 9953 8347 10011 8353
rect 9953 8313 9965 8347
rect 9999 8344 10011 8347
rect 11146 8344 11152 8356
rect 9999 8316 11152 8344
rect 9999 8313 10011 8316
rect 9953 8307 10011 8313
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 11606 8344 11612 8356
rect 11256 8316 11612 8344
rect 5074 8276 5080 8288
rect 5035 8248 5080 8276
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5537 8279 5595 8285
rect 5537 8276 5549 8279
rect 5224 8248 5549 8276
rect 5224 8236 5230 8248
rect 5537 8245 5549 8248
rect 5583 8245 5595 8279
rect 5537 8239 5595 8245
rect 10965 8279 11023 8285
rect 10965 8245 10977 8279
rect 11011 8276 11023 8279
rect 11256 8276 11284 8316
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 12912 8344 12940 8384
rect 13256 8381 13268 8415
rect 13302 8412 13314 8415
rect 15672 8412 15700 8588
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 18506 8576 18512 8628
rect 18564 8616 18570 8628
rect 20165 8619 20223 8625
rect 20165 8616 20177 8619
rect 18564 8588 20177 8616
rect 18564 8576 18570 8588
rect 20165 8585 20177 8588
rect 20211 8585 20223 8619
rect 20165 8579 20223 8585
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 20717 8619 20775 8625
rect 20717 8616 20729 8619
rect 20680 8588 20729 8616
rect 20680 8576 20686 8588
rect 20717 8585 20729 8588
rect 20763 8585 20775 8619
rect 20717 8579 20775 8585
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 17494 8480 17500 8492
rect 16991 8452 17500 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 18656 8452 18797 8480
rect 18656 8440 18662 8452
rect 18785 8449 18797 8452
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 13302 8384 15148 8412
rect 15672 8384 19012 8412
rect 13302 8381 13314 8384
rect 13256 8375 13314 8381
rect 15120 8356 15148 8384
rect 13998 8344 14004 8356
rect 12912 8316 14004 8344
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 14550 8344 14556 8356
rect 14463 8316 14556 8344
rect 14550 8304 14556 8316
rect 14608 8344 14614 8356
rect 14890 8347 14948 8353
rect 14890 8344 14902 8347
rect 14608 8316 14902 8344
rect 14608 8304 14614 8316
rect 14890 8313 14902 8316
rect 14936 8313 14948 8347
rect 14890 8307 14948 8313
rect 15102 8304 15108 8356
rect 15160 8304 15166 8356
rect 16666 8344 16672 8356
rect 16627 8316 16672 8344
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 11011 8248 11284 8276
rect 11011 8245 11023 8248
rect 10965 8239 11023 8245
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 15194 8276 15200 8288
rect 11940 8248 15200 8276
rect 11940 8236 11946 8248
rect 15194 8236 15200 8248
rect 15252 8236 15258 8288
rect 16022 8276 16028 8288
rect 15983 8248 16028 8276
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 16758 8276 16764 8288
rect 16719 8248 16764 8276
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 18984 8276 19012 8384
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 19392 8384 20545 8412
rect 19392 8372 19398 8384
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 20533 8375 20591 8381
rect 19052 8347 19110 8353
rect 19052 8313 19064 8347
rect 19098 8344 19110 8347
rect 20438 8344 20444 8356
rect 19098 8316 20444 8344
rect 19098 8313 19110 8316
rect 19052 8307 19110 8313
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 19242 8276 19248 8288
rect 18984 8248 19248 8276
rect 19242 8236 19248 8248
rect 19300 8236 19306 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 1544 8044 2605 8072
rect 1544 8032 1550 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 5074 8072 5080 8084
rect 3007 8044 5080 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 5626 8072 5632 8084
rect 5583 8044 5632 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 5813 8075 5871 8081
rect 5813 8041 5825 8075
rect 5859 8072 5871 8075
rect 5994 8072 6000 8084
rect 5859 8044 6000 8072
rect 5859 8041 5871 8044
rect 5813 8035 5871 8041
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 10410 8072 10416 8084
rect 10275 8044 10416 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 11204 8044 12541 8072
rect 11204 8032 11210 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 12529 8035 12587 8041
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12768 8044 13001 8072
rect 12768 8032 12774 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 14093 8075 14151 8081
rect 14093 8041 14105 8075
rect 14139 8072 14151 8075
rect 14274 8072 14280 8084
rect 14139 8044 14280 8072
rect 14139 8041 14151 8044
rect 14093 8035 14151 8041
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14516 8044 14565 8072
rect 14516 8032 14522 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14553 8035 14611 8041
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 16724 8044 17693 8072
rect 16724 8032 16730 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 4706 8004 4712 8016
rect 3099 7976 4712 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 5718 7964 5724 8016
rect 5776 8004 5782 8016
rect 6273 8007 6331 8013
rect 6273 8004 6285 8007
rect 5776 7976 6285 8004
rect 5776 7964 5782 7976
rect 6273 7973 6285 7976
rect 6319 7973 6331 8007
rect 6273 7967 6331 7973
rect 9858 7964 9864 8016
rect 9916 8004 9922 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9916 7976 10333 8004
rect 9916 7964 9922 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 11790 8004 11796 8016
rect 10321 7967 10379 7973
rect 10520 7976 11796 8004
rect 4154 7936 4160 7948
rect 4115 7908 4160 7936
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 4424 7939 4482 7945
rect 4424 7905 4436 7939
rect 4470 7936 4482 7939
rect 5534 7936 5540 7948
rect 4470 7908 5540 7936
rect 4470 7905 4482 7908
rect 4424 7899 4482 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 6144 7908 6193 7936
rect 6144 7896 6150 7908
rect 6181 7905 6193 7908
rect 6227 7936 6239 7939
rect 6227 7908 10364 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 3142 7868 3148 7880
rect 3103 7840 3148 7868
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 5552 7868 5580 7896
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 5552 7840 6377 7868
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 10042 7800 10048 7812
rect 5092 7772 10048 7800
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 5092 7732 5120 7772
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 10336 7800 10364 7908
rect 10520 7877 10548 7976
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 12897 8007 12955 8013
rect 12897 8004 12909 8007
rect 12676 7976 12909 8004
rect 12676 7964 12682 7976
rect 12897 7973 12909 7976
rect 12943 7973 12955 8007
rect 12897 7967 12955 7973
rect 14292 7976 14780 8004
rect 10873 7939 10931 7945
rect 10873 7905 10885 7939
rect 10919 7936 10931 7939
rect 10962 7936 10968 7948
rect 10919 7908 10968 7936
rect 10919 7905 10931 7908
rect 10873 7899 10931 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11140 7939 11198 7945
rect 11140 7905 11152 7939
rect 11186 7936 11198 7939
rect 11698 7936 11704 7948
rect 11186 7908 11704 7936
rect 11186 7905 11198 7908
rect 11140 7899 11198 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 14292 7936 14320 7976
rect 14458 7936 14464 7948
rect 12032 7908 14320 7936
rect 14419 7908 14464 7936
rect 12032 7896 12038 7908
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 14752 7936 14780 7976
rect 16022 7964 16028 8016
rect 16080 8004 16086 8016
rect 16270 8007 16328 8013
rect 16270 8004 16282 8007
rect 16080 7976 16282 8004
rect 16080 7964 16086 7976
rect 16270 7973 16282 7976
rect 16316 7973 16328 8007
rect 16270 7967 16328 7973
rect 19236 8007 19294 8013
rect 19236 7973 19248 8007
rect 19282 8004 19294 8007
rect 19518 8004 19524 8016
rect 19282 7976 19524 8004
rect 19282 7973 19294 7976
rect 19236 7967 19294 7973
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 16850 7936 16856 7948
rect 14752 7908 16856 7936
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 18012 7908 18061 7936
rect 18012 7896 18018 7908
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 18141 7939 18199 7945
rect 18141 7905 18153 7939
rect 18187 7936 18199 7939
rect 18506 7936 18512 7948
rect 18187 7908 18512 7936
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 18506 7896 18512 7908
rect 18564 7896 18570 7948
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18969 7939 19027 7945
rect 18969 7936 18981 7939
rect 18656 7908 18981 7936
rect 18656 7896 18662 7908
rect 18969 7905 18981 7908
rect 19015 7936 19027 7939
rect 19058 7936 19064 7948
rect 19015 7908 19064 7936
rect 19015 7905 19027 7908
rect 18969 7899 19027 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12400 7840 13093 7868
rect 12400 7828 12406 7840
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 14550 7828 14556 7880
rect 14608 7868 14614 7880
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 14608 7840 14657 7868
rect 14608 7828 14614 7840
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 15988 7840 16037 7868
rect 15988 7828 15994 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 10870 7800 10876 7812
rect 10336 7772 10876 7800
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 12526 7800 12532 7812
rect 12124 7772 12532 7800
rect 12124 7760 12130 7772
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 17402 7800 17408 7812
rect 17363 7772 17408 7800
rect 17402 7760 17408 7772
rect 17460 7800 17466 7812
rect 18248 7800 18276 7831
rect 20162 7828 20168 7880
rect 20220 7868 20226 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20220 7840 20913 7868
rect 20220 7828 20226 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 17460 7772 18276 7800
rect 17460 7760 17466 7772
rect 4120 7704 5120 7732
rect 9861 7735 9919 7741
rect 4120 7692 4126 7704
rect 9861 7701 9873 7735
rect 9907 7732 9919 7735
rect 11606 7732 11612 7744
rect 9907 7704 11612 7732
rect 9907 7701 9919 7704
rect 9861 7695 9919 7701
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 12250 7732 12256 7744
rect 12211 7704 12256 7732
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 16942 7732 16948 7744
rect 12400 7704 16948 7732
rect 12400 7692 12406 7704
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 20346 7732 20352 7744
rect 20307 7704 20352 7732
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 3973 7531 4031 7537
rect 3973 7497 3985 7531
rect 4019 7528 4031 7531
rect 5166 7528 5172 7540
rect 4019 7500 5172 7528
rect 4019 7497 4031 7500
rect 3973 7491 4031 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 11698 7528 11704 7540
rect 10560 7500 11560 7528
rect 11659 7500 11704 7528
rect 10560 7488 10566 7500
rect 5534 7460 5540 7472
rect 4632 7432 5540 7460
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 3602 7392 3608 7404
rect 992 7364 3608 7392
rect 992 7352 998 7364
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 4632 7401 4660 7432
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 11532 7460 11560 7500
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 13170 7528 13176 7540
rect 12492 7500 13176 7528
rect 12492 7488 12498 7500
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 15160 7500 15485 7528
rect 15160 7488 15166 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 16758 7528 16764 7540
rect 16255 7500 16764 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 18012 7500 18061 7528
rect 18012 7488 18018 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 20438 7528 20444 7540
rect 20399 7500 20444 7528
rect 18049 7491 18107 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 12342 7460 12348 7472
rect 11532 7432 12348 7460
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 13817 7463 13875 7469
rect 13817 7429 13829 7463
rect 13863 7460 13875 7463
rect 13906 7460 13912 7472
rect 13863 7432 13912 7460
rect 13863 7429 13875 7432
rect 13817 7423 13875 7429
rect 13906 7420 13912 7432
rect 13964 7420 13970 7472
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4982 7392 4988 7404
rect 4943 7364 4988 7392
rect 4617 7355 4675 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9732 7364 10333 7392
rect 9732 7352 9738 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 13924 7392 13952 7420
rect 16853 7395 16911 7401
rect 13924 7364 14228 7392
rect 10321 7355 10379 7361
rect 11882 7324 11888 7336
rect 10428 7296 11888 7324
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 10428 7256 10456 7296
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 12158 7324 12164 7336
rect 11992 7296 12164 7324
rect 4120 7228 10456 7256
rect 10588 7259 10646 7265
rect 4120 7216 4126 7228
rect 10588 7225 10600 7259
rect 10634 7256 10646 7259
rect 10870 7256 10876 7268
rect 10634 7228 10876 7256
rect 10634 7225 10646 7228
rect 10588 7219 10646 7225
rect 10870 7216 10876 7228
rect 10928 7216 10934 7268
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11992 7256 12020 7296
rect 12158 7284 12164 7296
rect 12216 7324 12222 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12216 7296 12449 7324
rect 12216 7284 12222 7296
rect 12437 7293 12449 7296
rect 12483 7324 12495 7327
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 12483 7296 14105 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14200 7324 14228 7364
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 17402 7392 17408 7404
rect 16899 7364 17408 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 18322 7352 18328 7404
rect 18380 7392 18386 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18380 7364 18613 7392
rect 18380 7352 18386 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 19058 7392 19064 7404
rect 19019 7364 19064 7392
rect 18601 7355 18659 7361
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 14349 7327 14407 7333
rect 14349 7324 14361 7327
rect 14200 7296 14361 7324
rect 14093 7287 14151 7293
rect 14349 7293 14361 7296
rect 14395 7324 14407 7327
rect 15930 7324 15936 7336
rect 14395 7296 15936 7324
rect 14395 7293 14407 7296
rect 14349 7287 14407 7293
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7324 18567 7327
rect 20806 7324 20812 7336
rect 18555 7296 20812 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 11112 7228 12020 7256
rect 11112 7216 11118 7228
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12682 7259 12740 7265
rect 12682 7256 12694 7259
rect 12308 7228 12694 7256
rect 12308 7216 12314 7228
rect 12682 7225 12694 7228
rect 12728 7225 12740 7259
rect 12682 7219 12740 7225
rect 13170 7216 13176 7268
rect 13228 7256 13234 7268
rect 18524 7256 18552 7287
rect 20806 7284 20812 7296
rect 20864 7284 20870 7336
rect 13228 7228 18552 7256
rect 19328 7259 19386 7265
rect 13228 7216 13234 7228
rect 19328 7225 19340 7259
rect 19374 7256 19386 7259
rect 20346 7256 20352 7268
rect 19374 7228 20352 7256
rect 19374 7225 19386 7228
rect 19328 7219 19386 7225
rect 20346 7216 20352 7228
rect 20404 7216 20410 7268
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4304 7160 4353 7188
rect 4304 7148 4310 7160
rect 4341 7157 4353 7160
rect 4387 7157 4399 7191
rect 4341 7151 4399 7157
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4798 7188 4804 7200
rect 4479 7160 4804 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 11974 7188 11980 7200
rect 9916 7160 11980 7188
rect 9916 7148 9922 7160
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 15286 7188 15292 7200
rect 12584 7160 15292 7188
rect 12584 7148 12590 7160
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 16574 7188 16580 7200
rect 16535 7160 16580 7188
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 17497 7191 17555 7197
rect 16724 7160 16769 7188
rect 16724 7148 16730 7160
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 18417 7191 18475 7197
rect 18417 7188 18429 7191
rect 17543 7160 18429 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 18417 7157 18429 7160
rect 18463 7157 18475 7191
rect 18417 7151 18475 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6984 11667 6987
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 11655 6956 12173 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 12161 6953 12173 6956
rect 12207 6953 12219 6987
rect 12161 6947 12219 6953
rect 12621 6987 12679 6993
rect 12621 6953 12633 6987
rect 12667 6984 12679 6987
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 12667 6956 13185 6984
rect 12667 6953 12679 6956
rect 12621 6947 12679 6953
rect 13173 6953 13185 6956
rect 13219 6953 13231 6987
rect 13630 6984 13636 6996
rect 13591 6956 13636 6984
rect 13173 6947 13231 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 14185 6987 14243 6993
rect 14185 6953 14197 6987
rect 14231 6984 14243 6987
rect 14458 6984 14464 6996
rect 14231 6956 14464 6984
rect 14231 6953 14243 6956
rect 14185 6947 14243 6953
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 14553 6987 14611 6993
rect 14553 6953 14565 6987
rect 14599 6984 14611 6987
rect 15289 6987 15347 6993
rect 15289 6984 15301 6987
rect 14599 6956 15301 6984
rect 14599 6953 14611 6956
rect 14553 6947 14611 6953
rect 15289 6953 15301 6956
rect 15335 6953 15347 6987
rect 15289 6947 15347 6953
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 15749 6987 15807 6993
rect 15749 6984 15761 6987
rect 15528 6956 15761 6984
rect 15528 6944 15534 6956
rect 15749 6953 15761 6956
rect 15795 6953 15807 6987
rect 15749 6947 15807 6953
rect 18049 6987 18107 6993
rect 18049 6953 18061 6987
rect 18095 6984 18107 6987
rect 18598 6984 18604 6996
rect 18095 6956 18604 6984
rect 18095 6953 18107 6956
rect 18049 6947 18107 6953
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 20162 6984 20168 6996
rect 20123 6956 20168 6984
rect 20162 6944 20168 6956
rect 20220 6944 20226 6996
rect 10980 6888 13216 6916
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 10980 6848 11008 6888
rect 4028 6820 11008 6848
rect 4028 6808 4034 6820
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 11112 6820 11529 6848
rect 11112 6808 11118 6820
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 12526 6848 12532 6860
rect 12487 6820 12532 6848
rect 11517 6811 11575 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 13188 6848 13216 6888
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 13541 6919 13599 6925
rect 13541 6916 13553 6919
rect 13412 6888 13553 6916
rect 13412 6876 13418 6888
rect 13541 6885 13553 6888
rect 13587 6916 13599 6919
rect 16761 6919 16819 6925
rect 16761 6916 16773 6919
rect 13587 6888 16773 6916
rect 13587 6885 13599 6888
rect 13541 6879 13599 6885
rect 16761 6885 16773 6888
rect 16807 6885 16819 6919
rect 18322 6916 18328 6928
rect 16761 6879 16819 6885
rect 17052 6888 18328 6916
rect 15470 6848 15476 6860
rect 13188 6820 15476 6848
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15654 6848 15660 6860
rect 15615 6820 15660 6848
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16448 6820 16681 6848
rect 16448 6808 16454 6820
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 16669 6811 16727 6817
rect 17052 6792 17080 6888
rect 18322 6876 18328 6888
rect 18380 6876 18386 6928
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6780 11851 6783
rect 12250 6780 12256 6792
rect 11839 6752 12256 6780
rect 11839 6749 11851 6752
rect 11793 6743 11851 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 4120 6684 11284 6712
rect 4120 6672 4126 6684
rect 11146 6644 11152 6656
rect 11107 6616 11152 6644
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 11256 6644 11284 6684
rect 11698 6672 11704 6724
rect 11756 6712 11762 6724
rect 12728 6712 12756 6743
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14642 6780 14648 6792
rect 13780 6752 13825 6780
rect 14603 6752 14648 6780
rect 13780 6740 13786 6752
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 15102 6780 15108 6792
rect 14875 6752 15108 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 15930 6780 15936 6792
rect 15891 6752 15936 6780
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 16080 6752 16865 6780
rect 16080 6740 16086 6752
rect 16853 6749 16865 6752
rect 16899 6780 16911 6783
rect 17034 6780 17040 6792
rect 16899 6752 17040 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 18138 6780 18144 6792
rect 18099 6752 18144 6780
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18340 6789 18368 6876
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 20070 6740 20076 6792
rect 20128 6780 20134 6792
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 20128 6752 20269 6780
rect 20128 6740 20134 6752
rect 20257 6749 20269 6752
rect 20303 6749 20315 6783
rect 20438 6780 20444 6792
rect 20399 6752 20444 6780
rect 20257 6743 20315 6749
rect 20438 6740 20444 6752
rect 20496 6740 20502 6792
rect 11756 6684 12756 6712
rect 16301 6715 16359 6721
rect 11756 6672 11762 6684
rect 16301 6681 16313 6715
rect 16347 6712 16359 6715
rect 16574 6712 16580 6724
rect 16347 6684 16580 6712
rect 16347 6681 16359 6684
rect 16301 6675 16359 6681
rect 16574 6672 16580 6684
rect 16632 6672 16638 6724
rect 17681 6715 17739 6721
rect 17681 6681 17693 6715
rect 17727 6712 17739 6715
rect 18506 6712 18512 6724
rect 17727 6684 18512 6712
rect 17727 6681 17739 6684
rect 17681 6675 17739 6681
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 19794 6712 19800 6724
rect 19755 6684 19800 6712
rect 19794 6672 19800 6684
rect 19852 6672 19858 6724
rect 12434 6644 12440 6656
rect 11256 6616 12440 6644
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 10965 6443 11023 6449
rect 10965 6409 10977 6443
rect 11011 6440 11023 6443
rect 11054 6440 11060 6452
rect 11011 6412 11060 6440
rect 11011 6409 11023 6412
rect 10965 6403 11023 6409
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 12526 6440 12532 6452
rect 12483 6412 12532 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14700 6412 14841 6440
rect 14700 6400 14706 6412
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 15194 6400 15200 6452
rect 15252 6440 15258 6452
rect 15654 6440 15660 6452
rect 15252 6412 15660 6440
rect 15252 6400 15258 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 16485 6443 16543 6449
rect 16485 6409 16497 6443
rect 16531 6440 16543 6443
rect 16666 6440 16672 6452
rect 16531 6412 16672 6440
rect 16531 6409 16543 6412
rect 16485 6403 16543 6409
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 20070 6440 20076 6452
rect 20031 6412 20076 6440
rect 20070 6400 20076 6412
rect 20128 6400 20134 6452
rect 5442 6332 5448 6384
rect 5500 6372 5506 6384
rect 17954 6372 17960 6384
rect 5500 6344 17960 6372
rect 5500 6332 5506 6344
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 11609 6307 11667 6313
rect 11609 6273 11621 6307
rect 11655 6304 11667 6307
rect 11698 6304 11704 6316
rect 11655 6276 11704 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 11940 6276 13093 6304
rect 11940 6264 11946 6276
rect 13081 6273 13093 6276
rect 13127 6304 13139 6307
rect 13722 6304 13728 6316
rect 13127 6276 13728 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6304 14427 6307
rect 15194 6304 15200 6316
rect 14415 6276 15200 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15473 6307 15531 6313
rect 15335 6276 15424 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 11333 6239 11391 6245
rect 11333 6236 11345 6239
rect 11204 6208 11345 6236
rect 11204 6196 11210 6208
rect 11333 6205 11345 6208
rect 11379 6205 11391 6239
rect 11333 6199 11391 6205
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6236 12955 6239
rect 12943 6208 14964 6236
rect 12943 6205 12955 6208
rect 12897 6199 12955 6205
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 11974 6168 11980 6180
rect 10652 6140 11980 6168
rect 10652 6128 10658 6140
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 12805 6171 12863 6177
rect 12805 6137 12817 6171
rect 12851 6168 12863 6171
rect 13814 6168 13820 6180
rect 12851 6140 13820 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 14936 6168 14964 6208
rect 15396 6168 15424 6276
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15930 6304 15936 6316
rect 15519 6276 15936 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 17034 6304 17040 6316
rect 16995 6276 17040 6304
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 20346 6264 20352 6316
rect 20404 6304 20410 6316
rect 20625 6307 20683 6313
rect 20625 6304 20637 6307
rect 20404 6276 20637 6304
rect 20404 6264 20410 6276
rect 20625 6273 20637 6276
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 16942 6236 16948 6248
rect 16899 6208 16948 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 18046 6168 18052 6180
rect 14936 6140 15332 6168
rect 15396 6140 18052 6168
rect 11422 6100 11428 6112
rect 11383 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 15194 6100 15200 6112
rect 15155 6072 15200 6100
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15304 6100 15332 6140
rect 18046 6128 18052 6140
rect 18104 6128 18110 6180
rect 16390 6100 16396 6112
rect 15304 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 16945 6103 17003 6109
rect 16945 6100 16957 6103
rect 16908 6072 16957 6100
rect 16908 6060 16914 6072
rect 16945 6069 16957 6072
rect 16991 6069 17003 6103
rect 19886 6100 19892 6112
rect 19847 6072 19892 6100
rect 16945 6063 17003 6069
rect 19886 6060 19892 6072
rect 19944 6100 19950 6112
rect 20441 6103 20499 6109
rect 20441 6100 20453 6103
rect 19944 6072 20453 6100
rect 19944 6060 19950 6072
rect 20441 6069 20453 6072
rect 20487 6069 20499 6103
rect 20441 6063 20499 6069
rect 20530 6060 20536 6112
rect 20588 6100 20594 6112
rect 20588 6072 20633 6100
rect 20588 6060 20594 6072
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 10321 5899 10379 5905
rect 10321 5865 10333 5899
rect 10367 5896 10379 5899
rect 11422 5896 11428 5908
rect 10367 5868 11428 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 19886 5896 19892 5908
rect 11532 5868 19892 5896
rect 3142 5788 3148 5840
rect 3200 5828 3206 5840
rect 11532 5828 11560 5868
rect 19886 5856 19892 5868
rect 19944 5856 19950 5908
rect 3200 5800 11560 5828
rect 11600 5831 11658 5837
rect 3200 5788 3206 5800
rect 11600 5797 11612 5831
rect 11646 5828 11658 5831
rect 11790 5828 11796 5840
rect 11646 5800 11796 5828
rect 11646 5797 11658 5800
rect 11600 5791 11658 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 11974 5788 11980 5840
rect 12032 5828 12038 5840
rect 17954 5828 17960 5840
rect 12032 5800 17960 5828
rect 12032 5788 12038 5800
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 10689 5763 10747 5769
rect 10689 5760 10701 5763
rect 4212 5732 10701 5760
rect 4212 5720 4218 5732
rect 10689 5729 10701 5732
rect 10735 5729 10747 5763
rect 11882 5760 11888 5772
rect 10689 5723 10747 5729
rect 10980 5732 11888 5760
rect 10980 5704 11008 5732
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 18138 5760 18144 5772
rect 15252 5732 18144 5760
rect 15252 5720 15258 5732
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 10652 5664 10793 5692
rect 10652 5652 10658 5664
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 10962 5692 10968 5704
rect 10923 5664 10968 5692
rect 10781 5655 10839 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11333 5695 11391 5701
rect 11333 5692 11345 5695
rect 11112 5664 11345 5692
rect 11112 5652 11118 5664
rect 11333 5661 11345 5664
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12713 5559 12771 5565
rect 12713 5556 12725 5559
rect 12032 5528 12725 5556
rect 12032 5516 12038 5528
rect 12713 5525 12725 5528
rect 12759 5525 12771 5559
rect 12713 5519 12771 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 11204 5324 11345 5352
rect 11204 5312 11210 5324
rect 11333 5321 11345 5324
rect 11379 5321 11391 5355
rect 11333 5315 11391 5321
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 18506 5352 18512 5364
rect 13872 5324 18512 5352
rect 13872 5312 13878 5324
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 4120 5188 11805 5216
rect 4120 5176 4126 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 11808 5148 11836 5179
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 11940 5188 11985 5216
rect 11940 5176 11946 5188
rect 17218 5148 17224 5160
rect 11808 5120 17224 5148
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 11701 5083 11759 5089
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 12437 5083 12495 5089
rect 12437 5080 12449 5083
rect 11747 5052 12449 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 12437 5049 12449 5052
rect 12483 5049 12495 5083
rect 12437 5043 12495 5049
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 5350 4128 5356 4140
rect 4120 4100 5356 4128
rect 4120 4088 4126 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 17954 4128 17960 4140
rect 12860 4100 17960 4128
rect 12860 4088 12866 4100
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 11054 3720 11060 3732
rect 10704 3692 11060 3720
rect 10704 3593 10732 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11790 3680 11796 3732
rect 11848 3720 11854 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 11848 3692 12081 3720
rect 11848 3680 11854 3692
rect 12069 3689 12081 3692
rect 12115 3689 12127 3723
rect 12069 3683 12127 3689
rect 10956 3655 11014 3661
rect 10956 3621 10968 3655
rect 11002 3652 11014 3655
rect 11146 3652 11152 3664
rect 11002 3624 11152 3652
rect 11002 3621 11014 3624
rect 10956 3615 11014 3621
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3553 10747 3587
rect 18966 3584 18972 3596
rect 10689 3547 10747 3553
rect 10796 3556 18972 3584
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 10796 3516 10824 3556
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 8720 3488 10824 3516
rect 8720 3476 8726 3488
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 3326 2048 3332 2100
rect 3384 2088 3390 2100
rect 4798 2088 4804 2100
rect 3384 2060 4804 2088
rect 3384 2048 3390 2060
rect 4798 2048 4804 2060
rect 4856 2048 4862 2100
rect 14090 2048 14096 2100
rect 14148 2088 14154 2100
rect 18506 2088 18512 2100
rect 14148 2060 18512 2088
rect 14148 2048 14154 2060
rect 18506 2048 18512 2060
rect 18564 2048 18570 2100
rect 3142 688 3148 740
rect 3200 728 3206 740
rect 4890 728 4896 740
rect 3200 700 4896 728
rect 3200 688 3206 700
rect 4890 688 4896 700
rect 4948 688 4954 740
rect 3326 280 3332 332
rect 3384 320 3390 332
rect 5258 320 5264 332
rect 3384 292 5264 320
rect 3384 280 3390 292
rect 5258 280 5264 292
rect 5316 280 5322 332
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 13452 20000 13504 20052
rect 13912 20000 13964 20052
rect 14464 20000 14516 20052
rect 15384 20000 15436 20052
rect 15936 20000 15988 20052
rect 17776 20000 17828 20052
rect 18236 20000 18288 20052
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20628 20000 20680 20052
rect 6644 19932 6696 19984
rect 3148 19864 3200 19916
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 12900 19864 12952 19916
rect 3240 19796 3292 19848
rect 12164 19796 12216 19848
rect 13544 19864 13596 19916
rect 14096 19864 14148 19916
rect 15476 19864 15528 19916
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 3332 19728 3384 19780
rect 16580 19864 16632 19916
rect 17316 19796 17368 19848
rect 17960 19864 18012 19916
rect 19892 19864 19944 19916
rect 19984 19907 20036 19916
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 19800 19796 19852 19848
rect 17132 19728 17184 19780
rect 19616 19771 19668 19780
rect 19616 19737 19625 19771
rect 19625 19737 19659 19771
rect 19659 19737 19668 19771
rect 19616 19728 19668 19737
rect 2504 19703 2556 19712
rect 2504 19669 2513 19703
rect 2513 19669 2547 19703
rect 2547 19669 2556 19703
rect 2504 19660 2556 19669
rect 3424 19660 3476 19712
rect 3608 19703 3660 19712
rect 3608 19669 3617 19703
rect 3617 19669 3651 19703
rect 3651 19669 3660 19703
rect 3608 19660 3660 19669
rect 12716 19703 12768 19712
rect 12716 19669 12725 19703
rect 12725 19669 12759 19703
rect 12759 19669 12768 19703
rect 12716 19660 12768 19669
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 3700 19499 3752 19508
rect 3700 19465 3709 19499
rect 3709 19465 3743 19499
rect 3743 19465 3752 19499
rect 3700 19456 3752 19465
rect 3792 19456 3844 19508
rect 17960 19456 18012 19508
rect 2780 19388 2832 19440
rect 2596 19295 2648 19304
rect 2596 19261 2605 19295
rect 2605 19261 2639 19295
rect 2639 19261 2648 19295
rect 2596 19252 2648 19261
rect 3700 19320 3752 19372
rect 3792 19252 3844 19304
rect 3884 19252 3936 19304
rect 2872 19116 2924 19168
rect 3056 19116 3108 19168
rect 3608 19116 3660 19168
rect 4528 19252 4580 19304
rect 5816 19388 5868 19440
rect 4712 19320 4764 19372
rect 8944 19320 8996 19372
rect 4804 19252 4856 19304
rect 9864 19252 9916 19304
rect 11428 19295 11480 19304
rect 11428 19261 11437 19295
rect 11437 19261 11471 19295
rect 11471 19261 11480 19295
rect 11428 19252 11480 19261
rect 11980 19320 12032 19372
rect 12164 19320 12216 19372
rect 12900 19320 12952 19372
rect 12532 19252 12584 19304
rect 13176 19295 13228 19304
rect 13176 19261 13185 19295
rect 13185 19261 13219 19295
rect 13219 19261 13228 19295
rect 13176 19252 13228 19261
rect 14188 19252 14240 19304
rect 14832 19252 14884 19304
rect 14924 19252 14976 19304
rect 19984 19388 20036 19440
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 17868 19320 17920 19372
rect 18972 19320 19024 19372
rect 4988 19116 5040 19168
rect 10508 19116 10560 19168
rect 13268 19184 13320 19236
rect 13452 19227 13504 19236
rect 13452 19193 13486 19227
rect 13486 19193 13504 19227
rect 16580 19252 16632 19304
rect 13452 19184 13504 19193
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 15016 19116 15068 19168
rect 15200 19116 15252 19168
rect 15384 19116 15436 19168
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 16120 19116 16172 19168
rect 18696 19252 18748 19304
rect 20352 19252 20404 19304
rect 19340 19227 19392 19236
rect 19340 19193 19349 19227
rect 19349 19193 19383 19227
rect 19383 19193 19392 19227
rect 19340 19184 19392 19193
rect 17592 19116 17644 19168
rect 17960 19116 18012 19168
rect 19248 19116 19300 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 2964 18912 3016 18964
rect 3056 18912 3108 18964
rect 7380 18912 7432 18964
rect 8300 18955 8352 18964
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 8760 18912 8812 18964
rect 10968 18912 11020 18964
rect 13452 18955 13504 18964
rect 2596 18844 2648 18896
rect 3700 18844 3752 18896
rect 4988 18844 5040 18896
rect 2228 18776 2280 18828
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 7012 18776 7064 18828
rect 7104 18776 7156 18828
rect 10324 18819 10376 18828
rect 10324 18785 10333 18819
rect 10333 18785 10367 18819
rect 10367 18785 10376 18819
rect 10324 18776 10376 18785
rect 12440 18844 12492 18896
rect 13176 18844 13228 18896
rect 13452 18921 13461 18955
rect 13461 18921 13495 18955
rect 13495 18921 13504 18955
rect 13452 18912 13504 18921
rect 15108 18912 15160 18964
rect 15660 18912 15712 18964
rect 20444 18955 20496 18964
rect 1124 18640 1176 18692
rect 3424 18708 3476 18760
rect 3608 18708 3660 18760
rect 6368 18751 6420 18760
rect 4712 18572 4764 18624
rect 6368 18717 6377 18751
rect 6377 18717 6411 18751
rect 6411 18717 6420 18751
rect 6368 18708 6420 18717
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 7288 18708 7340 18760
rect 9128 18708 9180 18760
rect 9680 18708 9732 18760
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 11612 18708 11664 18760
rect 9956 18683 10008 18692
rect 4896 18572 4948 18624
rect 5448 18572 5500 18624
rect 5908 18615 5960 18624
rect 5908 18581 5917 18615
rect 5917 18581 5951 18615
rect 5951 18581 5960 18615
rect 5908 18572 5960 18581
rect 9036 18572 9088 18624
rect 9956 18649 9965 18683
rect 9965 18649 9999 18683
rect 9999 18649 10008 18683
rect 9956 18640 10008 18649
rect 11704 18683 11756 18692
rect 11704 18649 11713 18683
rect 11713 18649 11747 18683
rect 11747 18649 11756 18683
rect 11704 18640 11756 18649
rect 13360 18776 13412 18828
rect 15384 18776 15436 18828
rect 15752 18844 15804 18896
rect 20076 18844 20128 18896
rect 20444 18921 20453 18955
rect 20453 18921 20487 18955
rect 20487 18921 20496 18955
rect 20444 18912 20496 18921
rect 22468 18844 22520 18896
rect 16580 18776 16632 18828
rect 17868 18819 17920 18828
rect 14004 18708 14056 18760
rect 14648 18751 14700 18760
rect 14648 18717 14657 18751
rect 14657 18717 14691 18751
rect 14691 18717 14700 18751
rect 14648 18708 14700 18717
rect 14832 18751 14884 18760
rect 14832 18717 14841 18751
rect 14841 18717 14875 18751
rect 14875 18717 14884 18751
rect 14832 18708 14884 18717
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 17868 18785 17902 18819
rect 17902 18785 17920 18819
rect 17868 18776 17920 18785
rect 18788 18776 18840 18828
rect 19248 18819 19300 18828
rect 19248 18785 19257 18819
rect 19257 18785 19291 18819
rect 19291 18785 19300 18819
rect 19248 18776 19300 18785
rect 19524 18751 19576 18760
rect 12072 18640 12124 18692
rect 15292 18640 15344 18692
rect 15844 18572 15896 18624
rect 15936 18572 15988 18624
rect 16580 18572 16632 18624
rect 16672 18572 16724 18624
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 19984 18776 20036 18828
rect 21548 18776 21600 18828
rect 18880 18640 18932 18692
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 2320 18368 2372 18420
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 4160 18300 4212 18352
rect 6184 18368 6236 18420
rect 6368 18368 6420 18420
rect 5632 18343 5684 18352
rect 5632 18309 5641 18343
rect 5641 18309 5675 18343
rect 5675 18309 5684 18343
rect 5632 18300 5684 18309
rect 6460 18300 6512 18352
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 5356 18232 5408 18284
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 7564 18232 7616 18284
rect 2228 18164 2280 18216
rect 2964 18164 3016 18216
rect 4160 18164 4212 18216
rect 5448 18164 5500 18216
rect 7104 18164 7156 18216
rect 8300 18368 8352 18420
rect 8392 18368 8444 18420
rect 10048 18368 10100 18420
rect 10600 18368 10652 18420
rect 12532 18411 12584 18420
rect 12532 18377 12541 18411
rect 12541 18377 12575 18411
rect 12575 18377 12584 18411
rect 12532 18368 12584 18377
rect 13176 18368 13228 18420
rect 11612 18300 11664 18352
rect 12716 18232 12768 18284
rect 13360 18232 13412 18284
rect 14004 18232 14056 18284
rect 15292 18368 15344 18420
rect 15568 18368 15620 18420
rect 15752 18368 15804 18420
rect 16304 18368 16356 18420
rect 17500 18368 17552 18420
rect 17776 18368 17828 18420
rect 17960 18368 18012 18420
rect 15844 18300 15896 18352
rect 16672 18300 16724 18352
rect 18880 18368 18932 18420
rect 19156 18368 19208 18420
rect 18236 18300 18288 18352
rect 20904 18343 20956 18352
rect 8116 18164 8168 18216
rect 17868 18232 17920 18284
rect 18880 18232 18932 18284
rect 19800 18232 19852 18284
rect 3792 18096 3844 18148
rect 4988 18096 5040 18148
rect 5356 18096 5408 18148
rect 16580 18164 16632 18216
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 16948 18164 17000 18216
rect 18788 18164 18840 18216
rect 19432 18207 19484 18216
rect 19432 18173 19441 18207
rect 19441 18173 19475 18207
rect 19475 18173 19484 18207
rect 19432 18164 19484 18173
rect 20904 18309 20913 18343
rect 20913 18309 20947 18343
rect 20947 18309 20956 18343
rect 20904 18300 20956 18309
rect 20720 18207 20772 18216
rect 20720 18173 20729 18207
rect 20729 18173 20763 18207
rect 20763 18173 20772 18207
rect 20720 18164 20772 18173
rect 664 18028 716 18080
rect 2596 18028 2648 18080
rect 9128 18096 9180 18148
rect 7748 18028 7800 18080
rect 8392 18028 8444 18080
rect 9772 18096 9824 18148
rect 10876 18096 10928 18148
rect 11612 18096 11664 18148
rect 11060 18028 11112 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 13084 18028 13136 18080
rect 14832 18139 14884 18148
rect 14832 18105 14866 18139
rect 14866 18105 14884 18139
rect 14832 18096 14884 18105
rect 15844 18096 15896 18148
rect 18052 18096 18104 18148
rect 14188 18028 14240 18080
rect 15200 18028 15252 18080
rect 18604 18028 18656 18080
rect 18788 18028 18840 18080
rect 19708 18028 19760 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 3056 17867 3108 17876
rect 3056 17833 3065 17867
rect 3065 17833 3099 17867
rect 3099 17833 3108 17867
rect 3056 17824 3108 17833
rect 4252 17824 4304 17876
rect 5080 17824 5132 17876
rect 7012 17867 7064 17876
rect 7012 17833 7021 17867
rect 7021 17833 7055 17867
rect 7055 17833 7064 17867
rect 7012 17824 7064 17833
rect 10416 17824 10468 17876
rect 11704 17824 11756 17876
rect 2688 17756 2740 17808
rect 9956 17756 10008 17808
rect 10508 17799 10560 17808
rect 10508 17765 10542 17799
rect 10542 17765 10560 17799
rect 10508 17756 10560 17765
rect 2136 17731 2188 17740
rect 2136 17697 2155 17731
rect 2155 17697 2188 17731
rect 2136 17688 2188 17697
rect 4252 17688 4304 17740
rect 5632 17731 5684 17740
rect 4620 17620 4672 17672
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 5632 17697 5666 17731
rect 5666 17697 5684 17731
rect 5632 17688 5684 17697
rect 7012 17688 7064 17740
rect 9312 17688 9364 17740
rect 9404 17688 9456 17740
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 9036 17663 9088 17672
rect 9036 17629 9045 17663
rect 9045 17629 9079 17663
rect 9079 17629 9088 17663
rect 9036 17620 9088 17629
rect 9772 17620 9824 17672
rect 10048 17688 10100 17740
rect 13728 17824 13780 17876
rect 14004 17824 14056 17876
rect 14280 17824 14332 17876
rect 14464 17824 14516 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15108 17756 15160 17808
rect 12532 17688 12584 17740
rect 14372 17688 14424 17740
rect 14556 17731 14608 17740
rect 14556 17697 14565 17731
rect 14565 17697 14599 17731
rect 14599 17697 14608 17731
rect 14556 17688 14608 17697
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 16212 17824 16264 17876
rect 20444 17824 20496 17876
rect 16580 17799 16632 17808
rect 16580 17765 16589 17799
rect 16589 17765 16623 17799
rect 16623 17765 16632 17799
rect 16580 17756 16632 17765
rect 18972 17756 19024 17808
rect 19432 17756 19484 17808
rect 16028 17688 16080 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 18052 17688 18104 17740
rect 19984 17731 20036 17740
rect 19984 17697 19993 17731
rect 19993 17697 20027 17731
rect 20027 17697 20036 17731
rect 19984 17688 20036 17697
rect 15016 17620 15068 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 15936 17620 15988 17672
rect 17960 17663 18012 17672
rect 17960 17629 17969 17663
rect 17969 17629 18003 17663
rect 18003 17629 18012 17663
rect 17960 17620 18012 17629
rect 9680 17552 9732 17604
rect 1768 17527 1820 17536
rect 1768 17493 1777 17527
rect 1777 17493 1811 17527
rect 1811 17493 1820 17527
rect 1768 17484 1820 17493
rect 2504 17484 2556 17536
rect 4160 17484 4212 17536
rect 6000 17484 6052 17536
rect 6736 17527 6788 17536
rect 6736 17493 6745 17527
rect 6745 17493 6779 17527
rect 6779 17493 6788 17527
rect 6736 17484 6788 17493
rect 6828 17484 6880 17536
rect 8852 17484 8904 17536
rect 9128 17484 9180 17536
rect 9956 17484 10008 17536
rect 12164 17552 12216 17604
rect 13636 17552 13688 17604
rect 17224 17552 17276 17604
rect 11612 17527 11664 17536
rect 11612 17493 11621 17527
rect 11621 17493 11655 17527
rect 11655 17493 11664 17527
rect 11612 17484 11664 17493
rect 13728 17484 13780 17536
rect 16580 17484 16632 17536
rect 17500 17484 17552 17536
rect 18604 17484 18656 17536
rect 19340 17527 19392 17536
rect 19340 17493 19349 17527
rect 19349 17493 19383 17527
rect 19383 17493 19392 17527
rect 19340 17484 19392 17493
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 2780 17280 2832 17332
rect 4804 17280 4856 17332
rect 5540 17280 5592 17332
rect 2504 17144 2556 17196
rect 5448 17212 5500 17264
rect 4988 17144 5040 17196
rect 7564 17280 7616 17332
rect 9312 17323 9364 17332
rect 9312 17289 9321 17323
rect 9321 17289 9355 17323
rect 9355 17289 9364 17323
rect 9312 17280 9364 17289
rect 10324 17323 10376 17332
rect 10324 17289 10333 17323
rect 10333 17289 10367 17323
rect 10367 17289 10376 17323
rect 10324 17280 10376 17289
rect 10508 17280 10560 17332
rect 19984 17280 20036 17332
rect 4896 17076 4948 17128
rect 5080 17119 5132 17128
rect 5080 17085 5089 17119
rect 5089 17085 5123 17119
rect 5123 17085 5132 17119
rect 6828 17212 6880 17264
rect 8208 17212 8260 17264
rect 12348 17212 12400 17264
rect 13636 17255 13688 17264
rect 5908 17144 5960 17196
rect 6736 17144 6788 17196
rect 9956 17187 10008 17196
rect 6000 17119 6052 17128
rect 5080 17076 5132 17085
rect 6000 17085 6009 17119
rect 6009 17085 6043 17119
rect 6043 17085 6052 17119
rect 6000 17076 6052 17085
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 2964 17008 3016 17060
rect 3516 17008 3568 17060
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 2596 16940 2648 16992
rect 4160 16940 4212 16992
rect 4804 16940 4856 16992
rect 5356 17008 5408 17060
rect 10600 17076 10652 17128
rect 11060 17076 11112 17128
rect 12440 17076 12492 17128
rect 9404 17008 9456 17060
rect 7748 16940 7800 16992
rect 13636 17221 13645 17255
rect 13645 17221 13679 17255
rect 13679 17221 13688 17255
rect 13636 17212 13688 17221
rect 14372 17212 14424 17264
rect 19616 17255 19668 17264
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 14280 17144 14332 17196
rect 19616 17221 19625 17255
rect 19625 17221 19659 17255
rect 19659 17221 19668 17255
rect 19616 17212 19668 17221
rect 13268 17076 13320 17128
rect 10692 16940 10744 16992
rect 10968 16940 11020 16992
rect 11428 16940 11480 16992
rect 12348 16940 12400 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 14280 17008 14332 17060
rect 15844 17119 15896 17128
rect 15844 17085 15853 17119
rect 15853 17085 15887 17119
rect 15887 17085 15896 17119
rect 15844 17076 15896 17085
rect 17960 17144 18012 17196
rect 16856 17076 16908 17128
rect 15476 17008 15528 17060
rect 16764 17008 16816 17060
rect 17408 17008 17460 17060
rect 19340 17076 19392 17128
rect 20168 17076 20220 17128
rect 19800 17008 19852 17060
rect 20444 17051 20496 17060
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 15016 16940 15068 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 17592 16940 17644 16992
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 20444 17017 20453 17051
rect 20453 17017 20487 17051
rect 20487 17017 20496 17051
rect 20444 17008 20496 17017
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 4252 16736 4304 16788
rect 4712 16736 4764 16788
rect 4896 16736 4948 16788
rect 6736 16736 6788 16788
rect 7564 16736 7616 16788
rect 10508 16779 10560 16788
rect 8208 16668 8260 16720
rect 8576 16668 8628 16720
rect 9220 16668 9272 16720
rect 3056 16600 3108 16652
rect 3884 16600 3936 16652
rect 5080 16600 5132 16652
rect 5908 16600 5960 16652
rect 6736 16600 6788 16652
rect 7380 16600 7432 16652
rect 7564 16600 7616 16652
rect 10508 16745 10517 16779
rect 10517 16745 10551 16779
rect 10551 16745 10560 16779
rect 10508 16736 10560 16745
rect 10968 16779 11020 16788
rect 10968 16745 10977 16779
rect 10977 16745 11011 16779
rect 11011 16745 11020 16779
rect 10968 16736 11020 16745
rect 11704 16736 11756 16788
rect 12256 16736 12308 16788
rect 14280 16736 14332 16788
rect 14464 16736 14516 16788
rect 16672 16736 16724 16788
rect 17408 16779 17460 16788
rect 17408 16745 17417 16779
rect 17417 16745 17451 16779
rect 17451 16745 17460 16779
rect 17408 16736 17460 16745
rect 18512 16736 18564 16788
rect 18696 16736 18748 16788
rect 12716 16668 12768 16720
rect 14832 16668 14884 16720
rect 20076 16668 20128 16720
rect 11428 16600 11480 16652
rect 11704 16600 11756 16652
rect 15016 16600 15068 16652
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 15936 16600 15988 16652
rect 16672 16600 16724 16652
rect 17868 16600 17920 16652
rect 19432 16600 19484 16652
rect 19800 16600 19852 16652
rect 1952 16575 2004 16584
rect 1952 16541 1961 16575
rect 1961 16541 1995 16575
rect 1995 16541 2004 16575
rect 1952 16532 2004 16541
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 5816 16532 5868 16584
rect 1584 16507 1636 16516
rect 1584 16473 1593 16507
rect 1593 16473 1627 16507
rect 1627 16473 1636 16507
rect 1584 16464 1636 16473
rect 5172 16464 5224 16516
rect 7380 16464 7432 16516
rect 8576 16464 8628 16516
rect 8668 16464 8720 16516
rect 2964 16396 3016 16448
rect 4988 16396 5040 16448
rect 5540 16396 5592 16448
rect 10140 16532 10192 16584
rect 10968 16532 11020 16584
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11980 16532 12032 16584
rect 12532 16532 12584 16584
rect 13268 16575 13320 16584
rect 13268 16541 13277 16575
rect 13277 16541 13311 16575
rect 13311 16541 13320 16575
rect 13268 16532 13320 16541
rect 15844 16532 15896 16584
rect 19616 16532 19668 16584
rect 20168 16575 20220 16584
rect 20168 16541 20177 16575
rect 20177 16541 20211 16575
rect 20211 16541 20220 16575
rect 20168 16532 20220 16541
rect 9588 16396 9640 16448
rect 10416 16396 10468 16448
rect 15752 16396 15804 16448
rect 16396 16396 16448 16448
rect 20720 16464 20772 16516
rect 17224 16396 17276 16448
rect 19892 16396 19944 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 3884 16235 3936 16244
rect 3884 16201 3893 16235
rect 3893 16201 3927 16235
rect 3927 16201 3936 16235
rect 3884 16192 3936 16201
rect 4160 16192 4212 16244
rect 5356 16192 5408 16244
rect 8668 16192 8720 16244
rect 11612 16192 11664 16244
rect 11704 16192 11756 16244
rect 12716 16192 12768 16244
rect 14372 16192 14424 16244
rect 16304 16192 16356 16244
rect 16672 16192 16724 16244
rect 16764 16192 16816 16244
rect 1952 16056 2004 16108
rect 4068 16124 4120 16176
rect 7288 16124 7340 16176
rect 11520 16124 11572 16176
rect 12532 16124 12584 16176
rect 13912 16124 13964 16176
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 11704 16056 11756 16108
rect 11888 16056 11940 16108
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 2320 15988 2372 16040
rect 2504 16031 2556 16040
rect 2504 15997 2513 16031
rect 2513 15997 2547 16031
rect 2547 15997 2556 16031
rect 2504 15988 2556 15997
rect 4988 15988 5040 16040
rect 5724 15988 5776 16040
rect 8668 16031 8720 16040
rect 8668 15997 8702 16031
rect 8702 15997 8720 16031
rect 2044 15963 2096 15972
rect 2044 15929 2053 15963
rect 2053 15929 2087 15963
rect 2087 15929 2096 15963
rect 2044 15920 2096 15929
rect 4068 15920 4120 15972
rect 1492 15852 1544 15904
rect 3332 15852 3384 15904
rect 4160 15895 4212 15904
rect 4160 15861 4169 15895
rect 4169 15861 4203 15895
rect 4203 15861 4212 15895
rect 4160 15852 4212 15861
rect 5448 15920 5500 15972
rect 8668 15988 8720 15997
rect 7012 15895 7064 15904
rect 7012 15861 7021 15895
rect 7021 15861 7055 15895
rect 7055 15861 7064 15895
rect 7012 15852 7064 15861
rect 7380 15895 7432 15904
rect 7380 15861 7389 15895
rect 7389 15861 7423 15895
rect 7423 15861 7432 15895
rect 7380 15852 7432 15861
rect 7472 15895 7524 15904
rect 7472 15861 7481 15895
rect 7481 15861 7515 15895
rect 7515 15861 7524 15895
rect 8852 15920 8904 15972
rect 7472 15852 7524 15861
rect 9496 15852 9548 15904
rect 11980 15988 12032 16040
rect 12624 15988 12676 16040
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 19064 16192 19116 16244
rect 18788 16124 18840 16176
rect 17960 16056 18012 16108
rect 18696 16056 18748 16108
rect 17684 15988 17736 16040
rect 12992 15920 13044 15972
rect 11152 15852 11204 15904
rect 11428 15895 11480 15904
rect 11428 15861 11437 15895
rect 11437 15861 11471 15895
rect 11471 15861 11480 15895
rect 11428 15852 11480 15861
rect 12164 15852 12216 15904
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 12440 15852 12492 15861
rect 14464 15852 14516 15904
rect 15016 15920 15068 15972
rect 17224 15920 17276 15972
rect 19616 15988 19668 16040
rect 19524 15920 19576 15972
rect 16120 15852 16172 15904
rect 16396 15852 16448 15904
rect 16488 15852 16540 15904
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 17040 15852 17092 15904
rect 19800 15920 19852 15972
rect 20168 15895 20220 15904
rect 20168 15861 20177 15895
rect 20177 15861 20211 15895
rect 20211 15861 20220 15895
rect 20168 15852 20220 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 4160 15648 4212 15700
rect 4068 15580 4120 15632
rect 5816 15648 5868 15700
rect 7472 15648 7524 15700
rect 8208 15691 8260 15700
rect 8208 15657 8217 15691
rect 8217 15657 8251 15691
rect 8251 15657 8260 15691
rect 8208 15648 8260 15657
rect 8852 15691 8904 15700
rect 8852 15657 8861 15691
rect 8861 15657 8895 15691
rect 8895 15657 8904 15691
rect 8852 15648 8904 15657
rect 11520 15648 11572 15700
rect 12164 15691 12216 15700
rect 12164 15657 12173 15691
rect 12173 15657 12207 15691
rect 12207 15657 12216 15691
rect 12164 15648 12216 15657
rect 5172 15580 5224 15632
rect 7104 15580 7156 15632
rect 8576 15580 8628 15632
rect 8760 15580 8812 15632
rect 9956 15580 10008 15632
rect 11428 15580 11480 15632
rect 16488 15691 16540 15700
rect 16488 15657 16497 15691
rect 16497 15657 16531 15691
rect 16531 15657 16540 15691
rect 16488 15648 16540 15657
rect 17500 15648 17552 15700
rect 19248 15648 19300 15700
rect 2044 15512 2096 15564
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 2688 15512 2740 15521
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 4252 15444 4304 15496
rect 6276 15512 6328 15564
rect 7748 15512 7800 15564
rect 8484 15512 8536 15564
rect 10048 15512 10100 15564
rect 10232 15512 10284 15564
rect 12440 15580 12492 15632
rect 17592 15580 17644 15632
rect 19064 15580 19116 15632
rect 11888 15512 11940 15564
rect 12624 15512 12676 15564
rect 13176 15555 13228 15564
rect 13176 15521 13185 15555
rect 13185 15521 13219 15555
rect 13219 15521 13228 15555
rect 13176 15512 13228 15521
rect 14556 15512 14608 15564
rect 11612 15444 11664 15496
rect 13268 15487 13320 15496
rect 3516 15419 3568 15428
rect 3516 15385 3525 15419
rect 3525 15385 3559 15419
rect 3559 15385 3568 15419
rect 3516 15376 3568 15385
rect 5356 15376 5408 15428
rect 7564 15419 7616 15428
rect 5632 15308 5684 15360
rect 7564 15385 7573 15419
rect 7573 15385 7607 15419
rect 7607 15385 7616 15419
rect 7564 15376 7616 15385
rect 12532 15376 12584 15428
rect 11980 15308 12032 15360
rect 12072 15308 12124 15360
rect 12256 15308 12308 15360
rect 12624 15308 12676 15360
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 15936 15444 15988 15496
rect 14280 15376 14332 15428
rect 13084 15308 13136 15360
rect 16672 15376 16724 15428
rect 16856 15444 16908 15496
rect 18788 15512 18840 15564
rect 19340 15555 19392 15564
rect 19340 15521 19349 15555
rect 19349 15521 19383 15555
rect 19383 15521 19392 15555
rect 19340 15512 19392 15521
rect 19616 15512 19668 15564
rect 17224 15444 17276 15496
rect 19248 15444 19300 15496
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 19524 15487 19576 15496
rect 19524 15453 19533 15487
rect 19533 15453 19567 15487
rect 19567 15453 19576 15487
rect 19524 15444 19576 15453
rect 16580 15308 16632 15360
rect 19156 15376 19208 15428
rect 20260 15444 20312 15496
rect 20076 15308 20128 15360
rect 20352 15308 20404 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2688 15104 2740 15156
rect 6276 15147 6328 15156
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 7380 15104 7432 15156
rect 11704 15104 11756 15156
rect 14556 15147 14608 15156
rect 1952 15079 2004 15088
rect 1952 15045 1961 15079
rect 1961 15045 1995 15079
rect 1995 15045 2004 15079
rect 1952 15036 2004 15045
rect 6184 15036 6236 15088
rect 3056 15011 3108 15020
rect 3056 14977 3065 15011
rect 3065 14977 3099 15011
rect 3099 14977 3108 15011
rect 3056 14968 3108 14977
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 5356 14968 5408 15020
rect 9220 15036 9272 15088
rect 7012 14968 7064 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 7748 14968 7800 15020
rect 8576 14968 8628 15020
rect 11152 15036 11204 15088
rect 13084 15036 13136 15088
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 17224 15079 17276 15088
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 12256 14968 12308 15020
rect 14556 14968 14608 15020
rect 17224 15045 17233 15079
rect 17233 15045 17267 15079
rect 17267 15045 17276 15079
rect 17224 15036 17276 15045
rect 18880 15036 18932 15088
rect 15844 15011 15896 15020
rect 15844 14977 15853 15011
rect 15853 14977 15887 15011
rect 15887 14977 15896 15011
rect 15844 14968 15896 14977
rect 2412 14900 2464 14952
rect 6368 14900 6420 14952
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 7196 14900 7248 14952
rect 8208 14900 8260 14952
rect 12440 14900 12492 14952
rect 8484 14832 8536 14884
rect 3700 14764 3752 14816
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 12716 14900 12768 14952
rect 14004 14832 14056 14884
rect 9956 14807 10008 14816
rect 9956 14773 9965 14807
rect 9965 14773 9999 14807
rect 9999 14773 10008 14807
rect 9956 14764 10008 14773
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 16764 14832 16816 14884
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 15476 14764 15528 14816
rect 17868 14832 17920 14884
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 18604 14900 18656 14952
rect 18696 14900 18748 14952
rect 20168 14832 20220 14884
rect 17500 14807 17552 14816
rect 17500 14773 17509 14807
rect 17509 14773 17543 14807
rect 17543 14773 17552 14807
rect 17500 14764 17552 14773
rect 19524 14764 19576 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 2872 14560 2924 14612
rect 204 14492 256 14544
rect 5172 14492 5224 14544
rect 1952 14424 2004 14476
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 3424 14424 3476 14476
rect 1400 14356 1452 14408
rect 3976 14356 4028 14408
rect 1768 14288 1820 14340
rect 2504 14288 2556 14340
rect 5448 14331 5500 14340
rect 5448 14297 5457 14331
rect 5457 14297 5491 14331
rect 5491 14297 5500 14331
rect 5448 14288 5500 14297
rect 4252 14220 4304 14272
rect 6276 14560 6328 14612
rect 7564 14492 7616 14544
rect 9312 14560 9364 14612
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 9956 14560 10008 14612
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 16304 14560 16356 14612
rect 16764 14603 16816 14612
rect 16764 14569 16773 14603
rect 16773 14569 16807 14603
rect 16807 14569 16816 14603
rect 16764 14560 16816 14569
rect 19248 14603 19300 14612
rect 10416 14492 10468 14544
rect 6460 14424 6512 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 9588 14356 9640 14408
rect 10600 14356 10652 14408
rect 8852 14288 8904 14340
rect 11980 14492 12032 14544
rect 13728 14492 13780 14544
rect 15476 14492 15528 14544
rect 16488 14492 16540 14544
rect 19248 14569 19257 14603
rect 19257 14569 19291 14603
rect 19291 14569 19300 14603
rect 19248 14560 19300 14569
rect 19340 14560 19392 14612
rect 20260 14560 20312 14612
rect 17316 14535 17368 14544
rect 17316 14501 17325 14535
rect 17325 14501 17359 14535
rect 17359 14501 17368 14535
rect 17316 14492 17368 14501
rect 11152 14467 11204 14476
rect 11152 14433 11186 14467
rect 11186 14433 11204 14467
rect 11152 14424 11204 14433
rect 11612 14424 11664 14476
rect 12256 14424 12308 14476
rect 14648 14467 14700 14476
rect 12624 14399 12676 14408
rect 6920 14220 6972 14272
rect 7380 14220 7432 14272
rect 8208 14220 8260 14272
rect 10324 14220 10376 14272
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 14648 14433 14657 14467
rect 14657 14433 14691 14467
rect 14691 14433 14700 14467
rect 14648 14424 14700 14433
rect 15936 14424 15988 14476
rect 15016 14356 15068 14408
rect 16948 14424 17000 14476
rect 18696 14492 18748 14544
rect 18880 14492 18932 14544
rect 20076 14535 20128 14544
rect 20076 14501 20085 14535
rect 20085 14501 20119 14535
rect 20119 14501 20128 14535
rect 20076 14492 20128 14501
rect 17224 14356 17276 14408
rect 18512 14424 18564 14476
rect 18604 14424 18656 14476
rect 20260 14424 20312 14476
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 11152 14220 11204 14272
rect 14004 14331 14056 14340
rect 14004 14297 14013 14331
rect 14013 14297 14047 14331
rect 14047 14297 14056 14331
rect 14004 14288 14056 14297
rect 17868 14220 17920 14272
rect 20536 14288 20588 14340
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 5448 14016 5500 14068
rect 3332 13880 3384 13932
rect 4712 13923 4764 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 2044 13812 2096 13864
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 5264 13812 5316 13864
rect 7196 14016 7248 14068
rect 8484 14016 8536 14068
rect 8852 14016 8904 14068
rect 9864 14016 9916 14068
rect 10600 14016 10652 14068
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 12440 14016 12492 14025
rect 15200 14016 15252 14068
rect 15936 14016 15988 14068
rect 16948 14016 17000 14068
rect 19432 14016 19484 14068
rect 7012 13948 7064 14000
rect 7748 13948 7800 14000
rect 11520 13948 11572 14000
rect 11888 13948 11940 14000
rect 12256 13948 12308 14000
rect 7564 13880 7616 13932
rect 9864 13880 9916 13932
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 3608 13744 3660 13796
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 4068 13676 4120 13728
rect 4988 13676 5040 13728
rect 9128 13812 9180 13864
rect 11980 13880 12032 13932
rect 13176 13948 13228 14000
rect 9680 13744 9732 13796
rect 10048 13744 10100 13796
rect 12256 13812 12308 13864
rect 12808 13812 12860 13864
rect 13176 13812 13228 13864
rect 14004 13880 14056 13932
rect 15016 13880 15068 13932
rect 10508 13787 10560 13796
rect 6736 13676 6788 13728
rect 7196 13676 7248 13728
rect 10508 13753 10542 13787
rect 10542 13753 10560 13787
rect 10508 13744 10560 13753
rect 10600 13744 10652 13796
rect 16580 13880 16632 13932
rect 16764 13880 16816 13932
rect 17132 13880 17184 13932
rect 17408 13880 17460 13932
rect 18696 13948 18748 14000
rect 16304 13812 16356 13864
rect 17960 13812 18012 13864
rect 19340 13812 19392 13864
rect 20168 13880 20220 13932
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 11796 13676 11848 13728
rect 13820 13676 13872 13728
rect 14188 13719 14240 13728
rect 14188 13685 14197 13719
rect 14197 13685 14231 13719
rect 14231 13685 14240 13719
rect 14188 13676 14240 13685
rect 16212 13744 16264 13796
rect 19800 13744 19852 13796
rect 15108 13719 15160 13728
rect 15108 13685 15117 13719
rect 15117 13685 15151 13719
rect 15151 13685 15160 13719
rect 15108 13676 15160 13685
rect 15200 13719 15252 13728
rect 15200 13685 15209 13719
rect 15209 13685 15243 13719
rect 15243 13685 15252 13719
rect 15200 13676 15252 13685
rect 18052 13676 18104 13728
rect 19248 13676 19300 13728
rect 19432 13676 19484 13728
rect 20352 13719 20404 13728
rect 20352 13685 20361 13719
rect 20361 13685 20395 13719
rect 20395 13685 20404 13719
rect 20352 13676 20404 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 3424 13472 3476 13524
rect 3608 13515 3660 13524
rect 3608 13481 3617 13515
rect 3617 13481 3651 13515
rect 3651 13481 3660 13515
rect 3608 13472 3660 13481
rect 4068 13515 4120 13524
rect 4068 13481 4077 13515
rect 4077 13481 4111 13515
rect 4111 13481 4120 13515
rect 4068 13472 4120 13481
rect 5264 13472 5316 13524
rect 7196 13472 7248 13524
rect 10232 13515 10284 13524
rect 4252 13404 4304 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 2044 13379 2096 13388
rect 2044 13345 2078 13379
rect 2078 13345 2096 13379
rect 2044 13336 2096 13345
rect 2596 13336 2648 13388
rect 3516 13336 3568 13388
rect 3884 13336 3936 13388
rect 9956 13404 10008 13456
rect 10232 13481 10241 13515
rect 10241 13481 10275 13515
rect 10275 13481 10284 13515
rect 10232 13472 10284 13481
rect 10600 13515 10652 13524
rect 10600 13481 10609 13515
rect 10609 13481 10643 13515
rect 10643 13481 10652 13515
rect 10600 13472 10652 13481
rect 11888 13472 11940 13524
rect 12440 13472 12492 13524
rect 11520 13404 11572 13456
rect 4712 13268 4764 13320
rect 3792 13200 3844 13252
rect 4068 13200 4120 13252
rect 9588 13336 9640 13388
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 6644 13311 6696 13320
rect 3608 13132 3660 13184
rect 5356 13200 5408 13252
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 7012 13268 7064 13320
rect 8576 13268 8628 13320
rect 12440 13336 12492 13388
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 13084 13404 13136 13456
rect 15384 13404 15436 13456
rect 16304 13472 16356 13524
rect 17500 13472 17552 13524
rect 17684 13472 17736 13524
rect 18512 13515 18564 13524
rect 18052 13404 18104 13456
rect 13268 13336 13320 13388
rect 14280 13336 14332 13388
rect 15292 13379 15344 13388
rect 10508 13268 10560 13320
rect 11980 13268 12032 13320
rect 12256 13268 12308 13320
rect 13452 13268 13504 13320
rect 12532 13200 12584 13252
rect 12808 13200 12860 13252
rect 8024 13132 8076 13184
rect 13360 13132 13412 13184
rect 13636 13268 13688 13320
rect 14004 13311 14056 13320
rect 14004 13277 14013 13311
rect 14013 13277 14047 13311
rect 14047 13277 14056 13311
rect 14004 13268 14056 13277
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 15936 13336 15988 13388
rect 16120 13336 16172 13388
rect 16212 13268 16264 13320
rect 16488 13336 16540 13388
rect 17224 13336 17276 13388
rect 17684 13336 17736 13388
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 18788 13515 18840 13524
rect 18788 13481 18797 13515
rect 18797 13481 18831 13515
rect 18831 13481 18840 13515
rect 18788 13472 18840 13481
rect 18880 13472 18932 13524
rect 20260 13515 20312 13524
rect 18420 13336 18472 13388
rect 20260 13481 20269 13515
rect 20269 13481 20303 13515
rect 20303 13481 20312 13515
rect 20260 13472 20312 13481
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 19432 13268 19484 13320
rect 17040 13200 17092 13252
rect 18788 13200 18840 13252
rect 13636 13132 13688 13184
rect 18604 13132 18656 13184
rect 18880 13132 18932 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 4160 12928 4212 12980
rect 4804 12928 4856 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 6644 12928 6696 12980
rect 8576 12928 8628 12980
rect 4344 12860 4396 12912
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 3240 12792 3292 12844
rect 4436 12792 4488 12844
rect 5356 12792 5408 12844
rect 7196 12792 7248 12844
rect 8024 12792 8076 12844
rect 9680 12928 9732 12980
rect 14188 12928 14240 12980
rect 14280 12928 14332 12980
rect 15108 12928 15160 12980
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 12716 12860 12768 12912
rect 12900 12860 12952 12912
rect 13084 12860 13136 12912
rect 11796 12835 11848 12844
rect 3884 12724 3936 12776
rect 3976 12724 4028 12776
rect 4252 12767 4304 12776
rect 4252 12733 4261 12767
rect 4261 12733 4295 12767
rect 4295 12733 4304 12767
rect 4252 12724 4304 12733
rect 7288 12724 7340 12776
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 3332 12699 3384 12708
rect 3332 12665 3341 12699
rect 3341 12665 3375 12699
rect 3375 12665 3384 12699
rect 3332 12656 3384 12665
rect 3700 12656 3752 12708
rect 4804 12656 4856 12708
rect 4896 12656 4948 12708
rect 5356 12699 5408 12708
rect 5356 12665 5365 12699
rect 5365 12665 5399 12699
rect 5399 12665 5408 12699
rect 5356 12656 5408 12665
rect 10876 12724 10928 12776
rect 8760 12656 8812 12708
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 11336 12724 11388 12776
rect 12256 12792 12308 12844
rect 12624 12792 12676 12844
rect 15384 12860 15436 12912
rect 15660 12860 15712 12912
rect 15016 12792 15068 12844
rect 15844 12792 15896 12844
rect 17224 12928 17276 12980
rect 17684 12971 17736 12980
rect 17684 12937 17693 12971
rect 17693 12937 17727 12971
rect 17727 12937 17736 12971
rect 17684 12928 17736 12937
rect 17960 12928 18012 12980
rect 18512 12928 18564 12980
rect 19984 12928 20036 12980
rect 18788 12860 18840 12912
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 15200 12724 15252 12776
rect 15384 12724 15436 12776
rect 18880 12724 18932 12776
rect 19432 12724 19484 12776
rect 6000 12588 6052 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 7656 12631 7708 12640
rect 7656 12597 7665 12631
rect 7665 12597 7699 12631
rect 7699 12597 7708 12631
rect 7656 12588 7708 12597
rect 10324 12631 10376 12640
rect 10324 12597 10333 12631
rect 10333 12597 10367 12631
rect 10367 12597 10376 12631
rect 10324 12588 10376 12597
rect 10692 12631 10744 12640
rect 10692 12597 10701 12631
rect 10701 12597 10735 12631
rect 10735 12597 10744 12631
rect 10692 12588 10744 12597
rect 10876 12588 10928 12640
rect 12348 12656 12400 12708
rect 13912 12656 13964 12708
rect 13636 12588 13688 12640
rect 15384 12631 15436 12640
rect 15384 12597 15393 12631
rect 15393 12597 15427 12631
rect 15427 12597 15436 12631
rect 15384 12588 15436 12597
rect 16304 12656 16356 12708
rect 17960 12656 18012 12708
rect 20076 12656 20128 12708
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2044 12384 2096 12436
rect 4344 12384 4396 12436
rect 5356 12384 5408 12436
rect 5540 12384 5592 12436
rect 5908 12384 5960 12436
rect 7656 12384 7708 12436
rect 10324 12384 10376 12436
rect 10692 12384 10744 12436
rect 10968 12384 11020 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 12808 12384 12860 12436
rect 13360 12427 13412 12436
rect 13360 12393 13369 12427
rect 13369 12393 13403 12427
rect 13403 12393 13412 12427
rect 13360 12384 13412 12393
rect 18788 12427 18840 12436
rect 3516 12359 3568 12368
rect 3516 12325 3525 12359
rect 3525 12325 3559 12359
rect 3559 12325 3568 12359
rect 3516 12316 3568 12325
rect 7196 12316 7248 12368
rect 7748 12316 7800 12368
rect 8668 12316 8720 12368
rect 12072 12316 12124 12368
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 19616 12384 19668 12436
rect 20168 12384 20220 12436
rect 17868 12316 17920 12368
rect 2596 12248 2648 12300
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 4252 12248 4304 12300
rect 5080 12248 5132 12300
rect 5264 12248 5316 12300
rect 5908 12248 5960 12300
rect 10968 12248 11020 12300
rect 11152 12248 11204 12300
rect 11336 12248 11388 12300
rect 11796 12248 11848 12300
rect 14280 12291 14332 12300
rect 14280 12257 14289 12291
rect 14289 12257 14323 12291
rect 14323 12257 14332 12291
rect 14280 12248 14332 12257
rect 15844 12248 15896 12300
rect 16028 12291 16080 12300
rect 16028 12257 16062 12291
rect 16062 12257 16080 12291
rect 16028 12248 16080 12257
rect 17224 12248 17276 12300
rect 19708 12248 19760 12300
rect 3700 12180 3752 12232
rect 4436 12180 4488 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 8760 12180 8812 12232
rect 6092 12112 6144 12164
rect 10508 12180 10560 12232
rect 13360 12180 13412 12232
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 12532 12112 12584 12164
rect 3792 12044 3844 12096
rect 7564 12087 7616 12096
rect 7564 12053 7573 12087
rect 7573 12053 7607 12087
rect 7607 12053 7616 12087
rect 7564 12044 7616 12053
rect 8300 12044 8352 12096
rect 8484 12044 8536 12096
rect 12900 12044 12952 12096
rect 13452 12044 13504 12096
rect 19432 12180 19484 12232
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 18972 12112 19024 12164
rect 19892 12112 19944 12164
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 2320 11840 2372 11892
rect 3240 11772 3292 11824
rect 2044 11704 2096 11756
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 5724 11815 5776 11824
rect 5724 11781 5733 11815
rect 5733 11781 5767 11815
rect 5767 11781 5776 11815
rect 5724 11772 5776 11781
rect 6092 11772 6144 11824
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 1952 11568 2004 11620
rect 3608 11568 3660 11620
rect 3976 11568 4028 11620
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 3792 11500 3844 11552
rect 5908 11636 5960 11688
rect 7564 11704 7616 11756
rect 8208 11704 8260 11756
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7104 11500 7156 11552
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 9036 11500 9088 11552
rect 12808 11840 12860 11892
rect 16028 11883 16080 11892
rect 16028 11849 16037 11883
rect 16037 11849 16071 11883
rect 16071 11849 16080 11883
rect 16028 11840 16080 11849
rect 17776 11840 17828 11892
rect 17960 11840 18012 11892
rect 20168 11840 20220 11892
rect 20996 11883 21048 11892
rect 20996 11849 21005 11883
rect 21005 11849 21039 11883
rect 21039 11849 21048 11883
rect 20996 11840 21048 11849
rect 11796 11772 11848 11824
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 9680 11704 9732 11756
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 13360 11704 13412 11756
rect 14280 11704 14332 11756
rect 18788 11704 18840 11756
rect 10508 11636 10560 11688
rect 10968 11636 11020 11688
rect 12716 11636 12768 11688
rect 14556 11636 14608 11688
rect 15660 11636 15712 11688
rect 17132 11636 17184 11688
rect 18696 11636 18748 11688
rect 19064 11636 19116 11688
rect 20812 11679 20864 11688
rect 20812 11645 20821 11679
rect 20821 11645 20855 11679
rect 20855 11645 20864 11679
rect 20812 11636 20864 11645
rect 9312 11611 9364 11620
rect 9312 11577 9321 11611
rect 9321 11577 9355 11611
rect 9355 11577 9364 11611
rect 9312 11568 9364 11577
rect 9496 11568 9548 11620
rect 15108 11568 15160 11620
rect 15292 11568 15344 11620
rect 19892 11568 19944 11620
rect 9404 11500 9456 11552
rect 10784 11500 10836 11552
rect 13176 11500 13228 11552
rect 13728 11500 13780 11552
rect 15384 11500 15436 11552
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2228 11296 2280 11348
rect 4252 11296 4304 11348
rect 4712 11296 4764 11348
rect 6552 11296 6604 11348
rect 8668 11339 8720 11348
rect 2504 11228 2556 11280
rect 5724 11228 5776 11280
rect 8300 11228 8352 11280
rect 6920 11203 6972 11212
rect 6920 11169 6954 11203
rect 6954 11169 6972 11203
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 8852 11296 8904 11348
rect 10600 11296 10652 11348
rect 10968 11296 11020 11348
rect 13636 11296 13688 11348
rect 14372 11296 14424 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16580 11296 16632 11348
rect 16948 11296 17000 11348
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 19248 11296 19300 11348
rect 19708 11339 19760 11348
rect 19708 11305 19717 11339
rect 19717 11305 19751 11339
rect 19751 11305 19760 11339
rect 19708 11296 19760 11305
rect 11704 11228 11756 11280
rect 12624 11271 12676 11280
rect 12624 11237 12658 11271
rect 12658 11237 12676 11271
rect 12624 11228 12676 11237
rect 14096 11228 14148 11280
rect 16120 11228 16172 11280
rect 20168 11228 20220 11280
rect 6920 11160 6972 11169
rect 2228 11092 2280 11144
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 3700 11092 3752 11144
rect 2136 11024 2188 11076
rect 3516 11024 3568 11076
rect 3792 11024 3844 11076
rect 5908 11092 5960 11144
rect 9128 11160 9180 11212
rect 12440 11160 12492 11212
rect 15200 11160 15252 11212
rect 6368 11067 6420 11076
rect 6368 11033 6377 11067
rect 6377 11033 6411 11067
rect 6411 11033 6420 11067
rect 6368 11024 6420 11033
rect 8484 11024 8536 11076
rect 9404 11024 9456 11076
rect 4804 10956 4856 11008
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 9588 11092 9640 11144
rect 12256 11092 12308 11144
rect 14924 11092 14976 11144
rect 15660 11024 15712 11076
rect 16212 11024 16264 11076
rect 16764 11024 16816 11076
rect 17776 11092 17828 11144
rect 18604 11160 18656 11212
rect 20076 11203 20128 11212
rect 20076 11169 20085 11203
rect 20085 11169 20119 11203
rect 20119 11169 20128 11203
rect 20076 11160 20128 11169
rect 19984 11092 20036 11144
rect 19892 11024 19944 11076
rect 11152 10956 11204 11008
rect 13544 10956 13596 11008
rect 16856 10956 16908 11008
rect 16948 10956 17000 11008
rect 17960 10956 18012 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 3884 10795 3936 10804
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 4068 10752 4120 10804
rect 10968 10752 11020 10804
rect 4620 10684 4672 10736
rect 9588 10684 9640 10736
rect 11612 10684 11664 10736
rect 1584 10616 1636 10668
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 3240 10616 3292 10668
rect 5908 10616 5960 10668
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8852 10616 8904 10668
rect 8944 10616 8996 10668
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 2872 10548 2924 10600
rect 3148 10548 3200 10600
rect 6368 10548 6420 10600
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 3700 10480 3752 10532
rect 5816 10480 5868 10532
rect 10968 10480 11020 10532
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 2596 10412 2648 10464
rect 4804 10412 4856 10464
rect 5356 10412 5408 10464
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6092 10455 6144 10464
rect 6092 10421 6101 10455
rect 6101 10421 6135 10455
rect 6135 10421 6144 10455
rect 6092 10412 6144 10421
rect 6552 10412 6604 10464
rect 7196 10412 7248 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 8852 10455 8904 10464
rect 7288 10412 7340 10421
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 8944 10412 8996 10464
rect 13544 10616 13596 10668
rect 14096 10616 14148 10668
rect 14556 10616 14608 10668
rect 14648 10616 14700 10668
rect 15752 10752 15804 10804
rect 16212 10795 16264 10804
rect 16212 10761 16221 10795
rect 16221 10761 16255 10795
rect 16255 10761 16264 10795
rect 16212 10752 16264 10761
rect 16672 10752 16724 10804
rect 18880 10752 18932 10804
rect 19156 10752 19208 10804
rect 19892 10795 19944 10804
rect 16856 10684 16908 10736
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 16948 10616 17000 10625
rect 11152 10548 11204 10600
rect 11520 10591 11572 10600
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 11704 10480 11756 10532
rect 14372 10480 14424 10532
rect 14924 10548 14976 10600
rect 16764 10548 16816 10600
rect 17960 10548 18012 10600
rect 18420 10548 18472 10600
rect 19892 10761 19901 10795
rect 19901 10761 19935 10795
rect 19935 10761 19944 10795
rect 19892 10752 19944 10761
rect 20076 10752 20128 10804
rect 20536 10616 20588 10668
rect 17408 10480 17460 10532
rect 18604 10480 18656 10532
rect 11152 10412 11204 10421
rect 12716 10412 12768 10464
rect 13176 10412 13228 10464
rect 13728 10412 13780 10464
rect 14096 10412 14148 10464
rect 16304 10412 16356 10464
rect 18328 10412 18380 10464
rect 18420 10412 18472 10464
rect 19064 10412 19116 10464
rect 19248 10412 19300 10464
rect 19708 10412 19760 10464
rect 20720 10455 20772 10464
rect 20720 10421 20729 10455
rect 20729 10421 20763 10455
rect 20763 10421 20772 10455
rect 20720 10412 20772 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1676 10208 1728 10260
rect 6736 10208 6788 10260
rect 7196 10251 7248 10260
rect 7196 10217 7205 10251
rect 7205 10217 7239 10251
rect 7239 10217 7248 10251
rect 7196 10208 7248 10217
rect 8300 10208 8352 10260
rect 9680 10208 9732 10260
rect 10968 10208 11020 10260
rect 13268 10208 13320 10260
rect 13912 10208 13964 10260
rect 15016 10208 15068 10260
rect 16120 10208 16172 10260
rect 17776 10251 17828 10260
rect 17776 10217 17785 10251
rect 17785 10217 17819 10251
rect 17819 10217 17828 10251
rect 17776 10208 17828 10217
rect 20720 10208 20772 10260
rect 3516 10140 3568 10192
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 3332 10072 3384 10081
rect 3884 10072 3936 10124
rect 4712 10140 4764 10192
rect 6368 10140 6420 10192
rect 4620 10072 4672 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 3700 10004 3752 10056
rect 8852 10072 8904 10124
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 7564 10004 7616 10056
rect 8208 10004 8260 10056
rect 8576 10004 8628 10056
rect 10692 10140 10744 10192
rect 9956 10115 10008 10124
rect 9956 10081 9990 10115
rect 9990 10081 10008 10115
rect 9956 10072 10008 10081
rect 12624 10140 12676 10192
rect 1952 9979 2004 9988
rect 1952 9945 1961 9979
rect 1961 9945 1995 9979
rect 1995 9945 2004 9979
rect 1952 9936 2004 9945
rect 3976 9868 4028 9920
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 8668 9868 8720 9920
rect 11796 9868 11848 9920
rect 11980 9911 12032 9920
rect 11980 9877 11989 9911
rect 11989 9877 12023 9911
rect 12023 9877 12032 9911
rect 11980 9868 12032 9877
rect 12348 10004 12400 10056
rect 13268 10072 13320 10124
rect 12808 10004 12860 10056
rect 14464 10140 14516 10192
rect 14924 10140 14976 10192
rect 16580 10140 16632 10192
rect 18052 10140 18104 10192
rect 19708 10140 19760 10192
rect 19892 10140 19944 10192
rect 13636 10072 13688 10124
rect 15752 10072 15804 10124
rect 16212 10072 16264 10124
rect 17500 10072 17552 10124
rect 18328 10072 18380 10124
rect 18696 10072 18748 10124
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 14004 10004 14056 10056
rect 14648 10004 14700 10056
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 13912 9868 13964 9920
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 17316 9868 17368 9920
rect 19248 10004 19300 10056
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 19432 9979 19484 9988
rect 19432 9945 19441 9979
rect 19441 9945 19475 9979
rect 19475 9945 19484 9979
rect 19432 9936 19484 9945
rect 19064 9868 19116 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 4068 9664 4120 9716
rect 8208 9707 8260 9716
rect 1860 9639 1912 9648
rect 1860 9605 1869 9639
rect 1869 9605 1903 9639
rect 1903 9605 1912 9639
rect 1860 9596 1912 9605
rect 2228 9639 2280 9648
rect 2228 9605 2237 9639
rect 2237 9605 2271 9639
rect 2271 9605 2280 9639
rect 2228 9596 2280 9605
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 12532 9664 12584 9716
rect 13912 9664 13964 9716
rect 11336 9596 11388 9648
rect 3516 9528 3568 9580
rect 3700 9528 3752 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 4160 9460 4212 9512
rect 2780 9392 2832 9444
rect 12348 9528 12400 9580
rect 13636 9596 13688 9648
rect 13728 9596 13780 9648
rect 4620 9460 4672 9512
rect 5908 9460 5960 9512
rect 9772 9460 9824 9512
rect 11152 9460 11204 9512
rect 11244 9460 11296 9512
rect 13544 9528 13596 9580
rect 14096 9528 14148 9580
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 15568 9528 15620 9580
rect 14740 9460 14792 9512
rect 15292 9460 15344 9512
rect 16304 9460 16356 9512
rect 16488 9596 16540 9648
rect 18880 9664 18932 9716
rect 19248 9596 19300 9648
rect 19984 9639 20036 9648
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 19984 9605 19993 9639
rect 19993 9605 20027 9639
rect 20027 9605 20036 9639
rect 19984 9596 20036 9605
rect 20536 9571 20588 9580
rect 3240 9324 3292 9376
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 5540 9392 5592 9444
rect 4896 9324 4948 9376
rect 7012 9392 7064 9444
rect 8484 9392 8536 9444
rect 8944 9392 8996 9444
rect 9588 9392 9640 9444
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10784 9324 10836 9376
rect 11612 9324 11664 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 14096 9324 14148 9376
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 15936 9392 15988 9444
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 18512 9435 18564 9444
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16948 9367 17000 9376
rect 16212 9324 16264 9333
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 16948 9324 17000 9333
rect 18512 9401 18546 9435
rect 18546 9401 18564 9435
rect 18512 9392 18564 9401
rect 19432 9392 19484 9444
rect 18420 9324 18472 9376
rect 18696 9324 18748 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 3516 9120 3568 9172
rect 3700 9120 3752 9172
rect 7288 9120 7340 9172
rect 1676 9052 1728 9104
rect 4068 9052 4120 9104
rect 11336 9120 11388 9172
rect 12900 9120 12952 9172
rect 13268 9163 13320 9172
rect 13268 9129 13277 9163
rect 13277 9129 13311 9163
rect 13311 9129 13320 9163
rect 13268 9120 13320 9129
rect 7564 9095 7616 9104
rect 7564 9061 7598 9095
rect 7598 9061 7616 9095
rect 7564 9052 7616 9061
rect 10140 9052 10192 9104
rect 10324 9052 10376 9104
rect 11244 9052 11296 9104
rect 13820 9120 13872 9172
rect 14280 9120 14332 9172
rect 15476 9120 15528 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 14188 9052 14240 9104
rect 16948 9052 17000 9104
rect 1492 9027 1544 9036
rect 1492 8993 1501 9027
rect 1501 8993 1535 9027
rect 1535 8993 1544 9027
rect 1492 8984 1544 8993
rect 2136 8984 2188 9036
rect 3056 8984 3108 9036
rect 3884 8984 3936 9036
rect 3240 8916 3292 8968
rect 4804 8916 4856 8968
rect 7012 8984 7064 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 5816 8916 5868 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 12072 8984 12124 9036
rect 12256 8984 12308 9036
rect 12532 8984 12584 9036
rect 5632 8848 5684 8900
rect 4712 8780 4764 8832
rect 5908 8780 5960 8832
rect 10876 8916 10928 8968
rect 13268 8984 13320 9036
rect 13452 8916 13504 8968
rect 13820 8959 13872 8968
rect 13820 8925 13829 8959
rect 13829 8925 13863 8959
rect 13863 8925 13872 8959
rect 13820 8916 13872 8925
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 15936 8984 15988 9036
rect 16212 8984 16264 9036
rect 17408 8984 17460 9036
rect 17868 8984 17920 9036
rect 18788 8984 18840 9036
rect 19800 8984 19852 9036
rect 14188 8916 14240 8968
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 19248 8916 19300 8968
rect 13912 8848 13964 8900
rect 14556 8848 14608 8900
rect 17224 8848 17276 8900
rect 18696 8848 18748 8900
rect 19892 8848 19944 8900
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 9956 8780 10008 8832
rect 10968 8780 11020 8832
rect 12072 8780 12124 8832
rect 12440 8780 12492 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 5540 8576 5592 8628
rect 10324 8576 10376 8628
rect 3884 8440 3936 8492
rect 2136 8304 2188 8356
rect 4160 8304 4212 8356
rect 4988 8304 5040 8356
rect 9956 8440 10008 8492
rect 11980 8576 12032 8628
rect 10968 8508 11020 8560
rect 10784 8440 10836 8492
rect 12164 8440 12216 8492
rect 12532 8440 12584 8492
rect 15016 8576 15068 8628
rect 16304 8619 16356 8628
rect 5632 8304 5684 8356
rect 11152 8304 11204 8356
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 5172 8236 5224 8288
rect 11612 8304 11664 8356
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 18512 8576 18564 8628
rect 20628 8576 20680 8628
rect 17500 8440 17552 8492
rect 18604 8440 18656 8492
rect 14004 8304 14056 8356
rect 14556 8347 14608 8356
rect 14556 8313 14565 8347
rect 14565 8313 14599 8347
rect 14599 8313 14608 8347
rect 14556 8304 14608 8313
rect 15108 8304 15160 8356
rect 16672 8347 16724 8356
rect 16672 8313 16681 8347
rect 16681 8313 16715 8347
rect 16715 8313 16724 8347
rect 16672 8304 16724 8313
rect 11888 8236 11940 8288
rect 15200 8236 15252 8288
rect 16028 8279 16080 8288
rect 16028 8245 16037 8279
rect 16037 8245 16071 8279
rect 16071 8245 16080 8279
rect 16028 8236 16080 8245
rect 16764 8279 16816 8288
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 19340 8372 19392 8424
rect 20444 8304 20496 8356
rect 19248 8236 19300 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 1492 8032 1544 8084
rect 5080 8032 5132 8084
rect 5632 8032 5684 8084
rect 6000 8032 6052 8084
rect 10416 8032 10468 8084
rect 11152 8032 11204 8084
rect 12716 8032 12768 8084
rect 14280 8032 14332 8084
rect 14464 8032 14516 8084
rect 16672 8032 16724 8084
rect 4712 7964 4764 8016
rect 5724 7964 5776 8016
rect 9864 7964 9916 8016
rect 4160 7939 4212 7948
rect 4160 7905 4169 7939
rect 4169 7905 4203 7939
rect 4203 7905 4212 7939
rect 4160 7896 4212 7905
rect 5540 7896 5592 7948
rect 6092 7896 6144 7948
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 4068 7692 4120 7744
rect 10048 7760 10100 7812
rect 11796 7964 11848 8016
rect 12624 7964 12676 8016
rect 10968 7896 11020 7948
rect 11704 7896 11756 7948
rect 11980 7896 12032 7948
rect 14464 7939 14516 7948
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 14464 7896 14516 7905
rect 16028 7964 16080 8016
rect 19524 7964 19576 8016
rect 16856 7896 16908 7948
rect 17960 7896 18012 7948
rect 18512 7896 18564 7948
rect 18604 7896 18656 7948
rect 19064 7896 19116 7948
rect 12348 7828 12400 7880
rect 14556 7828 14608 7880
rect 15936 7828 15988 7880
rect 10876 7760 10928 7812
rect 12072 7760 12124 7812
rect 12532 7760 12584 7812
rect 17408 7803 17460 7812
rect 17408 7769 17417 7803
rect 17417 7769 17451 7803
rect 17451 7769 17460 7803
rect 20168 7828 20220 7880
rect 17408 7760 17460 7769
rect 11612 7692 11664 7744
rect 12256 7735 12308 7744
rect 12256 7701 12265 7735
rect 12265 7701 12299 7735
rect 12299 7701 12308 7735
rect 12256 7692 12308 7701
rect 12348 7692 12400 7744
rect 16948 7692 17000 7744
rect 20352 7735 20404 7744
rect 20352 7701 20361 7735
rect 20361 7701 20395 7735
rect 20395 7701 20404 7735
rect 20352 7692 20404 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 5172 7488 5224 7540
rect 10508 7488 10560 7540
rect 11704 7531 11756 7540
rect 940 7352 992 7404
rect 3608 7352 3660 7404
rect 5540 7420 5592 7472
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 12440 7488 12492 7540
rect 13176 7488 13228 7540
rect 15108 7488 15160 7540
rect 16764 7488 16816 7540
rect 17960 7488 18012 7540
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 12348 7420 12400 7472
rect 13912 7420 13964 7472
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 9680 7352 9732 7404
rect 4068 7216 4120 7268
rect 11888 7284 11940 7336
rect 10876 7216 10928 7268
rect 11060 7216 11112 7268
rect 12164 7284 12216 7336
rect 17408 7352 17460 7404
rect 18328 7352 18380 7404
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 15936 7284 15988 7336
rect 12256 7216 12308 7268
rect 13176 7216 13228 7268
rect 20812 7284 20864 7336
rect 20352 7216 20404 7268
rect 4252 7148 4304 7200
rect 4804 7148 4856 7200
rect 9864 7148 9916 7200
rect 11980 7148 12032 7200
rect 12532 7148 12584 7200
rect 15292 7148 15344 7200
rect 16580 7191 16632 7200
rect 16580 7157 16589 7191
rect 16589 7157 16623 7191
rect 16623 7157 16632 7191
rect 16580 7148 16632 7157
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 14464 6944 14516 6996
rect 15476 6944 15528 6996
rect 18604 6944 18656 6996
rect 20168 6987 20220 6996
rect 20168 6953 20177 6987
rect 20177 6953 20211 6987
rect 20211 6953 20220 6987
rect 20168 6944 20220 6953
rect 3976 6808 4028 6860
rect 11060 6808 11112 6860
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 13360 6876 13412 6928
rect 15476 6808 15528 6860
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 16396 6808 16448 6860
rect 18328 6876 18380 6928
rect 12256 6740 12308 6792
rect 4068 6672 4120 6724
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 11704 6672 11756 6724
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 14648 6783 14700 6792
rect 13728 6740 13780 6749
rect 14648 6749 14657 6783
rect 14657 6749 14691 6783
rect 14691 6749 14700 6783
rect 14648 6740 14700 6749
rect 15108 6740 15160 6792
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 16028 6740 16080 6792
rect 17040 6740 17092 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 20076 6740 20128 6792
rect 20444 6783 20496 6792
rect 20444 6749 20453 6783
rect 20453 6749 20487 6783
rect 20487 6749 20496 6783
rect 20444 6740 20496 6749
rect 16580 6672 16632 6724
rect 18512 6672 18564 6724
rect 19800 6715 19852 6724
rect 19800 6681 19809 6715
rect 19809 6681 19843 6715
rect 19843 6681 19852 6715
rect 19800 6672 19852 6681
rect 12440 6604 12492 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 11060 6400 11112 6452
rect 12532 6400 12584 6452
rect 14648 6400 14700 6452
rect 15200 6400 15252 6452
rect 15660 6400 15712 6452
rect 16672 6400 16724 6452
rect 20076 6443 20128 6452
rect 20076 6409 20085 6443
rect 20085 6409 20119 6443
rect 20119 6409 20128 6443
rect 20076 6400 20128 6409
rect 5448 6332 5500 6384
rect 17960 6332 18012 6384
rect 11704 6264 11756 6316
rect 11888 6264 11940 6316
rect 13728 6264 13780 6316
rect 15200 6264 15252 6316
rect 11152 6196 11204 6248
rect 10600 6128 10652 6180
rect 11980 6128 12032 6180
rect 13820 6128 13872 6180
rect 15936 6264 15988 6316
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 20352 6264 20404 6316
rect 16948 6196 17000 6248
rect 11428 6103 11480 6112
rect 11428 6069 11437 6103
rect 11437 6069 11471 6103
rect 11471 6069 11480 6103
rect 11428 6060 11480 6069
rect 15200 6103 15252 6112
rect 15200 6069 15209 6103
rect 15209 6069 15243 6103
rect 15243 6069 15252 6103
rect 15200 6060 15252 6069
rect 18052 6128 18104 6180
rect 16396 6060 16448 6112
rect 16856 6060 16908 6112
rect 19892 6103 19944 6112
rect 19892 6069 19901 6103
rect 19901 6069 19935 6103
rect 19935 6069 19944 6103
rect 19892 6060 19944 6069
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 11428 5856 11480 5908
rect 3148 5788 3200 5840
rect 19892 5856 19944 5908
rect 11796 5788 11848 5840
rect 11980 5788 12032 5840
rect 17960 5788 18012 5840
rect 4160 5720 4212 5772
rect 11888 5720 11940 5772
rect 15200 5720 15252 5772
rect 18144 5720 18196 5772
rect 10600 5652 10652 5704
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 11060 5652 11112 5704
rect 11980 5516 12032 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 11152 5312 11204 5364
rect 13820 5312 13872 5364
rect 18512 5312 18564 5364
rect 4068 5176 4120 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 17224 5108 17276 5160
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 4068 4088 4120 4140
rect 5356 4088 5408 4140
rect 12808 4088 12860 4140
rect 17960 4088 18012 4140
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 11060 3680 11112 3732
rect 11796 3680 11848 3732
rect 11152 3612 11204 3664
rect 8668 3476 8720 3528
rect 18972 3544 19024 3596
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 3332 2048 3384 2100
rect 4804 2048 4856 2100
rect 14096 2048 14148 2100
rect 18512 2048 18564 2100
rect 3148 688 3200 740
rect 4896 688 4948 740
rect 3332 280 3384 332
rect 5264 280 5316 332
<< metal2 >>
rect 202 22320 258 22800
rect 662 22320 718 22800
rect 1122 22320 1178 22800
rect 1582 22320 1638 22800
rect 2042 22320 2098 22800
rect 2502 22320 2558 22800
rect 2778 22536 2834 22545
rect 2778 22471 2834 22480
rect 216 14550 244 22320
rect 676 18086 704 22320
rect 1136 18698 1164 22320
rect 1596 19009 1624 22320
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1950 19272 2006 19281
rect 2056 19258 2084 22320
rect 2516 19802 2544 22320
rect 2792 20058 2820 22471
rect 3054 22320 3110 22800
rect 3514 22320 3570 22800
rect 3974 22320 4030 22800
rect 4434 22320 4490 22800
rect 4894 22320 4950 22800
rect 5354 22320 5410 22800
rect 5906 22320 5962 22800
rect 6366 22320 6422 22800
rect 6826 22320 6882 22800
rect 7286 22320 7342 22800
rect 7746 22320 7802 22800
rect 8206 22320 8262 22800
rect 8758 22320 8814 22800
rect 9218 22320 9274 22800
rect 9678 22320 9734 22800
rect 10138 22320 10194 22800
rect 10598 22320 10654 22800
rect 11058 22320 11114 22800
rect 11610 22320 11666 22800
rect 12070 22320 12126 22800
rect 12530 22320 12586 22800
rect 12990 22320 13046 22800
rect 13450 22320 13506 22800
rect 13910 22320 13966 22800
rect 14462 22320 14518 22800
rect 14922 22320 14978 22800
rect 15382 22320 15438 22800
rect 15842 22320 15898 22800
rect 16302 22320 16358 22800
rect 16762 22320 16818 22800
rect 17314 22320 17370 22800
rect 17774 22320 17830 22800
rect 18234 22320 18290 22800
rect 18694 22320 18750 22800
rect 19154 22320 19210 22800
rect 19614 22320 19670 22800
rect 20166 22320 20222 22800
rect 20626 22320 20682 22800
rect 20718 22536 20774 22545
rect 20718 22471 20774 22480
rect 2962 22128 3018 22137
rect 2962 22063 3018 22072
rect 2870 21176 2926 21185
rect 2870 21111 2926 21120
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2516 19774 2728 19802
rect 2504 19712 2556 19718
rect 2504 19654 2556 19660
rect 2134 19272 2190 19281
rect 2056 19230 2134 19258
rect 1950 19207 2006 19216
rect 2134 19207 2190 19216
rect 1582 19000 1638 19009
rect 1964 18970 1992 19207
rect 1582 18935 1638 18944
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2516 18873 2544 19654
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2608 18902 2636 19246
rect 2596 18896 2648 18902
rect 1766 18864 1822 18873
rect 2502 18864 2558 18873
rect 1766 18799 1822 18808
rect 2228 18828 2280 18834
rect 1124 18692 1176 18698
rect 1124 18634 1176 18640
rect 1780 18426 1808 18799
rect 2228 18770 2280 18776
rect 2320 18828 2372 18834
rect 2596 18838 2648 18844
rect 2502 18799 2558 18808
rect 2320 18770 2372 18776
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 2240 18222 2268 18770
rect 2332 18426 2360 18770
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 664 18080 716 18086
rect 664 18022 716 18028
rect 1596 16697 1624 18158
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2134 17776 2190 17785
rect 2134 17711 2136 17720
rect 2188 17711 2190 17720
rect 2136 17682 2188 17688
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 1780 17377 1808 17478
rect 1766 17368 1822 17377
rect 1766 17303 1822 17312
rect 2516 17202 2544 17478
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 1952 16992 2004 16998
rect 1950 16960 1952 16969
rect 2004 16960 2006 16969
rect 1950 16895 2006 16904
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1952 16584 2004 16590
rect 1582 16552 1638 16561
rect 1952 16526 2004 16532
rect 1582 16487 1584 16496
rect 1636 16487 1638 16496
rect 1584 16458 1636 16464
rect 1964 16114 1992 16526
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 2516 16046 2544 17138
rect 2608 16998 2636 18022
rect 2700 17814 2728 19774
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 2792 19281 2820 19382
rect 2778 19272 2834 19281
rect 2778 19207 2834 19216
rect 2884 19174 2912 21111
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2976 18970 3004 22063
rect 3068 19174 3096 22320
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3068 18426 3096 18906
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3054 18320 3110 18329
rect 3054 18255 3110 18264
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2778 17912 2834 17921
rect 2778 17847 2834 17856
rect 2688 17808 2740 17814
rect 2688 17750 2740 17756
rect 2792 17338 2820 17847
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2976 17184 3004 18158
rect 3068 17882 3096 18255
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2792 17156 3004 17184
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 204 14544 256 14550
rect 204 14486 256 14492
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13870 1440 14350
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1504 11393 1532 15846
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1964 15609 1992 15642
rect 1950 15600 2006 15609
rect 2056 15570 2084 15914
rect 2332 15706 2360 15982
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 1950 15535 2006 15544
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 1952 15088 2004 15094
rect 1950 15056 1952 15065
rect 2004 15056 2006 15065
rect 1950 14991 2006 15000
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 1582 14648 1638 14657
rect 1582 14583 1638 14592
rect 1596 14074 1624 14583
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1780 13394 1808 14282
rect 1858 14104 1914 14113
rect 1964 14074 1992 14418
rect 1858 14039 1914 14048
rect 1952 14068 2004 14074
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1490 11384 1546 11393
rect 1490 11319 1546 11328
rect 1596 10674 1624 12174
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10266 1716 10406
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1872 9654 1900 14039
rect 1952 14010 2004 14016
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2056 13394 2084 13806
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2056 12442 2084 13330
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 2056 11762 2084 12378
rect 2332 11898 2360 13670
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2424 11665 2452 14894
rect 2516 14346 2544 15982
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2700 15162 2728 15506
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2410 11656 2466 11665
rect 1952 11620 2004 11626
rect 2410 11591 2466 11600
rect 1952 11562 2004 11568
rect 1964 9994 1992 11562
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11354 2268 11494
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2516 11286 2544 12786
rect 2608 12306 2636 13330
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2608 11150 2636 12242
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2148 10674 2176 11018
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9110 1716 9454
rect 1676 9104 1728 9110
rect 1676 9046 1728 9052
rect 2148 9042 2176 10610
rect 2240 9654 2268 11086
rect 2608 10470 2636 11086
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 10062 2636 10406
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2228 9648 2280 9654
rect 2792 9625 2820 17156
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2976 16454 3004 17002
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2976 15502 3004 16390
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3068 15026 3096 16594
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3160 14906 3188 19858
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 2976 14878 3188 14906
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 14618 2912 14758
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2228 9590 2280 9596
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2884 9466 2912 10542
rect 2792 9450 2912 9466
rect 2780 9444 2912 9450
rect 2832 9438 2912 9444
rect 2780 9386 2832 9392
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 1504 8090 1532 8978
rect 2148 8362 2176 8978
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 952 1057 980 7346
rect 2792 2009 2820 9386
rect 2976 5817 3004 14878
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3160 10606 3188 14418
rect 3252 13297 3280 19790
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 3344 15910 3372 19722
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 19145 3464 19654
rect 3422 19136 3478 19145
rect 3422 19071 3478 19080
rect 3424 18760 3476 18766
rect 3422 18728 3424 18737
rect 3476 18728 3478 18737
rect 3422 18663 3478 18672
rect 3528 17066 3556 22320
rect 3882 21584 3938 21593
rect 3882 21519 3938 21528
rect 3698 20632 3754 20641
rect 3698 20567 3754 20576
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3620 19281 3648 19654
rect 3712 19514 3740 20567
rect 3790 20224 3846 20233
rect 3790 20159 3846 20168
rect 3804 19514 3832 20159
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3790 19408 3846 19417
rect 3700 19372 3752 19378
rect 3790 19343 3846 19352
rect 3700 19314 3752 19320
rect 3606 19272 3662 19281
rect 3606 19207 3662 19216
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3712 19122 3740 19314
rect 3804 19310 3832 19343
rect 3896 19310 3924 21519
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3988 19258 4016 22320
rect 4448 19700 4476 22320
rect 4448 19672 4752 19700
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4724 19378 4752 19672
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4528 19304 4580 19310
rect 3988 19230 4108 19258
rect 4804 19304 4856 19310
rect 4580 19252 4804 19258
rect 4528 19246 4856 19252
rect 4540 19230 4844 19246
rect 3620 18884 3648 19110
rect 3712 19094 4016 19122
rect 3700 18896 3752 18902
rect 3620 18856 3700 18884
rect 3700 18838 3752 18844
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3514 16008 3570 16017
rect 3514 15943 3570 15952
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3528 15434 3556 15943
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3436 13954 3464 14418
rect 3344 13938 3464 13954
rect 3332 13932 3464 13938
rect 3384 13926 3464 13932
rect 3332 13874 3384 13880
rect 3436 13530 3464 13926
rect 3620 13802 3648 18702
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 3606 13696 3662 13705
rect 3606 13631 3662 13640
rect 3620 13530 3648 13631
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3238 13288 3294 13297
rect 3238 13223 3294 13232
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3252 11830 3280 12786
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3252 10674 3280 11766
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3344 10130 3372 12650
rect 3528 12374 3556 13330
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3620 12753 3648 13126
rect 3606 12744 3662 12753
rect 3712 12714 3740 14758
rect 3804 13258 3832 18090
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 3896 16250 3924 16594
rect 3988 16561 4016 19094
rect 3974 16552 4030 16561
rect 3974 16487 4030 16496
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 4080 16182 4108 19230
rect 4908 18630 4936 22320
rect 5262 19408 5318 19417
rect 5262 19343 5318 19352
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5000 18902 5028 19110
rect 4988 18896 5040 18902
rect 4988 18838 5040 18844
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4160 18352 4212 18358
rect 4212 18300 4292 18306
rect 4160 18294 4292 18300
rect 4172 18278 4292 18294
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4172 17542 4200 18158
rect 4264 17882 4292 18278
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16250 4200 16934
rect 4264 16794 4292 17682
rect 4620 17672 4672 17678
rect 4618 17640 4620 17649
rect 4672 17640 4674 17649
rect 4618 17575 4674 17584
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4724 16794 4752 18566
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4816 17338 4844 17614
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 5000 17202 5028 18090
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4896 17128 4948 17134
rect 4894 17096 4896 17105
rect 4948 17096 4950 17105
rect 4894 17031 4950 17040
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 4080 15638 4108 15914
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 15706 4200 15846
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 4080 15026 4108 15574
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3976 14408 4028 14414
rect 4080 14396 4108 14962
rect 4028 14368 4108 14396
rect 3976 14350 4028 14356
rect 4264 14278 4292 15438
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13530 4108 13670
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3896 12986 3924 13330
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3606 12679 3662 12688
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 3516 11076 3568 11082
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3068 8634 3096 8978
rect 3252 8974 3280 9318
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3068 8378 3096 8570
rect 3068 8350 3188 8378
rect 3160 7886 3188 8350
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3148 5840 3200 5846
rect 2962 5808 3018 5817
rect 3148 5782 3200 5788
rect 2962 5743 3018 5752
rect 3160 4865 3188 5782
rect 3146 4856 3202 4865
rect 3146 4791 3202 4800
rect 3344 3913 3372 10066
rect 3436 7290 3464 11047
rect 3516 11018 3568 11024
rect 3528 10198 3556 11018
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3528 9178 3556 9522
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3620 7410 3648 11562
rect 3712 11150 3740 12174
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11762 3832 12038
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3712 10538 3740 11086
rect 3804 11082 3832 11494
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3896 10810 3924 12718
rect 3988 11626 4016 12718
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 4080 10962 4108 13194
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3988 10934 4108 10962
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3988 10690 4016 10934
rect 4066 10840 4122 10849
rect 4066 10775 4068 10784
rect 4120 10775 4122 10784
rect 4068 10746 4120 10752
rect 3804 10662 4016 10690
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 3712 10062 3740 10474
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3712 9586 3740 9998
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3712 9178 3740 9318
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3804 7585 3832 10662
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3896 9042 3924 10066
rect 3974 10024 4030 10033
rect 3974 9959 4030 9968
rect 3988 9926 4016 9959
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 4080 9722 4108 10367
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4172 9518 4200 12922
rect 4264 12782 4292 13398
rect 4724 13326 4752 13874
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4816 12986 4844 16934
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4356 12442 4384 12854
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4264 11354 4292 12242
rect 4448 12238 4476 12786
rect 4816 12714 4844 12922
rect 4908 12714 4936 16730
rect 5000 16590 5028 17138
rect 5092 17134 5120 17818
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 16046 5028 16390
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5000 12986 5028 13670
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 5092 12306 5120 16594
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5184 15638 5212 16458
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5184 15178 5212 15574
rect 5276 15314 5304 19343
rect 5368 18290 5396 22320
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5828 18816 5856 19382
rect 5736 18788 5856 18816
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5460 18222 5488 18566
rect 5632 18352 5684 18358
rect 5632 18294 5684 18300
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5368 17678 5396 18090
rect 5538 17776 5594 17785
rect 5644 17746 5672 18294
rect 5538 17711 5594 17720
rect 5632 17740 5684 17746
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5368 17066 5396 17614
rect 5552 17338 5580 17711
rect 5632 17682 5684 17688
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5368 15434 5396 16186
rect 5460 15978 5488 17206
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5630 16416 5686 16425
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5552 15314 5580 16390
rect 5736 16402 5764 18788
rect 5920 18714 5948 22320
rect 6380 18850 6408 22320
rect 6840 20074 6868 22320
rect 5828 18686 5948 18714
rect 6288 18822 6408 18850
rect 6564 20046 6868 20074
rect 5828 16674 5856 18686
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5920 17202 5948 18566
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6012 17134 6040 17478
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 5828 16658 5948 16674
rect 5828 16652 5960 16658
rect 5828 16646 5908 16652
rect 5908 16594 5960 16600
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5906 16552 5962 16561
rect 5686 16374 5764 16402
rect 5630 16351 5686 16360
rect 5736 16046 5764 16374
rect 5828 16114 5856 16526
rect 5906 16487 5962 16496
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5828 15706 5856 16050
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5276 15286 5580 15314
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5184 15150 5488 15178
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 5184 13512 5212 14486
rect 5276 13870 5304 14758
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5264 13524 5316 13530
rect 5184 13484 5264 13512
rect 5264 13466 5316 13472
rect 5276 12306 5304 13466
rect 5368 13258 5396 14962
rect 5460 14346 5488 15150
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5368 12850 5396 13194
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5368 12442 5396 12650
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4724 11354 4752 12174
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4264 10305 4292 11290
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4250 10296 4306 10305
rect 4250 10231 4306 10240
rect 4250 10160 4306 10169
rect 4632 10130 4660 10678
rect 4724 10198 4752 11290
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4816 10470 4844 10950
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4250 10095 4306 10104
rect 4620 10124 4672 10130
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4160 9376 4212 9382
rect 4264 9330 4292 10095
rect 4620 10066 4672 10072
rect 4632 10010 4660 10066
rect 4632 9982 4752 10010
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4724 9704 4752 9982
rect 4632 9676 4752 9704
rect 4632 9518 4660 9676
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4212 9324 4292 9330
rect 4160 9318 4292 9324
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4172 9302 4292 9318
rect 4250 9208 4306 9217
rect 4250 9143 4306 9152
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3896 8498 3924 8978
rect 4080 8537 4108 9046
rect 4066 8528 4122 8537
rect 3884 8492 3936 8498
rect 4066 8463 4122 8472
rect 3884 8434 3936 8440
rect 3790 7576 3846 7585
rect 3790 7511 3846 7520
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3436 7262 3832 7290
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 2778 2000 2834 2009
rect 2778 1935 2834 1944
rect 3344 1601 3372 2042
rect 3330 1592 3386 1601
rect 3330 1527 3386 1536
rect 938 1048 994 1057
rect 938 983 994 992
rect 3148 740 3200 746
rect 3148 682 3200 688
rect 3160 649 3188 682
rect 3146 640 3202 649
rect 3146 575 3202 584
rect 3804 480 3832 7262
rect 3896 3505 3924 8434
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4080 7750 4108 8055
rect 4172 7954 4200 8298
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 7177 4108 7210
rect 4264 7206 4292 9143
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 8022 4752 8774
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4816 7206 4844 8910
rect 4252 7200 4304 7206
rect 4066 7168 4122 7177
rect 4252 7142 4304 7148
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4066 7103 4122 7112
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3988 6225 4016 6802
rect 4066 6760 4122 6769
rect 4066 6695 4068 6704
rect 4120 6695 4122 6704
rect 4068 6666 4120 6672
rect 3974 6216 4030 6225
rect 3974 6151 4030 6160
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4066 5264 4122 5273
rect 4066 5199 4068 5208
rect 4120 5199 4122 5208
rect 4068 5170 4120 5176
rect 4066 4312 4122 4321
rect 4172 4298 4200 5714
rect 4122 4270 4200 4298
rect 4066 4247 4122 4256
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3882 3496 3938 3505
rect 3882 3431 3938 3440
rect 4080 2961 4108 4082
rect 4066 2952 4122 2961
rect 4066 2887 4122 2896
rect 4264 2553 4292 7142
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4250 2544 4306 2553
rect 4250 2479 4306 2488
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4816 2106 4844 7142
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 4908 746 4936 9318
rect 4988 8356 5040 8362
rect 4988 8298 5040 8304
rect 5000 7410 5028 8298
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5092 8090 5120 8230
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5184 7546 5212 8230
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4896 740 4948 746
rect 4896 682 4948 688
rect 3332 332 3384 338
rect 3332 274 3384 280
rect 3344 241 3372 274
rect 3330 232 3386 241
rect 3330 167 3386 176
rect 3790 0 3846 480
rect 5276 338 5304 12242
rect 5460 12186 5488 14010
rect 5552 13326 5580 15286
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5368 12158 5488 12186
rect 5368 10470 5396 12158
rect 5552 10996 5580 12378
rect 5460 10968 5580 10996
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 4146 5396 10406
rect 5460 6390 5488 10968
rect 5644 10826 5672 15302
rect 5920 12442 5948 16487
rect 6196 15094 6224 18362
rect 6288 15688 6316 18822
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6380 18426 6408 18702
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6472 18358 6500 18702
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6288 15660 6408 15688
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6288 15162 6316 15506
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 6288 14618 6316 15098
rect 6380 14958 6408 15660
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6380 14498 6408 14894
rect 6380 14482 6500 14498
rect 6380 14476 6512 14482
rect 6380 14470 6460 14476
rect 6460 14418 6512 14424
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5724 11824 5776 11830
rect 5722 11792 5724 11801
rect 5776 11792 5778 11801
rect 5722 11727 5778 11736
rect 5736 11286 5764 11727
rect 5920 11694 5948 12242
rect 6012 11762 6040 12582
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6104 11830 6132 12106
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5920 11150 5948 11630
rect 6564 11354 6592 20046
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6656 13326 6684 19926
rect 7102 19000 7158 19009
rect 7102 18935 7158 18944
rect 7116 18834 7144 18935
rect 7300 18850 7328 22320
rect 7378 19136 7434 19145
rect 7378 19071 7434 19080
rect 7392 18970 7420 19071
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7104 18828 7156 18834
rect 7300 18822 7696 18850
rect 7104 18770 7156 18776
rect 7024 17882 7052 18770
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7300 18290 7328 18702
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6748 17202 6776 17478
rect 6840 17270 6868 17478
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 7024 17105 7052 17682
rect 7010 17096 7066 17105
rect 7010 17031 7066 17040
rect 7024 16980 7052 17031
rect 6932 16952 7052 16980
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6748 16658 6776 16730
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6932 14906 6960 16952
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 7024 15026 7052 15846
rect 7116 15638 7144 18158
rect 7576 17678 7604 18226
rect 7564 17672 7616 17678
rect 7194 17640 7250 17649
rect 7564 17614 7616 17620
rect 7194 17575 7250 17584
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 7208 14958 7236 17575
rect 7576 17338 7604 17614
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7576 16658 7604 16730
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7392 16522 7420 16594
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7196 14952 7248 14958
rect 6932 14878 7052 14906
rect 7196 14894 7248 14900
rect 7024 14804 7052 14878
rect 7196 14816 7248 14822
rect 7024 14776 7144 14804
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6656 12986 6684 13262
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 5644 10798 6040 10826
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10532 5868 10538
rect 5816 10474 5868 10480
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 8634 5580 9386
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5552 7954 5580 8570
rect 5644 8362 5672 8842
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 8090 5672 8298
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5736 8022 5764 10406
rect 5828 8974 5856 10474
rect 5920 9926 5948 10610
rect 6012 10282 6040 10798
rect 6380 10606 6408 11018
rect 6368 10600 6420 10606
rect 6090 10568 6146 10577
rect 6368 10542 6420 10548
rect 6090 10503 6146 10512
rect 6104 10470 6132 10503
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6012 10254 6132 10282
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5920 9518 5948 9862
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5906 9072 5962 9081
rect 5906 9007 5962 9016
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5920 8838 5948 9007
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 6012 8090 6040 8910
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 6104 7954 6132 10254
rect 6380 10198 6408 10542
rect 6564 10470 6592 11290
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6748 10266 6776 13670
rect 6826 11928 6882 11937
rect 6826 11863 6882 11872
rect 6840 11558 6868 11863
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6932 11218 6960 14214
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7024 13326 7052 13942
rect 7116 13433 7144 14776
rect 7196 14758 7248 14764
rect 7208 14074 7236 14758
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 13530 7236 13670
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7102 13424 7158 13433
rect 7102 13359 7158 13368
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7208 12374 7236 12786
rect 7300 12782 7328 16118
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7392 15162 7420 15846
rect 7484 15706 7512 15846
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7576 15434 7604 16050
rect 7564 15428 7616 15434
rect 7564 15370 7616 15376
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7484 14804 7512 14962
rect 7392 14776 7512 14804
rect 7392 14278 7420 14776
rect 7576 14550 7604 15370
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7576 13938 7604 14486
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7668 12646 7696 18822
rect 7760 18086 7788 22320
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8220 18408 8248 22320
rect 8772 18970 8800 22320
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8312 18426 8340 18906
rect 8036 18380 8248 18408
rect 8300 18420 8352 18426
rect 7748 18080 7800 18086
rect 8036 18068 8064 18380
rect 8300 18362 8352 18368
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8404 18306 8432 18362
rect 8128 18278 8432 18306
rect 8128 18222 8156 18278
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8392 18080 8444 18086
rect 8036 18040 8248 18068
rect 7748 18022 7800 18028
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17354 8248 18040
rect 8392 18022 8444 18028
rect 8220 17326 8340 17354
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 15570 7788 16934
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8220 16726 8248 17206
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8312 16572 8340 17326
rect 8220 16544 8340 16572
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15706 8248 16544
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7760 15026 7788 15506
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7760 14006 7788 14962
rect 8220 14958 8248 15642
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14278 8248 14758
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12850 8064 13126
rect 8024 12844 8076 12850
rect 8076 12804 8248 12832
rect 8024 12786 8076 12792
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7300 11880 7328 12582
rect 7668 12442 7696 12582
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7760 12374 7788 12718
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7116 11852 7328 11880
rect 7116 11558 7144 11852
rect 7576 11762 7604 12038
rect 8220 11762 8248 12804
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8206 11656 8262 11665
rect 8206 11591 8262 11600
rect 8220 11558 8248 11591
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8312 11286 8340 12038
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7208 10266 7236 10406
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7024 9042 7052 9386
rect 7300 9178 7328 10406
rect 7576 10062 7604 10610
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8312 10266 8340 10950
rect 8404 10606 8432 18022
rect 8850 17640 8906 17649
rect 8850 17575 8906 17584
rect 8864 17542 8892 17575
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8758 16688 8814 16697
rect 8588 16522 8616 16662
rect 8758 16623 8814 16632
rect 8576 16516 8628 16522
rect 8576 16458 8628 16464
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8680 16250 8708 16458
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8680 16046 8708 16186
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8772 15638 8800 16623
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8864 15706 8892 15914
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8496 14890 8524 15506
rect 8588 15026 8616 15574
rect 8772 15178 8800 15574
rect 8680 15150 8800 15178
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8496 14074 8524 14826
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 12102 8524 13806
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12986 8616 13262
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8680 12832 8708 15150
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8864 14074 8892 14282
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8680 12804 8892 12832
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8668 12368 8720 12374
rect 8666 12336 8668 12345
rect 8720 12336 8722 12345
rect 8666 12271 8722 12280
rect 8772 12238 8800 12650
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8484 12096 8536 12102
rect 8864 12084 8892 12804
rect 8484 12038 8536 12044
rect 8680 12056 8892 12084
rect 8680 11354 8708 12056
rect 8850 11656 8906 11665
rect 8850 11591 8906 11600
rect 8864 11354 8892 11591
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7576 9110 7604 9998
rect 8220 9722 8248 9998
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8496 9450 8524 11018
rect 8956 10674 8984 19314
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 17678 9076 18566
rect 9140 18154 9168 18702
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9140 17542 9168 18090
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9232 16726 9260 22320
rect 9692 18850 9720 22320
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9508 18822 9720 18850
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9324 17338 9352 17682
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9416 17066 9444 17682
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9508 16538 9536 18822
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 17610 9720 18702
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9784 17678 9812 18090
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9324 16510 9536 16538
rect 9220 15088 9272 15094
rect 9324 15076 9352 16510
rect 9588 16448 9640 16454
rect 9586 16416 9588 16425
rect 9640 16416 9642 16425
rect 9586 16351 9642 16360
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9272 15048 9352 15076
rect 9220 15030 9272 15036
rect 9324 14618 9352 15048
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9140 13870 9168 14350
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9508 13274 9536 15846
rect 9876 14618 9904 19246
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9968 18329 9996 18634
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9954 18320 10010 18329
rect 9954 18255 10010 18264
rect 9956 17808 10008 17814
rect 9954 17776 9956 17785
rect 10008 17776 10010 17785
rect 10060 17746 10088 18362
rect 9954 17711 10010 17720
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9968 17202 9996 17478
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10060 16114 10088 17682
rect 10152 16590 10180 22320
rect 10508 19168 10560 19174
rect 10414 19136 10470 19145
rect 10508 19110 10560 19116
rect 10414 19071 10470 19080
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10230 18728 10286 18737
rect 10230 18663 10286 18672
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9956 15632 10008 15638
rect 9954 15600 9956 15609
rect 10008 15600 10010 15609
rect 10060 15570 10088 16050
rect 10244 15570 10272 18663
rect 10336 17338 10364 18770
rect 10428 17882 10456 19071
rect 10520 18737 10548 19110
rect 10612 18850 10640 22320
rect 11072 19394 11100 22320
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11624 19530 11652 22320
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11624 19502 11928 19530
rect 11072 19366 11836 19394
rect 11428 19304 11480 19310
rect 11164 19264 11428 19292
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10612 18822 10824 18850
rect 10600 18760 10652 18766
rect 10506 18728 10562 18737
rect 10600 18702 10652 18708
rect 10506 18663 10562 18672
rect 10612 18426 10640 18702
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10428 17626 10456 17818
rect 10508 17808 10560 17814
rect 10612 17796 10640 18362
rect 10560 17768 10640 17796
rect 10508 17750 10560 17756
rect 10428 17598 10640 17626
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10414 17232 10470 17241
rect 10414 17167 10470 17176
rect 10428 16454 10456 17167
rect 10520 16794 10548 17274
rect 10612 17134 10640 17598
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 9954 15535 10010 15544
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14618 9996 14758
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 13394 9628 14350
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 13938 9904 14010
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9508 13246 9628 13274
rect 9494 12064 9550 12073
rect 9494 11999 9550 12008
rect 9310 11928 9366 11937
rect 9310 11863 9366 11872
rect 9324 11626 9352 11863
rect 9402 11792 9458 11801
rect 9402 11727 9404 11736
rect 9456 11727 9458 11736
rect 9404 11698 9456 11704
rect 9508 11626 9536 11999
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9036 11552 9088 11558
rect 9404 11552 9456 11558
rect 9088 11500 9404 11506
rect 9036 11494 9456 11500
rect 9048 11478 9444 11494
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9140 11121 9168 11154
rect 9600 11150 9628 13246
rect 9692 12986 9720 13738
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9588 11144 9640 11150
rect 9126 11112 9182 11121
rect 9588 11086 9640 11092
rect 9126 11047 9182 11056
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10674 9444 11018
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 8574 10568 8630 10577
rect 8864 10554 8892 10610
rect 8864 10526 8984 10554
rect 8574 10503 8630 10512
rect 8588 10062 8616 10503
rect 8956 10470 8984 10526
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8864 10130 8892 10406
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 8680 8838 8708 9862
rect 8956 9450 8984 10406
rect 9600 9450 9628 10678
rect 9692 10674 9720 11698
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9692 10266 9720 10610
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9692 10130 9720 10202
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9692 9602 9720 10066
rect 9692 9574 9812 9602
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9692 9042 9720 9574
rect 9784 9518 9812 9574
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 5552 7478 5580 7890
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8680 3534 8708 8774
rect 9692 7410 9720 8978
rect 9876 8022 9904 13874
rect 10060 13802 10088 15506
rect 10244 14600 10272 15506
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10244 14572 10364 14600
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10244 13530 10272 14418
rect 10336 14396 10364 14572
rect 10428 14550 10456 14758
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10336 14368 10456 14396
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10336 13977 10364 14214
rect 10322 13968 10378 13977
rect 10322 13903 10378 13912
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9968 11762 9996 13398
rect 10230 13288 10286 13297
rect 10230 13223 10286 13232
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9968 8838 9996 10066
rect 10244 9636 10272 13223
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 12442 10364 12582
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10244 9608 10364 9636
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10046 9208 10102 9217
rect 10046 9143 10102 9152
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8498 9996 8774
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9876 7206 9904 7958
rect 10060 7818 10088 9143
rect 10152 9110 10180 9318
rect 10336 9217 10364 9608
rect 10322 9208 10378 9217
rect 10322 9143 10378 9152
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10336 8634 10364 9046
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10428 8090 10456 14368
rect 10520 13802 10548 14962
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10612 14074 10640 14350
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10520 13326 10548 13738
rect 10612 13530 10640 13738
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10704 12646 10732 16934
rect 10796 12850 10824 18822
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10888 17202 10916 18090
rect 10980 17921 11008 18906
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10966 17912 11022 17921
rect 10966 17847 11022 17856
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 11072 17134 11100 18022
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10980 16794 11008 16934
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 11164 16674 11192 19264
rect 11428 19246 11480 19252
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11624 18358 11652 18702
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11716 18465 11744 18634
rect 11702 18456 11758 18465
rect 11702 18391 11758 18400
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11624 17762 11652 18090
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 17882 11744 18022
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11624 17734 11744 17762
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11072 16646 11192 16674
rect 11440 16658 11468 16934
rect 11428 16652 11480 16658
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10874 13560 10930 13569
rect 10874 13495 10930 13504
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11694 10548 12174
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10428 7528 10456 8026
rect 10508 7540 10560 7546
rect 10428 7500 10508 7528
rect 10508 7482 10560 7488
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 10612 6186 10640 11290
rect 10704 10198 10732 12378
rect 10796 11558 10824 12786
rect 10888 12782 10916 13495
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 8498 10824 9318
rect 10888 8974 10916 12582
rect 10980 12442 11008 16526
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10980 11694 11008 12242
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11354 11008 11630
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10980 10713 11008 10746
rect 10966 10704 11022 10713
rect 10966 10639 11022 10648
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10980 10266 11008 10474
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 8566 11008 8774
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 11072 7970 11100 16646
rect 11428 16594 11480 16600
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11164 15910 11192 16526
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11624 16250 11652 17478
rect 11716 16794 11744 17734
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11716 16250 11744 16594
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11520 16176 11572 16182
rect 11624 16153 11652 16186
rect 11520 16118 11572 16124
rect 11610 16144 11666 16153
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 15638 11468 15846
rect 11532 15706 11560 16118
rect 11610 16079 11666 16088
rect 11704 16108 11756 16114
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11624 15502 11652 16079
rect 11704 16050 11756 16056
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11716 15162 11744 16050
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11164 14482 11192 15030
rect 11716 14822 11744 15098
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 12306 11192 14214
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11532 13462 11560 13942
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11348 12306 11376 12718
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10606 11192 10950
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 10742 11652 14418
rect 11808 13818 11836 19366
rect 11900 16114 11928 19502
rect 11992 19378 12020 19858
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12084 19145 12112 22320
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12176 19378 12204 19790
rect 12544 19394 12572 22320
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12164 19372 12216 19378
rect 12544 19366 12664 19394
rect 12164 19314 12216 19320
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12070 19136 12126 19145
rect 12070 19071 12126 19080
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11992 16590 12020 17138
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11992 16046 12020 16526
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 12084 15586 12112 18634
rect 12452 18306 12480 18838
rect 12544 18426 12572 19246
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12452 18278 12572 18306
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17610 12204 18022
rect 12544 17746 12572 18278
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12360 17105 12388 17206
rect 12440 17128 12492 17134
rect 12346 17096 12402 17105
rect 12440 17070 12492 17076
rect 12346 17031 12402 17040
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15706 12204 15846
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 11888 15564 11940 15570
rect 12084 15558 12204 15586
rect 11888 15506 11940 15512
rect 11900 14006 11928 15506
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11992 14550 12020 15302
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11992 13938 12020 14486
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11716 13790 11836 13818
rect 11886 13832 11942 13841
rect 11716 11286 11744 13790
rect 11886 13767 11942 13776
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 12850 11836 13670
rect 11900 13530 11928 13767
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11808 11830 11836 12242
rect 11900 12220 11928 13466
rect 11992 13326 12020 13874
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12084 12374 12112 15302
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 11900 12192 12112 12220
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11152 10600 11204 10606
rect 11520 10600 11572 10606
rect 11152 10542 11204 10548
rect 11518 10568 11520 10577
rect 11572 10568 11574 10577
rect 11716 10538 11744 11222
rect 11518 10503 11574 10512
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 9518 11192 10406
rect 11794 10024 11850 10033
rect 11794 9959 11850 9968
rect 11808 9926 11836 9959
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11256 9110 11284 9454
rect 11348 9178 11376 9590
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8362 11652 9318
rect 11992 8634 12020 9862
rect 12084 9042 12112 12192
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12084 8480 12112 8774
rect 12176 8673 12204 15558
rect 12268 15366 12296 16730
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12268 14618 12296 14962
rect 12360 14929 12388 16934
rect 12452 15910 12480 17070
rect 12544 16590 12572 17682
rect 12636 17105 12664 19366
rect 12728 18290 12756 19654
rect 12912 19378 12940 19858
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12912 18057 12940 19314
rect 12898 18048 12954 18057
rect 12898 17983 12954 17992
rect 12622 17096 12678 17105
rect 13004 17082 13032 22320
rect 13464 20058 13492 22320
rect 13924 20058 13952 22320
rect 14476 20058 14504 22320
rect 14936 20346 14964 22320
rect 14936 20318 15056 20346
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13188 18902 13216 19246
rect 13268 19236 13320 19242
rect 13268 19178 13320 19184
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 13188 18426 13216 18838
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13096 17202 13124 18022
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12622 17031 12678 17040
rect 12820 17054 13032 17082
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12440 15632 12492 15638
rect 12438 15600 12440 15609
rect 12492 15600 12494 15609
rect 12438 15535 12494 15544
rect 12544 15434 12572 16118
rect 12636 16046 12664 17031
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12728 16250 12756 16662
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12636 15473 12664 15506
rect 12622 15464 12678 15473
rect 12532 15428 12584 15434
rect 12622 15399 12678 15408
rect 12532 15370 12584 15376
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12440 14952 12492 14958
rect 12346 14920 12402 14929
rect 12440 14894 12492 14900
rect 12636 14940 12664 15302
rect 12716 14952 12768 14958
rect 12636 14912 12716 14940
rect 12346 14855 12402 14864
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12268 14482 12296 14554
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12268 13870 12296 13942
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12256 13320 12308 13326
rect 12360 13297 12388 14855
rect 12452 14074 12480 14894
rect 12636 14414 12664 14912
rect 12716 14894 12768 14900
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12820 13870 12848 17054
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13569 12848 13806
rect 12806 13560 12862 13569
rect 12440 13524 12492 13530
rect 12806 13495 12862 13504
rect 12440 13466 12492 13472
rect 12452 13394 12480 13466
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12728 13297 12756 13330
rect 12256 13262 12308 13268
rect 12346 13288 12402 13297
rect 12268 12850 12296 13262
rect 12714 13288 12770 13297
rect 12346 13223 12402 13232
rect 12532 13252 12584 13258
rect 12912 13274 12940 16934
rect 12990 16144 13046 16153
rect 12990 16079 12992 16088
rect 13044 16079 13046 16088
rect 12992 16050 13044 16056
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 12820 13258 12940 13274
rect 12714 13223 12770 13232
rect 12808 13252 12940 13258
rect 12532 13194 12584 13200
rect 12860 13246 12940 13252
rect 12808 13194 12860 13200
rect 12544 13138 12572 13194
rect 12452 13110 12572 13138
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12452 12730 12480 13110
rect 12912 12918 12940 13246
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12360 12714 12480 12730
rect 12348 12708 12480 12714
rect 12400 12702 12480 12708
rect 12348 12650 12400 12656
rect 12636 12442 12664 12786
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12254 11248 12310 11257
rect 12254 11183 12310 11192
rect 12440 11212 12492 11218
rect 12268 11150 12296 11183
rect 12440 11154 12492 11160
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12360 9586 12388 9998
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12254 9208 12310 9217
rect 12254 9143 12310 9152
rect 12268 9042 12296 9143
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12162 8664 12218 8673
rect 12162 8599 12218 8608
rect 12164 8492 12216 8498
rect 12084 8452 12164 8480
rect 12164 8434 12216 8440
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11164 8090 11192 8298
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11796 8016 11848 8022
rect 10968 7948 11020 7954
rect 11072 7942 11192 7970
rect 11796 7958 11848 7964
rect 10968 7890 11020 7896
rect 10874 7848 10930 7857
rect 10980 7834 11008 7890
rect 10980 7806 11100 7834
rect 10874 7783 10876 7792
rect 10928 7783 10930 7792
rect 10876 7754 10928 7760
rect 11072 7274 11100 7806
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10612 5710 10640 6122
rect 10888 6066 10916 7210
rect 11072 7018 11100 7210
rect 10980 6990 11100 7018
rect 10980 6338 11008 6990
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11072 6458 11100 6802
rect 11164 6662 11192 7942
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11624 7041 11652 7686
rect 11716 7546 11744 7890
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11610 7032 11666 7041
rect 11610 6967 11666 6976
rect 11716 6730 11744 7482
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10980 6310 11100 6338
rect 11716 6322 11744 6666
rect 10888 6038 11008 6066
rect 10980 5710 11008 6038
rect 11072 5710 11100 6310
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 3738 11100 5646
rect 11164 5370 11192 6190
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5914 11468 6054
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11808 5846 11836 7958
rect 11900 7342 11928 8230
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11992 7206 12020 7890
rect 12070 7848 12126 7857
rect 12070 7783 12072 7792
rect 12124 7783 12126 7792
rect 12072 7754 12124 7760
rect 12176 7342 12204 8434
rect 12360 7886 12388 9522
rect 12452 8922 12480 11154
rect 12544 9722 12572 12106
rect 12636 11286 12664 12378
rect 12728 11694 12756 12854
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12820 12442 12848 12718
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12912 12186 12940 12718
rect 12820 12158 12940 12186
rect 12820 11898 12848 12158
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12912 11762 12940 12038
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12806 10704 12862 10713
rect 12806 10639 12862 10648
rect 12820 10606 12848 10639
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12530 9072 12586 9081
rect 12530 9007 12532 9016
rect 12584 9007 12586 9016
rect 12532 8978 12584 8984
rect 12452 8894 12572 8922
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8673 12480 8774
rect 12438 8664 12494 8673
rect 12438 8599 12494 8608
rect 12544 8498 12572 8894
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12636 8022 12664 10134
rect 12728 8090 12756 10406
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12268 7274 12296 7686
rect 12360 7478 12388 7686
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 12268 6798 12296 7210
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12452 6662 12480 7482
rect 12544 7206 12572 7754
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12544 6458 12572 6802
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11808 3738 11836 5782
rect 11900 5778 11928 6258
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11992 5846 12020 6122
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11900 5522 11928 5714
rect 11980 5568 12032 5574
rect 11900 5516 11980 5522
rect 11900 5510 12032 5516
rect 11900 5494 12020 5510
rect 11900 5234 11928 5494
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 12820 4146 12848 9998
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9178 12940 9318
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13004 9081 13032 15914
rect 13096 15366 13124 17138
rect 13280 17134 13308 19178
rect 13372 18834 13400 19790
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18970 13492 19178
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13360 18284 13412 18290
rect 13464 18272 13492 18906
rect 13412 18244 13492 18272
rect 13360 18226 13412 18232
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13096 13462 13124 15030
rect 13188 14006 13216 15506
rect 13280 15502 13308 16526
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 15065 13308 15438
rect 13266 15056 13322 15065
rect 13266 14991 13322 15000
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 12990 9072 13046 9081
rect 12990 9007 13046 9016
rect 13096 8945 13124 12854
rect 13188 11558 13216 13806
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13082 8936 13138 8945
rect 13082 8871 13138 8880
rect 13188 7546 13216 10406
rect 13280 10266 13308 13330
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12442 13400 13126
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13372 11762 13400 12174
rect 13464 12102 13492 13262
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13556 11234 13584 19858
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 14016 18290 14044 18702
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13818 17912 13874 17921
rect 13728 17876 13780 17882
rect 14016 17882 14044 18226
rect 13818 17847 13874 17856
rect 14004 17876 14056 17882
rect 13728 17818 13780 17824
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13648 17270 13676 17546
rect 13740 17542 13768 17818
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13740 13954 13768 14486
rect 13648 13926 13768 13954
rect 13648 13326 13676 13926
rect 13832 13818 13860 17847
rect 14004 17818 14056 17824
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13740 13790 13860 13818
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12646 13676 13126
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13740 11642 13768 13790
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13648 11614 13768 11642
rect 13648 11354 13676 11614
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13372 11206 13584 11234
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9178 13308 10066
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13188 7274 13216 7482
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 11164 898 11192 3606
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11164 870 11376 898
rect 11348 480 11376 870
rect 13280 649 13308 8978
rect 13372 6934 13400 11206
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10674 13584 10950
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10062 13584 10610
rect 13740 10606 13768 11494
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9586 13584 9998
rect 13648 9654 13676 10066
rect 13740 9654 13768 10406
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13544 9580 13596 9586
rect 13464 9540 13544 9568
rect 13464 9058 13492 9540
rect 13544 9522 13596 9528
rect 13740 9217 13768 9590
rect 13832 9466 13860 13670
rect 13924 12832 13952 16118
rect 14004 14884 14056 14890
rect 14004 14826 14056 14832
rect 14016 14346 14044 14826
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 13938 14044 14282
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14016 13326 14044 13874
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14108 12866 14136 19858
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14832 19304 14884 19310
rect 14924 19304 14976 19310
rect 14884 19264 14924 19292
rect 14832 19246 14884 19252
rect 15028 19292 15056 20318
rect 15396 20058 15424 22320
rect 15856 20074 15884 22320
rect 15856 20058 15976 20074
rect 15384 20052 15436 20058
rect 15856 20052 15988 20058
rect 15856 20046 15936 20052
rect 15384 19994 15436 20000
rect 15936 19994 15988 20000
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15028 19264 15128 19292
rect 14924 19246 14976 19252
rect 14200 18086 14228 19246
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 15016 19168 15068 19174
rect 15100 19156 15128 19264
rect 15200 19168 15252 19174
rect 15100 19128 15148 19156
rect 15016 19110 15068 19116
rect 14568 18952 14596 19110
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14568 18924 14872 18952
rect 14844 18766 14872 18924
rect 15028 18850 15056 19110
rect 15120 18970 15148 19128
rect 15200 19110 15252 19116
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15212 18850 15240 19110
rect 15396 18952 15424 19110
rect 15028 18822 15240 18850
rect 15304 18924 15424 18952
rect 14648 18760 14700 18766
rect 14646 18728 14648 18737
rect 14832 18760 14884 18766
rect 14700 18728 14702 18737
rect 14832 18702 14884 18708
rect 14646 18663 14702 18672
rect 14844 18154 14872 18702
rect 15304 18698 15332 18924
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 14200 16130 14228 18022
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14462 17912 14518 17921
rect 14280 17876 14332 17882
rect 14684 17904 14980 17924
rect 14462 17847 14464 17856
rect 14280 17818 14332 17824
rect 14516 17847 14518 17856
rect 14464 17818 14516 17824
rect 14292 17202 14320 17818
rect 15108 17808 15160 17814
rect 15106 17776 15108 17785
rect 15160 17776 15162 17785
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14556 17740 14608 17746
rect 15106 17711 15162 17720
rect 14556 17682 14608 17688
rect 14384 17270 14412 17682
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14384 17082 14412 17206
rect 14568 17105 14596 17682
rect 15016 17672 15068 17678
rect 15212 17660 15240 18022
rect 15304 17882 15332 18362
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15212 17632 15332 17660
rect 15016 17614 15068 17620
rect 14554 17096 14610 17105
rect 14280 17060 14332 17066
rect 14384 17054 14504 17082
rect 14280 17002 14332 17008
rect 14292 16794 14320 17002
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14384 16250 14412 16934
rect 14476 16794 14504 17054
rect 14554 17031 14610 17040
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14568 16561 14596 17031
rect 15028 16998 15056 17614
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14554 16552 14610 16561
rect 14554 16487 14610 16496
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14200 16102 14412 16130
rect 14278 15464 14334 15473
rect 14278 15399 14280 15408
rect 14332 15399 14334 15408
rect 14280 15370 14332 15376
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14200 12986 14228 13670
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14292 12986 14320 13330
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14108 12838 14228 12866
rect 13924 12804 14044 12832
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13924 10266 13952 12650
rect 14016 12322 14044 12804
rect 14016 12294 14136 12322
rect 14108 11286 14136 12294
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14108 10674 14136 11222
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9722 13952 9862
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13832 9438 13952 9466
rect 13924 9382 13952 9438
rect 13912 9376 13964 9382
rect 13818 9344 13874 9353
rect 13912 9318 13964 9324
rect 13818 9279 13874 9288
rect 13726 9208 13782 9217
rect 13832 9178 13860 9279
rect 13726 9143 13782 9152
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13464 9030 13768 9058
rect 13464 8974 13492 9030
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13740 8922 13768 9030
rect 13820 8968 13872 8974
rect 13740 8916 13820 8922
rect 13740 8910 13872 8916
rect 13740 8894 13860 8910
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13924 7478 13952 8842
rect 14016 8362 14044 9998
rect 14108 9586 14136 10406
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13634 7032 13690 7041
rect 13634 6967 13636 6976
rect 13688 6967 13690 6976
rect 13636 6938 13688 6944
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6322 13768 6734
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13832 5370 13860 6122
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 14108 2106 14136 9318
rect 14200 9110 14228 12838
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 11762 14320 12242
rect 14384 12238 14412 16102
rect 14844 16046 14872 16662
rect 15028 16658 15056 16934
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15028 16114 15056 16594
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14384 10538 14412 11290
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14278 10432 14334 10441
rect 14278 10367 14334 10376
rect 14292 9178 14320 10367
rect 14476 10198 14504 15846
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15028 15609 15056 15914
rect 15014 15600 15070 15609
rect 14556 15564 14608 15570
rect 15014 15535 15070 15544
rect 14556 15506 14608 15512
rect 14568 15162 14596 15506
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14568 15026 14596 15098
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 14385 14688 14418
rect 15016 14408 15068 14414
rect 14646 14376 14702 14385
rect 15016 14350 15068 14356
rect 14646 14311 14702 14320
rect 15028 13938 15056 14350
rect 15212 14074 15240 14758
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15028 12850 15056 13874
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15200 13728 15252 13734
rect 15304 13716 15332 17632
rect 15252 13688 15332 13716
rect 15200 13670 15252 13676
rect 15120 12986 15148 13670
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15212 12866 15240 13670
rect 15396 13462 15424 18770
rect 15488 17184 15516 19858
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18426 15608 19110
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15672 18465 15700 18906
rect 15764 18902 15792 19314
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15658 18456 15714 18465
rect 15568 18420 15620 18426
rect 15764 18426 15792 18838
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15948 18630 15976 18702
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15936 18624 15988 18630
rect 16132 18601 16160 19110
rect 15936 18566 15988 18572
rect 16118 18592 16174 18601
rect 15658 18391 15714 18400
rect 15752 18420 15804 18426
rect 15568 18362 15620 18368
rect 15752 18362 15804 18368
rect 15856 18358 15884 18566
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15660 17740 15712 17746
rect 15712 17700 15792 17728
rect 15660 17682 15712 17688
rect 15488 17156 15608 17184
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16658 15516 17002
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14550 15516 14758
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15120 12838 15240 12866
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14568 10826 14596 11630
rect 15120 11626 15148 12838
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15212 11218 15240 12718
rect 15304 11778 15332 13330
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15396 12782 15424 12854
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15396 11914 15424 12582
rect 15396 11886 15516 11914
rect 15304 11750 15424 11778
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15304 11354 15332 11562
rect 15396 11558 15424 11750
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14568 10798 14688 10826
rect 14660 10674 14688 10798
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14568 10044 14596 10610
rect 14936 10606 14964 11086
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 14648 10056 14700 10062
rect 14568 10016 14648 10044
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14188 8968 14240 8974
rect 14186 8936 14188 8945
rect 14240 8936 14242 8945
rect 14186 8871 14242 8880
rect 14200 2553 14228 8871
rect 14292 8090 14320 8978
rect 14476 8090 14504 9318
rect 14568 8906 14596 10016
rect 14648 9998 14700 10004
rect 14738 9616 14794 9625
rect 14738 9551 14794 9560
rect 14752 9518 14780 9551
rect 14740 9512 14792 9518
rect 14936 9489 14964 10134
rect 14740 9454 14792 9460
rect 14922 9480 14978 9489
rect 14922 9415 14978 9424
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 15028 8634 15056 10202
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15120 8362 15148 9522
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14476 7002 14504 7890
rect 14568 7886 14596 8298
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 15120 7546 15148 8298
rect 15212 8294 15240 11154
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15304 9518 15332 9862
rect 15488 9625 15516 11886
rect 15474 9616 15530 9625
rect 15580 9586 15608 17156
rect 15764 16454 15792 17700
rect 15856 17678 15884 18090
rect 15948 17678 15976 18566
rect 16118 18527 16174 18536
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15844 17128 15896 17134
rect 15948 17116 15976 17614
rect 15896 17088 15976 17116
rect 15844 17070 15896 17076
rect 15856 16590 15884 17070
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15672 12918 15700 15982
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15672 11082 15700 11630
rect 15764 11121 15792 16390
rect 15948 15502 15976 16594
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15842 15056 15898 15065
rect 15842 14991 15844 15000
rect 15896 14991 15898 15000
rect 15844 14962 15896 14968
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15948 14074 15976 14418
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 12306 15884 12786
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15750 11112 15806 11121
rect 15660 11076 15712 11082
rect 15750 11047 15806 11056
rect 15660 11018 15712 11024
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15764 10130 15792 10746
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15474 9551 15530 9560
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15948 9450 15976 13330
rect 16040 12424 16068 17682
rect 16132 17524 16160 18527
rect 16316 18426 16344 22320
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16592 19310 16620 19858
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16592 18630 16620 18770
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16684 18358 16712 18566
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16224 17649 16252 17818
rect 16592 17814 16620 18158
rect 16580 17808 16632 17814
rect 16580 17750 16632 17756
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16210 17640 16266 17649
rect 16210 17575 16266 17584
rect 16132 17496 16252 17524
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16132 13394 16160 15846
rect 16224 14498 16252 17496
rect 16316 16250 16344 17682
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16302 16008 16358 16017
rect 16302 15943 16358 15952
rect 16316 14618 16344 15943
rect 16408 15910 16436 16390
rect 16592 15994 16620 17478
rect 16776 17184 16804 22320
rect 17328 19938 17356 22320
rect 17498 22128 17554 22137
rect 17498 22063 17554 22072
rect 17236 19910 17356 19938
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16684 17156 16804 17184
rect 16684 16794 16712 17156
rect 16868 17134 16896 18158
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 16250 16712 16594
rect 16776 16250 16804 17002
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16592 15966 16804 15994
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16500 15706 16528 15846
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16684 15434 16712 15846
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16488 14544 16540 14550
rect 16224 14470 16436 14498
rect 16488 14486 16540 14492
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16224 13326 16252 13738
rect 16316 13530 16344 13806
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16304 12708 16356 12714
rect 16304 12650 16356 12656
rect 16040 12396 16160 12424
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 16040 11898 16068 12242
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16132 11286 16160 12396
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16132 10266 16160 11222
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16224 10810 16252 11018
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16316 10577 16344 12650
rect 16302 10568 16358 10577
rect 16302 10503 16358 10512
rect 16316 10470 16344 10503
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 16224 9382 16252 10066
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 15120 6798 15148 7482
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14660 6458 14688 6734
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15212 6322 15240 6394
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15304 6202 15332 7142
rect 15488 7002 15516 9114
rect 16224 9042 16252 9318
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 15948 7886 15976 8978
rect 16316 8634 16344 9454
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 8022 16068 8230
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15488 6866 15516 6938
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 6458 15700 6802
rect 15948 6798 15976 7278
rect 16040 6798 16068 7958
rect 16408 6866 16436 14470
rect 16500 13394 16528 14486
rect 16592 13938 16620 15302
rect 16776 15008 16804 15966
rect 16856 15496 16908 15502
rect 16960 15484 16988 18158
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16908 15456 16988 15484
rect 16856 15438 16908 15444
rect 16684 14980 16804 15008
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16684 13512 16712 14980
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16776 14618 16804 14826
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16776 13938 16804 14554
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16868 13841 16896 15438
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16960 14074 16988 14418
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16854 13832 16910 13841
rect 16854 13767 16910 13776
rect 16684 13484 16988 13512
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16592 10198 16620 11290
rect 16684 10810 16712 11494
rect 16960 11354 16988 13484
rect 17052 13258 17080 15846
rect 17144 13938 17172 19722
rect 17236 17610 17264 19910
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 15978 17264 16390
rect 17224 15972 17276 15978
rect 17224 15914 17276 15920
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17236 15094 17264 15438
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17328 14550 17356 19790
rect 17512 18426 17540 22063
rect 17788 20058 17816 22320
rect 18248 20058 18276 22320
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17972 19514 18000 19858
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 18708 19394 18736 22320
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 18524 19366 18736 19394
rect 18972 19372 19024 19378
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17512 17082 17540 17478
rect 17604 17241 17632 19110
rect 17774 18864 17830 18873
rect 17880 18834 17908 19314
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17774 18799 17830 18808
rect 17868 18828 17920 18834
rect 17788 18426 17816 18799
rect 17868 18770 17920 18776
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17880 18290 17908 18770
rect 17972 18426 18000 19110
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18236 18352 18288 18358
rect 18234 18320 18236 18329
rect 18288 18320 18290 18329
rect 17868 18284 17920 18290
rect 18234 18255 18290 18264
rect 17868 18226 17920 18232
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 18064 17746 18092 18090
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17590 17232 17646 17241
rect 17972 17202 18000 17614
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17590 17167 17646 17176
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17408 17060 17460 17066
rect 17512 17054 17632 17082
rect 17408 17002 17460 17008
rect 17420 16794 17448 17002
rect 17604 16998 17632 17054
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17866 16960 17922 16969
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17512 15706 17540 16934
rect 17866 16895 17922 16904
rect 17880 16658 17908 16895
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17972 16114 18000 17138
rect 18524 16794 18552 19366
rect 19168 19360 19196 22320
rect 19246 21176 19302 21185
rect 19246 21111 19302 21120
rect 18972 19314 19024 19320
rect 19076 19332 19196 19360
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18616 18086 18644 18119
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17377 18644 17478
rect 18602 17368 18658 17377
rect 18602 17303 18658 17312
rect 18708 16794 18736 19246
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18800 18222 18828 18770
rect 18880 18692 18932 18698
rect 18984 18680 19012 19314
rect 18932 18652 19012 18680
rect 18880 18634 18932 18640
rect 18878 18456 18934 18465
rect 18878 18391 18880 18400
rect 18932 18391 18934 18400
rect 18880 18362 18932 18368
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18788 18216 18840 18222
rect 18892 18193 18920 18226
rect 18788 18158 18840 18164
rect 18878 18184 18934 18193
rect 18878 18119 18934 18128
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18800 16182 18828 18022
rect 18878 17912 18934 17921
rect 18878 17847 18934 17856
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17592 15632 17644 15638
rect 17592 15574 17644 15580
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17316 14544 17368 14550
rect 17316 14486 17368 14492
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17236 13394 17264 14350
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17236 12986 17264 13330
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17236 12306 17264 12922
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16776 10606 16804 11018
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16868 10742 16896 10950
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16960 10674 16988 10950
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 17144 10010 17172 11630
rect 17420 10690 17448 13874
rect 17512 13530 17540 14758
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17328 10662 17448 10690
rect 17144 9982 17264 10010
rect 16488 9648 16540 9654
rect 16486 9616 16488 9625
rect 16540 9616 16542 9625
rect 16486 9551 16542 9560
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16960 9110 16988 9318
rect 16948 9104 17000 9110
rect 16948 9046 17000 9052
rect 17236 8906 17264 9982
rect 17328 9926 17356 10662
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17420 9586 17448 10474
rect 17604 10146 17632 15574
rect 17696 13530 17724 15982
rect 17866 15600 17922 15609
rect 17866 15535 17922 15544
rect 17774 15056 17830 15065
rect 17774 14991 17830 15000
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17696 12986 17724 13330
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17788 11898 17816 14991
rect 17880 14890 17908 15535
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18708 14958 18736 16050
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18328 14952 18380 14958
rect 18326 14920 18328 14929
rect 18604 14952 18656 14958
rect 18380 14920 18382 14929
rect 17868 14884 17920 14890
rect 18604 14894 18656 14900
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18326 14855 18382 14864
rect 17868 14826 17920 14832
rect 18616 14482 18644 14894
rect 18708 14550 18736 14894
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 12374 17908 14214
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18418 13968 18474 13977
rect 18418 13903 18474 13912
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17972 12986 18000 13806
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 18064 13462 18092 13670
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 18432 13394 18460 13903
rect 18524 13530 18552 14418
rect 18602 14104 18658 14113
rect 18602 14039 18658 14048
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18420 13388 18472 13394
rect 18472 13348 18552 13376
rect 18420 13330 18472 13336
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12986 18552 13348
rect 18616 13190 18644 14039
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17972 11898 18000 12650
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18708 11694 18736 13942
rect 18800 13530 18828 15506
rect 18892 15094 18920 17847
rect 18984 17814 19012 18652
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 19076 16250 19104 19332
rect 19154 19272 19210 19281
rect 19154 19207 19210 19216
rect 19168 18426 19196 19207
rect 19260 19174 19288 21111
rect 19628 19904 19656 22320
rect 20180 20346 20208 22320
rect 20640 21706 20668 22320
rect 20548 21678 20668 21706
rect 20442 20632 20498 20641
rect 20442 20567 20498 20576
rect 20088 20318 20208 20346
rect 19892 19916 19944 19922
rect 19628 19876 19748 19904
rect 19614 19816 19670 19825
rect 19614 19751 19616 19760
rect 19668 19751 19670 19760
rect 19616 19722 19668 19728
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19260 15706 19288 18770
rect 19352 17626 19380 19178
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19444 17814 19472 18158
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19352 17598 19472 17626
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19352 17134 19380 17478
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19444 16658 19472 17598
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19536 15978 19564 18702
rect 19720 18086 19748 19876
rect 19892 19858 19944 19864
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19812 18290 19840 19790
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19628 16590 19656 17206
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19812 16658 19840 17002
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19628 16046 19656 16526
rect 19904 16454 19932 19858
rect 19996 19446 20024 19858
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 20088 18902 20116 20318
rect 20166 20224 20222 20233
rect 20166 20159 20222 20168
rect 20180 20058 20208 20159
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20076 18896 20128 18902
rect 20076 18838 20128 18844
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19996 18737 20024 18770
rect 19982 18728 20038 18737
rect 19982 18663 20038 18672
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19996 17338 20024 17682
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16726 20116 16934
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 20180 16590 20208 17070
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19064 15632 19116 15638
rect 19064 15574 19116 15580
rect 18880 15088 18932 15094
rect 18880 15030 18932 15036
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18892 13530 18920 14486
rect 18970 13696 19026 13705
rect 18970 13631 19026 13640
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18800 12918 18828 13194
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18800 12442 18828 12854
rect 18892 12782 18920 13126
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18800 11762 18828 12378
rect 18984 12288 19012 13631
rect 19076 13297 19104 15574
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 19062 13288 19118 13297
rect 19062 13223 19118 13232
rect 18892 12260 19012 12288
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11393 18460 11494
rect 18418 11384 18474 11393
rect 17776 11348 17828 11354
rect 18418 11319 18474 11328
rect 17776 11290 17828 11296
rect 17788 11257 17816 11290
rect 17774 11248 17830 11257
rect 17774 11183 17830 11192
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17788 10266 17816 11086
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10606 18000 10950
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18432 10470 18460 10542
rect 18616 10538 18644 11154
rect 18892 10810 18920 12260
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 18052 10192 18104 10198
rect 17500 10124 17552 10130
rect 17604 10118 18000 10146
rect 18052 10134 18104 10140
rect 17500 10066 17552 10072
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17512 9178 17540 10066
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16684 8090 16712 8298
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16776 7546 16804 8230
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15948 6322 15976 6734
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15212 6174 15332 6202
rect 15212 6118 15240 6174
rect 16408 6118 16436 6802
rect 16592 6730 16620 7142
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16684 6458 16712 7142
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16868 6118 16896 7890
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 6254 16988 7686
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17052 6322 17080 6734
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15212 5778 15240 6054
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 17236 5166 17264 8842
rect 17420 7818 17448 8978
rect 17512 8498 17540 9114
rect 17972 9081 18000 10118
rect 18064 10033 18092 10134
rect 18340 10130 18368 10406
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18050 10024 18106 10033
rect 18050 9959 18106 9968
rect 18432 9908 18460 10406
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18432 9880 18552 9908
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18524 9568 18552 9880
rect 18432 9540 18644 9568
rect 18432 9382 18460 9540
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 17774 9072 17830 9081
rect 17958 9072 18014 9081
rect 17868 9036 17920 9042
rect 17830 9016 17868 9024
rect 17774 9007 17868 9016
rect 17788 8996 17868 9007
rect 17958 9007 18014 9016
rect 17868 8978 17920 8984
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17420 7410 17448 7754
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14186 2544 14242 2553
rect 14186 2479 14242 2488
rect 14096 2100 14148 2106
rect 14096 2042 14148 2048
rect 17880 1057 17908 8978
rect 18524 8974 18552 9386
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18524 8634 18552 8910
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18616 8498 18644 9540
rect 18708 9466 18736 10066
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18892 9722 18920 9998
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 18708 9438 18828 9466
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 8906 18736 9318
rect 18800 9042 18828 9438
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 7954 18644 8434
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 17972 7546 18000 7890
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18340 6934 18368 7346
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18144 6792 18196 6798
rect 18142 6760 18144 6769
rect 18196 6760 18198 6769
rect 17972 6718 18142 6746
rect 17972 6390 18000 6718
rect 18524 6730 18552 7890
rect 18602 7576 18658 7585
rect 18602 7511 18658 7520
rect 18616 7002 18644 7511
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18142 6695 18198 6704
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 18142 6216 18198 6225
rect 18052 6180 18104 6186
rect 18142 6151 18198 6160
rect 18052 6122 18104 6128
rect 17960 5840 18012 5846
rect 18064 5817 18092 6122
rect 17960 5782 18012 5788
rect 18050 5808 18106 5817
rect 17972 5273 18000 5782
rect 18156 5778 18184 6151
rect 18050 5743 18106 5752
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 18524 4865 18552 5306
rect 18510 4856 18566 4865
rect 18510 4791 18566 4800
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17972 3505 18000 4082
rect 17958 3496 18014 3505
rect 17958 3431 18014 3440
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18512 2100 18564 2106
rect 18512 2042 18564 2048
rect 18524 1601 18552 2042
rect 18510 1592 18566 1601
rect 18510 1527 18566 1536
rect 17866 1048 17922 1057
rect 17866 983 17922 992
rect 13266 640 13322 649
rect 13266 575 13322 584
rect 5264 332 5316 338
rect 5264 274 5316 280
rect 11334 0 11390 480
rect 18800 241 18828 8978
rect 18892 2009 18920 9658
rect 18984 8537 19012 12106
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19076 10470 19104 11630
rect 19168 10810 19196 15370
rect 19260 14618 19288 15438
rect 19352 14618 19380 15506
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19444 14074 19472 15438
rect 19536 14822 19564 15438
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19260 12753 19288 13670
rect 19246 12744 19302 12753
rect 19246 12679 19302 12688
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19260 10656 19288 11290
rect 19168 10628 19288 10656
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19076 9353 19104 9862
rect 19062 9344 19118 9353
rect 19062 9279 19118 9288
rect 18970 8528 19026 8537
rect 18970 8463 19026 8472
rect 19076 8072 19104 9279
rect 18984 8044 19104 8072
rect 18984 7290 19012 8044
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19076 7410 19104 7890
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 18984 7262 19104 7290
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18878 2000 18934 2009
rect 18878 1935 18934 1944
rect 18984 480 19012 3538
rect 19076 2961 19104 7262
rect 19168 7177 19196 10628
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 10062 19288 10406
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9654 19288 9998
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19260 8974 19288 9590
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19352 8430 19380 13806
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19444 13433 19472 13670
rect 19430 13424 19486 13433
rect 19430 13359 19486 13368
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12782 19472 13262
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 9994 19472 12174
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19260 8294 19288 8325
rect 19248 8288 19300 8294
rect 19444 8242 19472 9386
rect 19300 8236 19472 8242
rect 19248 8230 19472 8236
rect 19260 8214 19472 8230
rect 19154 7168 19210 7177
rect 19154 7103 19210 7112
rect 19260 3913 19288 8214
rect 19536 8022 19564 14758
rect 19628 12442 19656 15506
rect 19812 13802 19840 15914
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20088 14550 20116 15302
rect 20180 14890 20208 15846
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20180 14414 20208 14826
rect 20272 14618 20300 15438
rect 20364 15366 20392 19246
rect 20456 18970 20484 20567
rect 20548 19009 20576 21678
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20640 20058 20668 21519
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20732 19174 20760 22471
rect 21086 22320 21142 22800
rect 21546 22320 21602 22800
rect 22006 22320 22062 22800
rect 22466 22320 22522 22800
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20534 19000 20590 19009
rect 20444 18964 20496 18970
rect 20534 18935 20590 18944
rect 20444 18906 20496 18912
rect 21100 18465 21128 22320
rect 21560 18834 21588 22320
rect 22020 19145 22048 22320
rect 22006 19136 22062 19145
rect 22006 19071 22062 19080
rect 22480 18902 22508 22320
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21086 18456 21142 18465
rect 21086 18391 21142 18400
rect 20904 18352 20956 18358
rect 20902 18320 20904 18329
rect 20956 18320 20958 18329
rect 20902 18255 20958 18264
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20456 17066 20484 17818
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20180 13938 20208 14350
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 20272 13530 20300 14418
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19720 11354 19748 12242
rect 19892 12164 19944 12170
rect 19996 12152 20024 12922
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 20088 12322 20116 12650
rect 20180 12442 20208 13330
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20088 12294 20208 12322
rect 20180 12238 20208 12294
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 19944 12124 20024 12152
rect 19892 12106 19944 12112
rect 20180 11898 20208 12174
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 19892 11620 19944 11626
rect 19892 11562 19944 11568
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19904 11082 19932 11562
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19904 10810 19932 11018
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19720 10198 19748 10406
rect 19904 10198 19932 10746
rect 19708 10192 19760 10198
rect 19708 10134 19760 10140
rect 19892 10192 19944 10198
rect 19892 10134 19944 10140
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19812 6730 19840 8978
rect 19904 8906 19932 9998
rect 19996 9654 20024 11086
rect 20088 10810 20116 11154
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 20180 9489 20208 11222
rect 20166 9480 20222 9489
rect 20166 9415 20222 9424
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 20364 8129 20392 13670
rect 20456 12345 20484 17002
rect 20732 16522 20760 18158
rect 20994 16552 21050 16561
rect 20720 16516 20772 16522
rect 20994 16487 21050 16496
rect 20720 16458 20772 16464
rect 20626 14648 20682 14657
rect 20626 14583 20682 14592
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20548 13938 20576 14282
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20442 12336 20498 12345
rect 20442 12271 20498 12280
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20548 9586 20576 10610
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20640 8634 20668 14583
rect 21008 11898 21036 16487
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 10266 20760 10406
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20350 8120 20406 8129
rect 20350 8055 20406 8064
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20180 7002 20208 7822
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20364 7274 20392 7686
rect 20456 7546 20484 8298
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20352 7268 20404 7274
rect 20352 7210 20404 7216
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19800 6724 19852 6730
rect 19800 6666 19852 6672
rect 20088 6458 20116 6734
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20364 6322 20392 7210
rect 20456 6798 20484 7482
rect 20824 7342 20852 11630
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 19904 5914 19932 6054
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 20548 4321 20576 6054
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 19246 3904 19302 3913
rect 19246 3839 19302 3848
rect 19062 2952 19118 2961
rect 19062 2887 19118 2896
rect 18786 232 18842 241
rect 18786 167 18842 176
rect 18970 0 19026 480
<< via2 >>
rect 2778 22480 2834 22536
rect 1950 19760 2006 19816
rect 1950 19216 2006 19272
rect 20718 22480 20774 22536
rect 2962 22072 3018 22128
rect 2870 21120 2926 21176
rect 2134 19216 2190 19272
rect 1582 18944 1638 19000
rect 1766 18808 1822 18864
rect 2502 18808 2558 18864
rect 2134 17740 2190 17776
rect 2134 17720 2136 17740
rect 2136 17720 2188 17740
rect 2188 17720 2190 17740
rect 1766 17312 1822 17368
rect 1950 16940 1952 16960
rect 1952 16940 2004 16960
rect 2004 16940 2006 16960
rect 1950 16904 2006 16940
rect 1582 16632 1638 16688
rect 1582 16516 1638 16552
rect 1582 16496 1584 16516
rect 1584 16496 1636 16516
rect 1636 16496 1638 16516
rect 2778 19216 2834 19272
rect 3054 18264 3110 18320
rect 2778 17856 2834 17912
rect 1950 15544 2006 15600
rect 1950 15036 1952 15056
rect 1952 15036 2004 15056
rect 2004 15036 2006 15056
rect 1950 15000 2006 15036
rect 1582 14592 1638 14648
rect 1858 14048 1914 14104
rect 1490 11328 1546 11384
rect 2410 11600 2466 11656
rect 2778 9560 2834 9616
rect 3422 19080 3478 19136
rect 3422 18708 3424 18728
rect 3424 18708 3476 18728
rect 3476 18708 3478 18728
rect 3422 18672 3478 18708
rect 3882 21528 3938 21584
rect 3698 20576 3754 20632
rect 3790 20168 3846 20224
rect 3790 19352 3846 19408
rect 3606 19216 3662 19272
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 3514 15952 3570 16008
rect 3606 13640 3662 13696
rect 3238 13232 3294 13288
rect 3606 12688 3662 12744
rect 3974 16496 4030 16552
rect 5262 19352 5318 19408
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4618 17620 4620 17640
rect 4620 17620 4672 17640
rect 4672 17620 4674 17640
rect 4618 17584 4674 17620
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4894 17076 4896 17096
rect 4896 17076 4948 17096
rect 4948 17076 4950 17096
rect 4894 17040 4950 17076
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3422 11056 3478 11112
rect 2962 5752 3018 5808
rect 3146 4800 3202 4856
rect 4066 10804 4122 10840
rect 4066 10784 4068 10804
rect 4068 10784 4120 10804
rect 4120 10784 4122 10804
rect 4066 10376 4122 10432
rect 3974 9968 4030 10024
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 5538 17720 5594 17776
rect 5630 16360 5686 16416
rect 5906 16496 5962 16552
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4250 10240 4306 10296
rect 4250 10104 4306 10160
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4250 9152 4306 9208
rect 4066 8472 4122 8528
rect 3790 7520 3846 7576
rect 3330 3848 3386 3904
rect 2778 1944 2834 2000
rect 3330 1536 3386 1592
rect 938 992 994 1048
rect 3146 584 3202 640
rect 4066 8064 4122 8120
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4066 7112 4122 7168
rect 4066 6724 4122 6760
rect 4066 6704 4068 6724
rect 4068 6704 4120 6724
rect 4120 6704 4122 6724
rect 3974 6160 4030 6216
rect 4066 5228 4122 5264
rect 4066 5208 4068 5228
rect 4068 5208 4120 5228
rect 4120 5208 4122 5228
rect 4066 4256 4122 4312
rect 3882 3440 3938 3496
rect 4066 2896 4122 2952
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4250 2488 4306 2544
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 3330 176 3386 232
rect 5722 11772 5724 11792
rect 5724 11772 5776 11792
rect 5776 11772 5778 11792
rect 5722 11736 5778 11772
rect 7102 18944 7158 19000
rect 7378 19080 7434 19136
rect 7010 17040 7066 17096
rect 7194 17584 7250 17640
rect 6090 10512 6146 10568
rect 5906 9016 5962 9072
rect 6826 11872 6882 11928
rect 7102 13368 7158 13424
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 8206 11600 8262 11656
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8850 17584 8906 17640
rect 8758 16632 8814 16688
rect 8666 12316 8668 12336
rect 8668 12316 8720 12336
rect 8720 12316 8722 12336
rect 8666 12280 8722 12316
rect 8850 11600 8906 11656
rect 9586 16396 9588 16416
rect 9588 16396 9640 16416
rect 9640 16396 9642 16416
rect 9586 16360 9642 16396
rect 9954 18264 10010 18320
rect 9954 17756 9956 17776
rect 9956 17756 10008 17776
rect 10008 17756 10010 17776
rect 9954 17720 10010 17756
rect 10414 19080 10470 19136
rect 10230 18672 10286 18728
rect 9954 15580 9956 15600
rect 9956 15580 10008 15600
rect 10008 15580 10010 15600
rect 9954 15544 10010 15580
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 10506 18672 10562 18728
rect 10414 17176 10470 17232
rect 9494 12008 9550 12064
rect 9310 11872 9366 11928
rect 9402 11756 9458 11792
rect 9402 11736 9404 11756
rect 9404 11736 9456 11756
rect 9456 11736 9458 11756
rect 9126 11056 9182 11112
rect 8574 10512 8630 10568
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 10322 13912 10378 13968
rect 10230 13232 10286 13288
rect 10046 9152 10102 9208
rect 10322 9152 10378 9208
rect 10966 17856 11022 17912
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11702 18400 11758 18456
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 10874 13504 10930 13560
rect 10966 10648 11022 10704
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11610 16088 11666 16144
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 12070 19080 12126 19136
rect 12346 17040 12402 17096
rect 11886 13776 11942 13832
rect 11518 10548 11520 10568
rect 11520 10548 11572 10568
rect 11572 10548 11574 10568
rect 11518 10512 11574 10548
rect 11794 9968 11850 10024
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 12898 17992 12954 18048
rect 12622 17040 12678 17096
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 12438 15580 12440 15600
rect 12440 15580 12492 15600
rect 12492 15580 12494 15600
rect 12438 15544 12494 15580
rect 12622 15408 12678 15464
rect 12346 14864 12402 14920
rect 12806 13504 12862 13560
rect 12346 13232 12402 13288
rect 12714 13232 12770 13288
rect 12990 16108 13046 16144
rect 12990 16088 12992 16108
rect 12992 16088 13044 16108
rect 13044 16088 13046 16108
rect 12254 11192 12310 11248
rect 12254 9152 12310 9208
rect 12162 8608 12218 8664
rect 10874 7812 10930 7848
rect 10874 7792 10876 7812
rect 10876 7792 10928 7812
rect 10928 7792 10930 7812
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11610 6976 11666 7032
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 12070 7812 12126 7848
rect 12070 7792 12072 7812
rect 12072 7792 12124 7812
rect 12124 7792 12126 7812
rect 12806 10648 12862 10704
rect 12530 9036 12586 9072
rect 12530 9016 12532 9036
rect 12532 9016 12584 9036
rect 12584 9016 12586 9036
rect 12438 8608 12494 8664
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 13266 15000 13322 15056
rect 12990 9016 13046 9072
rect 13082 8880 13138 8936
rect 13818 17856 13874 17912
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14646 18708 14648 18728
rect 14648 18708 14700 18728
rect 14700 18708 14702 18728
rect 14646 18672 14702 18708
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14462 17876 14518 17912
rect 14462 17856 14464 17876
rect 14464 17856 14516 17876
rect 14516 17856 14518 17876
rect 15106 17756 15108 17776
rect 15108 17756 15160 17776
rect 15160 17756 15162 17776
rect 15106 17720 15162 17756
rect 14554 17040 14610 17096
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14554 16496 14610 16552
rect 14278 15428 14334 15464
rect 14278 15408 14280 15428
rect 14280 15408 14332 15428
rect 14332 15408 14334 15428
rect 13818 9288 13874 9344
rect 13726 9152 13782 9208
rect 13634 6996 13690 7032
rect 13634 6976 13636 6996
rect 13636 6976 13688 6996
rect 13688 6976 13690 6996
rect 14278 10376 14334 10432
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 15014 15544 15070 15600
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14646 14320 14702 14376
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 15658 18400 15714 18456
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14186 8916 14188 8936
rect 14188 8916 14240 8936
rect 14240 8916 14242 8936
rect 14186 8880 14242 8916
rect 14738 9560 14794 9616
rect 14922 9424 14978 9480
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 15474 9560 15530 9616
rect 16118 18536 16174 18592
rect 15842 15020 15898 15056
rect 15842 15000 15844 15020
rect 15844 15000 15896 15020
rect 15896 15000 15898 15020
rect 15750 11056 15806 11112
rect 16210 17584 16266 17640
rect 16302 15952 16358 16008
rect 17498 22072 17554 22128
rect 16302 10512 16358 10568
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 16854 13776 16910 13832
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17774 18808 17830 18864
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18234 18300 18236 18320
rect 18236 18300 18288 18320
rect 18288 18300 18290 18320
rect 18234 18264 18290 18300
rect 17590 17176 17646 17232
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17866 16904 17922 16960
rect 19246 21120 19302 21176
rect 18602 18128 18658 18184
rect 18602 17312 18658 17368
rect 18878 18420 18934 18456
rect 18878 18400 18880 18420
rect 18880 18400 18932 18420
rect 18932 18400 18934 18420
rect 18878 18128 18934 18184
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18878 17856 18934 17912
rect 16486 9596 16488 9616
rect 16488 9596 16540 9616
rect 16540 9596 16542 9616
rect 16486 9560 16542 9596
rect 17866 15544 17922 15600
rect 17774 15000 17830 15056
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18326 14900 18328 14920
rect 18328 14900 18380 14920
rect 18380 14900 18382 14920
rect 18326 14864 18382 14900
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18418 13912 18474 13968
rect 18602 14048 18658 14104
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 19154 19216 19210 19272
rect 20442 20576 20498 20632
rect 19614 19780 19670 19816
rect 19614 19760 19616 19780
rect 19616 19760 19668 19780
rect 19668 19760 19670 19780
rect 20166 20168 20222 20224
rect 19982 18672 20038 18728
rect 18970 13640 19026 13696
rect 19062 13232 19118 13288
rect 18418 11328 18474 11384
rect 17774 11192 17830 11248
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 18050 9968 18106 10024
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17774 9016 17830 9072
rect 17958 9016 18014 9072
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 14186 2488 14242 2544
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18142 6740 18144 6760
rect 18144 6740 18196 6760
rect 18196 6740 18198 6760
rect 18142 6704 18198 6740
rect 18602 7520 18658 7576
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18142 6160 18198 6216
rect 18050 5752 18106 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 17958 5208 18014 5264
rect 18510 4800 18566 4856
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17958 3440 18014 3496
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18510 1536 18566 1592
rect 17866 992 17922 1048
rect 13266 584 13322 640
rect 19246 12688 19302 12744
rect 19062 9288 19118 9344
rect 18970 8472 19026 8528
rect 18878 1944 18934 2000
rect 19430 13368 19486 13424
rect 19154 7112 19210 7168
rect 20626 21528 20682 21584
rect 20534 18944 20590 19000
rect 22006 19080 22062 19136
rect 21086 18400 21142 18456
rect 20902 18300 20904 18320
rect 20904 18300 20956 18320
rect 20956 18300 20958 18320
rect 20902 18264 20958 18300
rect 20166 9424 20222 9480
rect 20994 16496 21050 16552
rect 20626 14592 20682 14648
rect 20442 12280 20498 12336
rect 20350 8064 20406 8120
rect 20534 4256 20590 4312
rect 19246 3848 19302 3904
rect 19062 2896 19118 2952
rect 18786 176 18842 232
<< metal3 >>
rect 0 22538 480 22568
rect 2773 22538 2839 22541
rect 0 22536 2839 22538
rect 0 22480 2778 22536
rect 2834 22480 2839 22536
rect 0 22478 2839 22480
rect 0 22448 480 22478
rect 2773 22475 2839 22478
rect 20713 22538 20779 22541
rect 22320 22538 22800 22568
rect 20713 22536 22800 22538
rect 20713 22480 20718 22536
rect 20774 22480 22800 22536
rect 20713 22478 22800 22480
rect 20713 22475 20779 22478
rect 22320 22448 22800 22478
rect 0 22130 480 22160
rect 2957 22130 3023 22133
rect 0 22128 3023 22130
rect 0 22072 2962 22128
rect 3018 22072 3023 22128
rect 0 22070 3023 22072
rect 0 22040 480 22070
rect 2957 22067 3023 22070
rect 17493 22130 17559 22133
rect 22320 22130 22800 22160
rect 17493 22128 22800 22130
rect 17493 22072 17498 22128
rect 17554 22072 22800 22128
rect 17493 22070 22800 22072
rect 17493 22067 17559 22070
rect 22320 22040 22800 22070
rect 0 21586 480 21616
rect 3877 21586 3943 21589
rect 0 21584 3943 21586
rect 0 21528 3882 21584
rect 3938 21528 3943 21584
rect 0 21526 3943 21528
rect 0 21496 480 21526
rect 3877 21523 3943 21526
rect 20621 21586 20687 21589
rect 22320 21586 22800 21616
rect 20621 21584 22800 21586
rect 20621 21528 20626 21584
rect 20682 21528 22800 21584
rect 20621 21526 22800 21528
rect 20621 21523 20687 21526
rect 22320 21496 22800 21526
rect 0 21178 480 21208
rect 2865 21178 2931 21181
rect 0 21176 2931 21178
rect 0 21120 2870 21176
rect 2926 21120 2931 21176
rect 0 21118 2931 21120
rect 0 21088 480 21118
rect 2865 21115 2931 21118
rect 19241 21178 19307 21181
rect 22320 21178 22800 21208
rect 19241 21176 22800 21178
rect 19241 21120 19246 21176
rect 19302 21120 22800 21176
rect 19241 21118 22800 21120
rect 19241 21115 19307 21118
rect 22320 21088 22800 21118
rect 0 20634 480 20664
rect 3693 20634 3759 20637
rect 0 20632 3759 20634
rect 0 20576 3698 20632
rect 3754 20576 3759 20632
rect 0 20574 3759 20576
rect 0 20544 480 20574
rect 3693 20571 3759 20574
rect 20437 20634 20503 20637
rect 22320 20634 22800 20664
rect 20437 20632 22800 20634
rect 20437 20576 20442 20632
rect 20498 20576 22800 20632
rect 20437 20574 22800 20576
rect 20437 20571 20503 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 3785 20226 3851 20229
rect 0 20224 3851 20226
rect 0 20168 3790 20224
rect 3846 20168 3851 20224
rect 0 20166 3851 20168
rect 0 20136 480 20166
rect 3785 20163 3851 20166
rect 20161 20226 20227 20229
rect 22320 20226 22800 20256
rect 20161 20224 22800 20226
rect 20161 20168 20166 20224
rect 20222 20168 22800 20224
rect 20161 20166 22800 20168
rect 20161 20163 20227 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 480 19758
rect 1945 19755 2011 19758
rect 19609 19818 19675 19821
rect 22320 19818 22800 19848
rect 19609 19816 22800 19818
rect 19609 19760 19614 19816
rect 19670 19760 22800 19816
rect 19609 19758 22800 19760
rect 19609 19755 19675 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 3785 19410 3851 19413
rect 5257 19410 5323 19413
rect 3785 19408 5323 19410
rect 3785 19352 3790 19408
rect 3846 19352 5262 19408
rect 5318 19352 5323 19408
rect 3785 19350 5323 19352
rect 3785 19347 3851 19350
rect 5257 19347 5323 19350
rect 0 19274 480 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 480 19214
rect 1945 19211 2011 19214
rect 2129 19274 2195 19277
rect 2773 19274 2839 19277
rect 2129 19272 2839 19274
rect 2129 19216 2134 19272
rect 2190 19216 2778 19272
rect 2834 19216 2839 19272
rect 2129 19214 2839 19216
rect 2129 19211 2195 19214
rect 2773 19211 2839 19214
rect 3601 19274 3667 19277
rect 19149 19274 19215 19277
rect 22320 19274 22800 19304
rect 3601 19272 17234 19274
rect 3601 19216 3606 19272
rect 3662 19216 17234 19272
rect 3601 19214 17234 19216
rect 3601 19211 3667 19214
rect 3417 19138 3483 19141
rect 7373 19138 7439 19141
rect 3417 19136 7439 19138
rect 3417 19080 3422 19136
rect 3478 19080 7378 19136
rect 7434 19080 7439 19136
rect 3417 19078 7439 19080
rect 3417 19075 3483 19078
rect 7373 19075 7439 19078
rect 10409 19138 10475 19141
rect 12065 19138 12131 19141
rect 10409 19136 12131 19138
rect 10409 19080 10414 19136
rect 10470 19080 12070 19136
rect 12126 19080 12131 19136
rect 10409 19078 12131 19080
rect 17174 19138 17234 19214
rect 19149 19272 22800 19274
rect 19149 19216 19154 19272
rect 19210 19216 22800 19272
rect 19149 19214 22800 19216
rect 19149 19211 19215 19214
rect 22320 19184 22800 19214
rect 22001 19138 22067 19141
rect 17174 19136 22067 19138
rect 17174 19080 22006 19136
rect 22062 19080 22067 19136
rect 17174 19078 22067 19080
rect 10409 19075 10475 19078
rect 12065 19075 12131 19078
rect 22001 19075 22067 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 1577 19002 1643 19005
rect 7097 19002 7163 19005
rect 20529 19002 20595 19005
rect 1577 19000 7163 19002
rect 1577 18944 1582 19000
rect 1638 18944 7102 19000
rect 7158 18944 7163 19000
rect 1577 18942 7163 18944
rect 1577 18939 1643 18942
rect 7097 18939 7163 18942
rect 16438 19000 20595 19002
rect 16438 18944 20534 19000
rect 20590 18944 20595 19000
rect 16438 18942 20595 18944
rect 0 18866 480 18896
rect 1761 18866 1827 18869
rect 0 18864 1827 18866
rect 0 18808 1766 18864
rect 1822 18808 1827 18864
rect 0 18806 1827 18808
rect 0 18776 480 18806
rect 1761 18803 1827 18806
rect 2497 18866 2563 18869
rect 16438 18866 16498 18942
rect 20529 18939 20595 18942
rect 2497 18864 16498 18866
rect 2497 18808 2502 18864
rect 2558 18808 16498 18864
rect 2497 18806 16498 18808
rect 17769 18866 17835 18869
rect 22320 18866 22800 18896
rect 17769 18864 22800 18866
rect 17769 18808 17774 18864
rect 17830 18808 22800 18864
rect 17769 18806 22800 18808
rect 2497 18803 2563 18806
rect 17769 18803 17835 18806
rect 22320 18776 22800 18806
rect 3417 18730 3483 18733
rect 10225 18730 10291 18733
rect 3417 18728 10291 18730
rect 3417 18672 3422 18728
rect 3478 18672 10230 18728
rect 10286 18672 10291 18728
rect 3417 18670 10291 18672
rect 3417 18667 3483 18670
rect 10225 18667 10291 18670
rect 10501 18730 10567 18733
rect 10501 18728 11714 18730
rect 10501 18672 10506 18728
rect 10562 18672 11714 18728
rect 10501 18670 11714 18672
rect 10501 18667 10567 18670
rect 11654 18594 11714 18670
rect 12934 18668 12940 18732
rect 13004 18730 13010 18732
rect 14641 18730 14707 18733
rect 19977 18730 20043 18733
rect 13004 18728 20043 18730
rect 13004 18672 14646 18728
rect 14702 18672 19982 18728
rect 20038 18672 20043 18728
rect 13004 18670 20043 18672
rect 13004 18668 13010 18670
rect 14641 18667 14707 18670
rect 19977 18667 20043 18670
rect 16113 18594 16179 18597
rect 11654 18592 16179 18594
rect 11654 18536 16118 18592
rect 16174 18536 16179 18592
rect 11654 18534 16179 18536
rect 16113 18531 16179 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 11697 18458 11763 18461
rect 15653 18458 15719 18461
rect 11697 18456 15719 18458
rect 11697 18400 11702 18456
rect 11758 18400 15658 18456
rect 15714 18400 15719 18456
rect 11697 18398 15719 18400
rect 11697 18395 11763 18398
rect 15653 18395 15719 18398
rect 18873 18458 18939 18461
rect 21081 18458 21147 18461
rect 18873 18456 21147 18458
rect 18873 18400 18878 18456
rect 18934 18400 21086 18456
rect 21142 18400 21147 18456
rect 18873 18398 21147 18400
rect 18873 18395 18939 18398
rect 21081 18395 21147 18398
rect 0 18322 480 18352
rect 3049 18322 3115 18325
rect 0 18320 3115 18322
rect 0 18264 3054 18320
rect 3110 18264 3115 18320
rect 0 18262 3115 18264
rect 0 18232 480 18262
rect 3049 18259 3115 18262
rect 9949 18322 10015 18325
rect 18229 18322 18295 18325
rect 9949 18320 18295 18322
rect 9949 18264 9954 18320
rect 10010 18264 18234 18320
rect 18290 18264 18295 18320
rect 9949 18262 18295 18264
rect 9949 18259 10015 18262
rect 18229 18259 18295 18262
rect 20897 18322 20963 18325
rect 22320 18322 22800 18352
rect 20897 18320 22800 18322
rect 20897 18264 20902 18320
rect 20958 18264 22800 18320
rect 20897 18262 22800 18264
rect 20897 18259 20963 18262
rect 22320 18232 22800 18262
rect 18597 18186 18663 18189
rect 18873 18186 18939 18189
rect 18597 18184 18939 18186
rect 18597 18128 18602 18184
rect 18658 18128 18878 18184
rect 18934 18128 18939 18184
rect 18597 18126 18939 18128
rect 18597 18123 18663 18126
rect 18873 18123 18939 18126
rect 12893 18050 12959 18053
rect 13118 18050 13124 18052
rect 12893 18048 13124 18050
rect 12893 17992 12898 18048
rect 12954 17992 13124 18048
rect 12893 17990 13124 17992
rect 12893 17987 12959 17990
rect 13118 17988 13124 17990
rect 13188 17988 13194 18052
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 2773 17914 2839 17917
rect 0 17912 2839 17914
rect 0 17856 2778 17912
rect 2834 17856 2839 17912
rect 0 17854 2839 17856
rect 0 17824 480 17854
rect 2773 17851 2839 17854
rect 10961 17914 11027 17917
rect 13813 17914 13879 17917
rect 14457 17914 14523 17917
rect 10961 17912 14523 17914
rect 10961 17856 10966 17912
rect 11022 17856 13818 17912
rect 13874 17856 14462 17912
rect 14518 17856 14523 17912
rect 10961 17854 14523 17856
rect 10961 17851 11027 17854
rect 13813 17851 13879 17854
rect 14457 17851 14523 17854
rect 18873 17914 18939 17917
rect 22320 17914 22800 17944
rect 18873 17912 22800 17914
rect 18873 17856 18878 17912
rect 18934 17856 22800 17912
rect 18873 17854 22800 17856
rect 18873 17851 18939 17854
rect 22320 17824 22800 17854
rect 2129 17778 2195 17781
rect 5533 17778 5599 17781
rect 2129 17776 5599 17778
rect 2129 17720 2134 17776
rect 2190 17720 5538 17776
rect 5594 17720 5599 17776
rect 2129 17718 5599 17720
rect 2129 17715 2195 17718
rect 5533 17715 5599 17718
rect 9949 17778 10015 17781
rect 15101 17778 15167 17781
rect 9949 17776 15167 17778
rect 9949 17720 9954 17776
rect 10010 17720 15106 17776
rect 15162 17720 15167 17776
rect 9949 17718 15167 17720
rect 9949 17715 10015 17718
rect 15101 17715 15167 17718
rect 4613 17642 4679 17645
rect 7189 17642 7255 17645
rect 4613 17640 7255 17642
rect 4613 17584 4618 17640
rect 4674 17584 7194 17640
rect 7250 17584 7255 17640
rect 4613 17582 7255 17584
rect 4613 17579 4679 17582
rect 7189 17579 7255 17582
rect 8845 17642 8911 17645
rect 16205 17642 16271 17645
rect 8845 17640 16271 17642
rect 8845 17584 8850 17640
rect 8906 17584 16210 17640
rect 16266 17584 16271 17640
rect 8845 17582 16271 17584
rect 8845 17579 8911 17582
rect 16205 17579 16271 17582
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1761 17370 1827 17373
rect 0 17368 1827 17370
rect 0 17312 1766 17368
rect 1822 17312 1827 17368
rect 0 17310 1827 17312
rect 0 17280 480 17310
rect 1761 17307 1827 17310
rect 18597 17370 18663 17373
rect 22320 17370 22800 17400
rect 18597 17368 22800 17370
rect 18597 17312 18602 17368
rect 18658 17312 22800 17368
rect 18597 17310 22800 17312
rect 18597 17307 18663 17310
rect 22320 17280 22800 17310
rect 10409 17234 10475 17237
rect 17585 17234 17651 17237
rect 17718 17234 17724 17236
rect 10409 17232 17724 17234
rect 10409 17176 10414 17232
rect 10470 17176 17590 17232
rect 17646 17176 17724 17232
rect 10409 17174 17724 17176
rect 10409 17171 10475 17174
rect 17585 17171 17651 17174
rect 17718 17172 17724 17174
rect 17788 17172 17794 17236
rect 4889 17098 4955 17101
rect 7005 17098 7071 17101
rect 4889 17096 7071 17098
rect 4889 17040 4894 17096
rect 4950 17040 7010 17096
rect 7066 17040 7071 17096
rect 4889 17038 7071 17040
rect 4889 17035 4955 17038
rect 7005 17035 7071 17038
rect 12341 17098 12407 17101
rect 12617 17098 12683 17101
rect 12341 17096 12683 17098
rect 12341 17040 12346 17096
rect 12402 17040 12622 17096
rect 12678 17040 12683 17096
rect 12341 17038 12683 17040
rect 12341 17035 12407 17038
rect 12617 17035 12683 17038
rect 14549 17098 14615 17101
rect 18638 17098 18644 17100
rect 14549 17096 18644 17098
rect 14549 17040 14554 17096
rect 14610 17040 18644 17096
rect 14549 17038 18644 17040
rect 14549 17035 14615 17038
rect 18638 17036 18644 17038
rect 18708 17036 18714 17100
rect 0 16962 480 16992
rect 1945 16962 2011 16965
rect 0 16960 2011 16962
rect 0 16904 1950 16960
rect 2006 16904 2011 16960
rect 0 16902 2011 16904
rect 0 16872 480 16902
rect 1945 16899 2011 16902
rect 17861 16962 17927 16965
rect 22320 16962 22800 16992
rect 17861 16960 22800 16962
rect 17861 16904 17866 16960
rect 17922 16904 22800 16960
rect 17861 16902 22800 16904
rect 17861 16899 17927 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 1577 16690 1643 16693
rect 8753 16690 8819 16693
rect 1577 16688 8819 16690
rect 1577 16632 1582 16688
rect 1638 16632 8758 16688
rect 8814 16632 8819 16688
rect 1577 16630 8819 16632
rect 1577 16627 1643 16630
rect 8753 16627 8819 16630
rect 0 16554 480 16584
rect 1577 16554 1643 16557
rect 0 16552 1643 16554
rect 0 16496 1582 16552
rect 1638 16496 1643 16552
rect 0 16494 1643 16496
rect 0 16464 480 16494
rect 1577 16491 1643 16494
rect 3969 16554 4035 16557
rect 5901 16554 5967 16557
rect 14549 16554 14615 16557
rect 3969 16552 14615 16554
rect 3969 16496 3974 16552
rect 4030 16496 5906 16552
rect 5962 16496 14554 16552
rect 14610 16496 14615 16552
rect 3969 16494 14615 16496
rect 3969 16491 4035 16494
rect 5901 16491 5967 16494
rect 14549 16491 14615 16494
rect 20989 16554 21055 16557
rect 22320 16554 22800 16584
rect 20989 16552 22800 16554
rect 20989 16496 20994 16552
rect 21050 16496 22800 16552
rect 20989 16494 22800 16496
rect 20989 16491 21055 16494
rect 22320 16464 22800 16494
rect 5625 16418 5691 16421
rect 9581 16418 9647 16421
rect 5625 16416 9647 16418
rect 5625 16360 5630 16416
rect 5686 16360 9586 16416
rect 9642 16360 9647 16416
rect 5625 16358 9647 16360
rect 5625 16355 5691 16358
rect 9581 16355 9647 16358
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 11605 16146 11671 16149
rect 12985 16146 13051 16149
rect 11605 16144 13051 16146
rect 11605 16088 11610 16144
rect 11666 16088 12990 16144
rect 13046 16088 13051 16144
rect 11605 16086 13051 16088
rect 11605 16083 11671 16086
rect 12985 16083 13051 16086
rect 0 16010 480 16040
rect 3509 16010 3575 16013
rect 0 16008 3575 16010
rect 0 15952 3514 16008
rect 3570 15952 3575 16008
rect 0 15950 3575 15952
rect 0 15920 480 15950
rect 3509 15947 3575 15950
rect 16297 16010 16363 16013
rect 22320 16010 22800 16040
rect 16297 16008 22800 16010
rect 16297 15952 16302 16008
rect 16358 15952 22800 16008
rect 16297 15950 22800 15952
rect 16297 15947 16363 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 1945 15602 2011 15605
rect 0 15600 2011 15602
rect 0 15544 1950 15600
rect 2006 15544 2011 15600
rect 0 15542 2011 15544
rect 0 15512 480 15542
rect 1945 15539 2011 15542
rect 9949 15602 10015 15605
rect 12433 15602 12499 15605
rect 9949 15600 12499 15602
rect 9949 15544 9954 15600
rect 10010 15544 12438 15600
rect 12494 15544 12499 15600
rect 9949 15542 12499 15544
rect 9949 15539 10015 15542
rect 12433 15539 12499 15542
rect 15009 15602 15075 15605
rect 15142 15602 15148 15604
rect 15009 15600 15148 15602
rect 15009 15544 15014 15600
rect 15070 15544 15148 15600
rect 15009 15542 15148 15544
rect 15009 15539 15075 15542
rect 15142 15540 15148 15542
rect 15212 15540 15218 15604
rect 17861 15602 17927 15605
rect 22320 15602 22800 15632
rect 17861 15600 22800 15602
rect 17861 15544 17866 15600
rect 17922 15544 22800 15600
rect 17861 15542 22800 15544
rect 17861 15539 17927 15542
rect 22320 15512 22800 15542
rect 12617 15466 12683 15469
rect 14273 15466 14339 15469
rect 12617 15464 14339 15466
rect 12617 15408 12622 15464
rect 12678 15408 14278 15464
rect 14334 15408 14339 15464
rect 12617 15406 14339 15408
rect 12617 15403 12683 15406
rect 14273 15403 14339 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 1945 15058 2011 15061
rect 0 15056 2011 15058
rect 0 15000 1950 15056
rect 2006 15000 2011 15056
rect 0 14998 2011 15000
rect 0 14968 480 14998
rect 1945 14995 2011 14998
rect 13261 15058 13327 15061
rect 15837 15058 15903 15061
rect 13261 15056 15903 15058
rect 13261 15000 13266 15056
rect 13322 15000 15842 15056
rect 15898 15000 15903 15056
rect 13261 14998 15903 15000
rect 13261 14995 13327 14998
rect 15837 14995 15903 14998
rect 17769 15058 17835 15061
rect 22320 15058 22800 15088
rect 17769 15056 22800 15058
rect 17769 15000 17774 15056
rect 17830 15000 22800 15056
rect 17769 14998 22800 15000
rect 17769 14995 17835 14998
rect 22320 14968 22800 14998
rect 12341 14922 12407 14925
rect 18321 14922 18387 14925
rect 12341 14920 18387 14922
rect 12341 14864 12346 14920
rect 12402 14864 18326 14920
rect 18382 14864 18387 14920
rect 12341 14862 18387 14864
rect 12341 14859 12407 14862
rect 18321 14859 18387 14862
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1577 14650 1643 14653
rect 0 14648 1643 14650
rect 0 14592 1582 14648
rect 1638 14592 1643 14648
rect 0 14590 1643 14592
rect 0 14560 480 14590
rect 1577 14587 1643 14590
rect 20621 14650 20687 14653
rect 22320 14650 22800 14680
rect 20621 14648 22800 14650
rect 20621 14592 20626 14648
rect 20682 14592 22800 14648
rect 20621 14590 22800 14592
rect 20621 14587 20687 14590
rect 22320 14560 22800 14590
rect 14406 14316 14412 14380
rect 14476 14378 14482 14380
rect 14641 14378 14707 14381
rect 14476 14376 14707 14378
rect 14476 14320 14646 14376
rect 14702 14320 14707 14376
rect 14476 14318 14707 14320
rect 14476 14316 14482 14318
rect 14641 14315 14707 14318
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1853 14106 1919 14109
rect 0 14104 1919 14106
rect 0 14048 1858 14104
rect 1914 14048 1919 14104
rect 0 14046 1919 14048
rect 0 14016 480 14046
rect 1853 14043 1919 14046
rect 18597 14106 18663 14109
rect 22320 14106 22800 14136
rect 18597 14104 22800 14106
rect 18597 14048 18602 14104
rect 18658 14048 22800 14104
rect 18597 14046 22800 14048
rect 18597 14043 18663 14046
rect 22320 14016 22800 14046
rect 10317 13970 10383 13973
rect 18413 13970 18479 13973
rect 10317 13968 18479 13970
rect 10317 13912 10322 13968
rect 10378 13912 18418 13968
rect 18474 13912 18479 13968
rect 10317 13910 18479 13912
rect 10317 13907 10383 13910
rect 18413 13907 18479 13910
rect 11881 13834 11947 13837
rect 16849 13834 16915 13837
rect 11881 13832 16915 13834
rect 11881 13776 11886 13832
rect 11942 13776 16854 13832
rect 16910 13776 16915 13832
rect 11881 13774 16915 13776
rect 11881 13771 11947 13774
rect 16849 13771 16915 13774
rect 0 13698 480 13728
rect 3601 13698 3667 13701
rect 0 13696 3667 13698
rect 0 13640 3606 13696
rect 3662 13640 3667 13696
rect 0 13638 3667 13640
rect 0 13608 480 13638
rect 3601 13635 3667 13638
rect 18965 13698 19031 13701
rect 22320 13698 22800 13728
rect 18965 13696 22800 13698
rect 18965 13640 18970 13696
rect 19026 13640 22800 13696
rect 18965 13638 22800 13640
rect 18965 13635 19031 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 10869 13562 10935 13565
rect 12801 13562 12867 13565
rect 10869 13560 12867 13562
rect 10869 13504 10874 13560
rect 10930 13504 12806 13560
rect 12862 13504 12867 13560
rect 10869 13502 12867 13504
rect 10869 13499 10935 13502
rect 12801 13499 12867 13502
rect 7097 13426 7163 13429
rect 19425 13426 19491 13429
rect 7097 13424 19491 13426
rect 7097 13368 7102 13424
rect 7158 13368 19430 13424
rect 19486 13368 19491 13424
rect 7097 13366 19491 13368
rect 7097 13363 7163 13366
rect 19425 13363 19491 13366
rect 0 13290 480 13320
rect 3233 13290 3299 13293
rect 0 13288 3299 13290
rect 0 13232 3238 13288
rect 3294 13232 3299 13288
rect 0 13230 3299 13232
rect 0 13200 480 13230
rect 3233 13227 3299 13230
rect 10225 13290 10291 13293
rect 12341 13290 12407 13293
rect 10225 13288 12407 13290
rect 10225 13232 10230 13288
rect 10286 13232 12346 13288
rect 12402 13232 12407 13288
rect 10225 13230 12407 13232
rect 10225 13227 10291 13230
rect 12341 13227 12407 13230
rect 12709 13290 12775 13293
rect 14406 13290 14412 13292
rect 12709 13288 14412 13290
rect 12709 13232 12714 13288
rect 12770 13232 14412 13288
rect 12709 13230 14412 13232
rect 12709 13227 12775 13230
rect 14406 13228 14412 13230
rect 14476 13228 14482 13292
rect 19057 13290 19123 13293
rect 22320 13290 22800 13320
rect 19057 13288 22800 13290
rect 19057 13232 19062 13288
rect 19118 13232 22800 13288
rect 19057 13230 22800 13232
rect 19057 13227 19123 13230
rect 22320 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 3601 12746 3667 12749
rect 0 12744 3667 12746
rect 0 12688 3606 12744
rect 3662 12688 3667 12744
rect 0 12686 3667 12688
rect 0 12656 480 12686
rect 3601 12683 3667 12686
rect 19241 12746 19307 12749
rect 22320 12746 22800 12776
rect 19241 12744 22800 12746
rect 19241 12688 19246 12744
rect 19302 12688 22800 12744
rect 19241 12686 22800 12688
rect 19241 12683 19307 12686
rect 22320 12656 22800 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 8661 12338 8727 12341
rect 0 12336 8727 12338
rect 0 12280 8666 12336
rect 8722 12280 8727 12336
rect 0 12278 8727 12280
rect 0 12248 480 12278
rect 8661 12275 8727 12278
rect 20437 12338 20503 12341
rect 22320 12338 22800 12368
rect 20437 12336 22800 12338
rect 20437 12280 20442 12336
rect 20498 12280 22800 12336
rect 20437 12278 22800 12280
rect 20437 12275 20503 12278
rect 22320 12248 22800 12278
rect 9489 12066 9555 12069
rect 4846 12064 9555 12066
rect 4846 12008 9494 12064
rect 9550 12008 9555 12064
rect 4846 12006 9555 12008
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 0 11794 480 11824
rect 4846 11794 4906 12006
rect 9489 12003 9555 12006
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 6821 11930 6887 11933
rect 9305 11930 9371 11933
rect 6821 11928 9371 11930
rect 6821 11872 6826 11928
rect 6882 11872 9310 11928
rect 9366 11872 9371 11928
rect 6821 11870 9371 11872
rect 6821 11867 6887 11870
rect 9305 11867 9371 11870
rect 0 11734 4906 11794
rect 5717 11794 5783 11797
rect 9397 11794 9463 11797
rect 5717 11792 9463 11794
rect 5717 11736 5722 11792
rect 5778 11736 9402 11792
rect 9458 11736 9463 11792
rect 5717 11734 9463 11736
rect 0 11704 480 11734
rect 5717 11731 5783 11734
rect 9397 11731 9463 11734
rect 17718 11732 17724 11796
rect 17788 11794 17794 11796
rect 22320 11794 22800 11824
rect 17788 11734 22800 11794
rect 17788 11732 17794 11734
rect 22320 11704 22800 11734
rect 2405 11658 2471 11661
rect 8201 11658 8267 11661
rect 8845 11658 8911 11661
rect 2405 11656 8911 11658
rect 2405 11600 2410 11656
rect 2466 11600 8206 11656
rect 8262 11600 8850 11656
rect 8906 11600 8911 11656
rect 2405 11598 8911 11600
rect 2405 11595 2471 11598
rect 8201 11595 8267 11598
rect 8845 11595 8911 11598
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 480 11326
rect 1485 11323 1551 11326
rect 18413 11386 18479 11389
rect 22320 11386 22800 11416
rect 18413 11384 22800 11386
rect 18413 11328 18418 11384
rect 18474 11328 22800 11384
rect 18413 11326 22800 11328
rect 18413 11323 18479 11326
rect 22320 11296 22800 11326
rect 12249 11250 12315 11253
rect 17769 11250 17835 11253
rect 12249 11248 17835 11250
rect 12249 11192 12254 11248
rect 12310 11192 17774 11248
rect 17830 11192 17835 11248
rect 12249 11190 17835 11192
rect 12249 11187 12315 11190
rect 17769 11187 17835 11190
rect 3417 11114 3483 11117
rect 9121 11114 9187 11117
rect 3417 11112 9187 11114
rect 3417 11056 3422 11112
rect 3478 11056 9126 11112
rect 9182 11056 9187 11112
rect 3417 11054 9187 11056
rect 3417 11051 3483 11054
rect 9121 11051 9187 11054
rect 15745 11114 15811 11117
rect 15745 11112 18568 11114
rect 15745 11056 15750 11112
rect 15806 11056 18568 11112
rect 15745 11054 18568 11056
rect 15745 11051 15811 11054
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 18508 10842 18568 11054
rect 22320 10842 22800 10872
rect 18508 10782 22800 10842
rect 0 10752 480 10782
rect 4061 10779 4127 10782
rect 22320 10752 22800 10782
rect 10961 10706 11027 10709
rect 12801 10706 12867 10709
rect 12934 10706 12940 10708
rect 10961 10704 12940 10706
rect 10961 10648 10966 10704
rect 11022 10648 12806 10704
rect 12862 10648 12940 10704
rect 10961 10646 12940 10648
rect 10961 10643 11027 10646
rect 12801 10643 12867 10646
rect 12934 10644 12940 10646
rect 13004 10644 13010 10708
rect 6085 10570 6151 10573
rect 8569 10570 8635 10573
rect 6085 10568 8635 10570
rect 6085 10512 6090 10568
rect 6146 10512 8574 10568
rect 8630 10512 8635 10568
rect 6085 10510 8635 10512
rect 6085 10507 6151 10510
rect 8569 10507 8635 10510
rect 11513 10570 11579 10573
rect 16297 10570 16363 10573
rect 11513 10568 16363 10570
rect 11513 10512 11518 10568
rect 11574 10512 16302 10568
rect 16358 10512 16363 10568
rect 11513 10510 16363 10512
rect 11513 10507 11579 10510
rect 16297 10507 16363 10510
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 14273 10434 14339 10437
rect 14406 10434 14412 10436
rect 14273 10432 14412 10434
rect 14273 10376 14278 10432
rect 14334 10376 14412 10432
rect 14273 10374 14412 10376
rect 14273 10371 14339 10374
rect 14406 10372 14412 10374
rect 14476 10372 14482 10436
rect 22320 10434 22800 10464
rect 15886 10374 22800 10434
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 4102 10236 4108 10300
rect 4172 10298 4178 10300
rect 4245 10298 4311 10301
rect 4172 10296 4311 10298
rect 4172 10240 4250 10296
rect 4306 10240 4311 10296
rect 4172 10238 4311 10240
rect 4172 10236 4178 10238
rect 4245 10235 4311 10238
rect 4245 10162 4311 10165
rect 13118 10162 13124 10164
rect 4245 10160 13124 10162
rect 4245 10104 4250 10160
rect 4306 10104 13124 10160
rect 4245 10102 13124 10104
rect 4245 10099 4311 10102
rect 13118 10100 13124 10102
rect 13188 10162 13194 10164
rect 15886 10162 15946 10374
rect 22320 10344 22800 10374
rect 13188 10102 15946 10162
rect 13188 10100 13194 10102
rect 0 10026 480 10056
rect 3969 10026 4035 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 480 9966
rect 3969 9963 4035 9966
rect 11789 10026 11855 10029
rect 15142 10026 15148 10028
rect 11789 10024 15148 10026
rect 11789 9968 11794 10024
rect 11850 9968 15148 10024
rect 11789 9966 15148 9968
rect 11789 9963 11855 9966
rect 15142 9964 15148 9966
rect 15212 10026 15218 10028
rect 18045 10026 18111 10029
rect 15212 10024 18111 10026
rect 15212 9968 18050 10024
rect 18106 9968 18111 10024
rect 15212 9966 18111 9968
rect 15212 9964 15218 9966
rect 18045 9963 18111 9966
rect 18638 9964 18644 10028
rect 18708 10026 18714 10028
rect 22320 10026 22800 10056
rect 18708 9966 22800 10026
rect 18708 9964 18714 9966
rect 22320 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 2773 9618 2839 9621
rect 1534 9616 2839 9618
rect 1534 9560 2778 9616
rect 2834 9560 2839 9616
rect 1534 9558 2839 9560
rect 0 9482 480 9512
rect 1534 9482 1594 9558
rect 2773 9555 2839 9558
rect 14733 9618 14799 9621
rect 15469 9618 15535 9621
rect 16481 9618 16547 9621
rect 14733 9616 16547 9618
rect 14733 9560 14738 9616
rect 14794 9560 15474 9616
rect 15530 9560 16486 9616
rect 16542 9560 16547 9616
rect 14733 9558 16547 9560
rect 14733 9555 14799 9558
rect 15469 9555 15535 9558
rect 16481 9555 16547 9558
rect 14917 9482 14983 9485
rect 20161 9482 20227 9485
rect 22320 9482 22800 9512
rect 0 9422 1594 9482
rect 13816 9480 15210 9482
rect 13816 9424 14922 9480
rect 14978 9424 15210 9480
rect 13816 9422 15210 9424
rect 0 9392 480 9422
rect 13816 9349 13876 9422
rect 14917 9419 14983 9422
rect 13813 9344 13879 9349
rect 13813 9288 13818 9344
rect 13874 9288 13879 9344
rect 13813 9283 13879 9288
rect 15150 9346 15210 9422
rect 20161 9480 22800 9482
rect 20161 9424 20166 9480
rect 20222 9424 22800 9480
rect 20161 9422 22800 9424
rect 20161 9419 20227 9422
rect 22320 9392 22800 9422
rect 19057 9346 19123 9349
rect 15150 9344 19123 9346
rect 15150 9288 19062 9344
rect 19118 9288 19123 9344
rect 15150 9286 19123 9288
rect 19057 9283 19123 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 4102 9148 4108 9212
rect 4172 9210 4178 9212
rect 4245 9210 4311 9213
rect 4172 9208 4311 9210
rect 4172 9152 4250 9208
rect 4306 9152 4311 9208
rect 4172 9150 4311 9152
rect 4172 9148 4178 9150
rect 4245 9147 4311 9150
rect 10041 9210 10107 9213
rect 10317 9210 10383 9213
rect 10041 9208 10383 9210
rect 10041 9152 10046 9208
rect 10102 9152 10322 9208
rect 10378 9152 10383 9208
rect 10041 9150 10383 9152
rect 10041 9147 10107 9150
rect 10317 9147 10383 9150
rect 12249 9210 12315 9213
rect 13721 9210 13787 9213
rect 12249 9208 13787 9210
rect 12249 9152 12254 9208
rect 12310 9152 13726 9208
rect 13782 9152 13787 9208
rect 12249 9150 13787 9152
rect 12249 9147 12315 9150
rect 13721 9147 13787 9150
rect 0 9074 480 9104
rect 5901 9074 5967 9077
rect 0 9072 5967 9074
rect 0 9016 5906 9072
rect 5962 9016 5967 9072
rect 0 9014 5967 9016
rect 0 8984 480 9014
rect 5901 9011 5967 9014
rect 12525 9074 12591 9077
rect 12985 9074 13051 9077
rect 17769 9074 17835 9077
rect 12525 9072 17835 9074
rect 12525 9016 12530 9072
rect 12586 9016 12990 9072
rect 13046 9016 17774 9072
rect 17830 9016 17835 9072
rect 12525 9014 17835 9016
rect 12525 9011 12591 9014
rect 12985 9011 13051 9014
rect 17769 9011 17835 9014
rect 17953 9074 18019 9077
rect 22320 9074 22800 9104
rect 17953 9072 22800 9074
rect 17953 9016 17958 9072
rect 18014 9016 22800 9072
rect 17953 9014 22800 9016
rect 17953 9011 18019 9014
rect 22320 8984 22800 9014
rect 13077 8938 13143 8941
rect 14181 8938 14247 8941
rect 13077 8936 14247 8938
rect 13077 8880 13082 8936
rect 13138 8880 14186 8936
rect 14242 8880 14247 8936
rect 13077 8878 14247 8880
rect 13077 8875 13143 8878
rect 14181 8875 14247 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 12157 8666 12223 8669
rect 12433 8666 12499 8669
rect 12157 8664 12499 8666
rect 12157 8608 12162 8664
rect 12218 8608 12438 8664
rect 12494 8608 12499 8664
rect 12157 8606 12499 8608
rect 12157 8603 12223 8606
rect 12433 8603 12499 8606
rect 0 8530 480 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 480 8470
rect 4061 8467 4127 8470
rect 18965 8530 19031 8533
rect 22320 8530 22800 8560
rect 18965 8528 22800 8530
rect 18965 8472 18970 8528
rect 19026 8472 22800 8528
rect 18965 8470 22800 8472
rect 18965 8467 19031 8470
rect 22320 8440 22800 8470
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 480 8062
rect 4061 8059 4127 8062
rect 20345 8122 20411 8125
rect 22320 8122 22800 8152
rect 20345 8120 22800 8122
rect 20345 8064 20350 8120
rect 20406 8064 22800 8120
rect 20345 8062 22800 8064
rect 20345 8059 20411 8062
rect 22320 8032 22800 8062
rect 10869 7850 10935 7853
rect 12065 7850 12131 7853
rect 10869 7848 12131 7850
rect 10869 7792 10874 7848
rect 10930 7792 12070 7848
rect 12126 7792 12131 7848
rect 10869 7790 12131 7792
rect 10869 7787 10935 7790
rect 12065 7787 12131 7790
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3785 7578 3851 7581
rect 0 7576 3851 7578
rect 0 7520 3790 7576
rect 3846 7520 3851 7576
rect 0 7518 3851 7520
rect 0 7488 480 7518
rect 3785 7515 3851 7518
rect 18597 7578 18663 7581
rect 22320 7578 22800 7608
rect 18597 7576 22800 7578
rect 18597 7520 18602 7576
rect 18658 7520 22800 7576
rect 18597 7518 22800 7520
rect 18597 7515 18663 7518
rect 22320 7488 22800 7518
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 19149 7170 19215 7173
rect 22320 7170 22800 7200
rect 19149 7168 22800 7170
rect 19149 7112 19154 7168
rect 19210 7112 22800 7168
rect 19149 7110 22800 7112
rect 19149 7107 19215 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 11605 7034 11671 7037
rect 13629 7034 13695 7037
rect 11605 7032 13695 7034
rect 11605 6976 11610 7032
rect 11666 6976 13634 7032
rect 13690 6976 13695 7032
rect 11605 6974 13695 6976
rect 11605 6971 11671 6974
rect 13629 6971 13695 6974
rect 0 6762 480 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 480 6702
rect 4061 6699 4127 6702
rect 18137 6762 18203 6765
rect 22320 6762 22800 6792
rect 18137 6760 22800 6762
rect 18137 6704 18142 6760
rect 18198 6704 22800 6760
rect 18137 6702 22800 6704
rect 18137 6699 18203 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 480 6248
rect 3969 6218 4035 6221
rect 0 6216 4035 6218
rect 0 6160 3974 6216
rect 4030 6160 4035 6216
rect 0 6158 4035 6160
rect 0 6128 480 6158
rect 3969 6155 4035 6158
rect 18137 6218 18203 6221
rect 22320 6218 22800 6248
rect 18137 6216 22800 6218
rect 18137 6160 18142 6216
rect 18198 6160 22800 6216
rect 18137 6158 22800 6160
rect 18137 6155 18203 6158
rect 22320 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 2957 5810 3023 5813
rect 0 5808 3023 5810
rect 0 5752 2962 5808
rect 3018 5752 3023 5808
rect 0 5750 3023 5752
rect 0 5720 480 5750
rect 2957 5747 3023 5750
rect 18045 5810 18111 5813
rect 22320 5810 22800 5840
rect 18045 5808 22800 5810
rect 18045 5752 18050 5808
rect 18106 5752 22800 5808
rect 18045 5750 22800 5752
rect 18045 5747 18111 5750
rect 22320 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 480 5206
rect 4061 5203 4127 5206
rect 17953 5266 18019 5269
rect 22320 5266 22800 5296
rect 17953 5264 22800 5266
rect 17953 5208 17958 5264
rect 18014 5208 22800 5264
rect 17953 5206 22800 5208
rect 17953 5203 18019 5206
rect 22320 5176 22800 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 3141 4858 3207 4861
rect 0 4856 3207 4858
rect 0 4800 3146 4856
rect 3202 4800 3207 4856
rect 0 4798 3207 4800
rect 0 4768 480 4798
rect 3141 4795 3207 4798
rect 18505 4858 18571 4861
rect 22320 4858 22800 4888
rect 18505 4856 22800 4858
rect 18505 4800 18510 4856
rect 18566 4800 22800 4856
rect 18505 4798 22800 4800
rect 18505 4795 18571 4798
rect 22320 4768 22800 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 480 4254
rect 4061 4251 4127 4254
rect 20529 4314 20595 4317
rect 22320 4314 22800 4344
rect 20529 4312 22800 4314
rect 20529 4256 20534 4312
rect 20590 4256 22800 4312
rect 20529 4254 22800 4256
rect 20529 4251 20595 4254
rect 22320 4224 22800 4254
rect 0 3906 480 3936
rect 3325 3906 3391 3909
rect 0 3904 3391 3906
rect 0 3848 3330 3904
rect 3386 3848 3391 3904
rect 0 3846 3391 3848
rect 0 3816 480 3846
rect 3325 3843 3391 3846
rect 19241 3906 19307 3909
rect 22320 3906 22800 3936
rect 19241 3904 22800 3906
rect 19241 3848 19246 3904
rect 19302 3848 22800 3904
rect 19241 3846 22800 3848
rect 19241 3843 19307 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 0 3498 480 3528
rect 3877 3498 3943 3501
rect 0 3496 3943 3498
rect 0 3440 3882 3496
rect 3938 3440 3943 3496
rect 0 3438 3943 3440
rect 0 3408 480 3438
rect 3877 3435 3943 3438
rect 17953 3498 18019 3501
rect 22320 3498 22800 3528
rect 17953 3496 22800 3498
rect 17953 3440 17958 3496
rect 18014 3440 22800 3496
rect 17953 3438 22800 3440
rect 17953 3435 18019 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 480 2984
rect 4061 2954 4127 2957
rect 0 2952 4127 2954
rect 0 2896 4066 2952
rect 4122 2896 4127 2952
rect 0 2894 4127 2896
rect 0 2864 480 2894
rect 4061 2891 4127 2894
rect 19057 2954 19123 2957
rect 22320 2954 22800 2984
rect 19057 2952 22800 2954
rect 19057 2896 19062 2952
rect 19118 2896 22800 2952
rect 19057 2894 22800 2896
rect 19057 2891 19123 2894
rect 22320 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 4245 2546 4311 2549
rect 0 2544 4311 2546
rect 0 2488 4250 2544
rect 4306 2488 4311 2544
rect 0 2486 4311 2488
rect 0 2456 480 2486
rect 4245 2483 4311 2486
rect 14181 2546 14247 2549
rect 22320 2546 22800 2576
rect 14181 2544 22800 2546
rect 14181 2488 14186 2544
rect 14242 2488 22800 2544
rect 14181 2486 22800 2488
rect 14181 2483 14247 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 2773 2002 2839 2005
rect 0 2000 2839 2002
rect 0 1944 2778 2000
rect 2834 1944 2839 2000
rect 0 1942 2839 1944
rect 0 1912 480 1942
rect 2773 1939 2839 1942
rect 18873 2002 18939 2005
rect 22320 2002 22800 2032
rect 18873 2000 22800 2002
rect 18873 1944 18878 2000
rect 18934 1944 22800 2000
rect 18873 1942 22800 1944
rect 18873 1939 18939 1942
rect 22320 1912 22800 1942
rect 0 1594 480 1624
rect 3325 1594 3391 1597
rect 0 1592 3391 1594
rect 0 1536 3330 1592
rect 3386 1536 3391 1592
rect 0 1534 3391 1536
rect 0 1504 480 1534
rect 3325 1531 3391 1534
rect 18505 1594 18571 1597
rect 22320 1594 22800 1624
rect 18505 1592 22800 1594
rect 18505 1536 18510 1592
rect 18566 1536 22800 1592
rect 18505 1534 22800 1536
rect 18505 1531 18571 1534
rect 22320 1504 22800 1534
rect 0 1050 480 1080
rect 933 1050 999 1053
rect 0 1048 999 1050
rect 0 992 938 1048
rect 994 992 999 1048
rect 0 990 999 992
rect 0 960 480 990
rect 933 987 999 990
rect 17861 1050 17927 1053
rect 22320 1050 22800 1080
rect 17861 1048 22800 1050
rect 17861 992 17866 1048
rect 17922 992 22800 1048
rect 17861 990 22800 992
rect 17861 987 17927 990
rect 22320 960 22800 990
rect 0 642 480 672
rect 3141 642 3207 645
rect 0 640 3207 642
rect 0 584 3146 640
rect 3202 584 3207 640
rect 0 582 3207 584
rect 0 552 480 582
rect 3141 579 3207 582
rect 13261 642 13327 645
rect 22320 642 22800 672
rect 13261 640 22800 642
rect 13261 584 13266 640
rect 13322 584 22800 640
rect 13261 582 22800 584
rect 13261 579 13327 582
rect 22320 552 22800 582
rect 0 234 480 264
rect 3325 234 3391 237
rect 0 232 3391 234
rect 0 176 3330 232
rect 3386 176 3391 232
rect 0 174 3391 176
rect 0 144 480 174
rect 3325 171 3391 174
rect 18781 234 18847 237
rect 22320 234 22800 264
rect 18781 232 22800 234
rect 18781 176 18786 232
rect 18842 176 22800 232
rect 18781 174 22800 176
rect 18781 171 18847 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 12940 18668 13004 18732
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 13124 17988 13188 18052
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 17724 17172 17788 17236
rect 18644 17036 18708 17100
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 15148 15540 15212 15604
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 14412 14316 14476 14380
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 14412 13228 14476 13292
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 17724 11732 17788 11796
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 12940 10644 13004 10708
rect 14412 10372 14476 10436
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4108 10236 4172 10300
rect 13124 10100 13188 10164
rect 15148 9964 15212 10028
rect 18644 9964 18708 10028
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4108 9148 4172 9212
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4107 10300 4173 10301
rect 4107 10236 4108 10300
rect 4172 10236 4173 10300
rect 4107 10235 4173 10236
rect 4110 9213 4170 10235
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4107 9212 4173 9213
rect 4107 9148 4108 9212
rect 4172 9148 4173 9212
rect 4107 9147 4173 9148
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 12939 18732 13005 18733
rect 12939 18668 12940 18732
rect 13004 18668 13005 18732
rect 12939 18667 13005 18668
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 12942 10709 13002 18667
rect 13123 18052 13189 18053
rect 13123 17988 13124 18052
rect 13188 17988 13189 18052
rect 13123 17987 13189 17988
rect 12939 10708 13005 10709
rect 12939 10644 12940 10708
rect 13004 10644 13005 10708
rect 12939 10643 13005 10644
rect 13126 10165 13186 17987
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 17723 17236 17789 17237
rect 17723 17172 17724 17236
rect 17788 17172 17789 17236
rect 17723 17171 17789 17172
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 15147 15604 15213 15605
rect 15147 15540 15148 15604
rect 15212 15540 15213 15604
rect 15147 15539 15213 15540
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14411 14380 14477 14381
rect 14411 14316 14412 14380
rect 14476 14316 14477 14380
rect 14411 14315 14477 14316
rect 14414 13293 14474 14315
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14411 13292 14477 13293
rect 14411 13228 14412 13292
rect 14476 13228 14477 13292
rect 14411 13227 14477 13228
rect 14414 10437 14474 13227
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14411 10436 14477 10437
rect 14411 10372 14412 10436
rect 14476 10372 14477 10436
rect 14411 10371 14477 10372
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 13123 10164 13189 10165
rect 13123 10100 13124 10164
rect 13188 10100 13189 10164
rect 13123 10099 13189 10100
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 9280 14992 10304
rect 15150 10029 15210 15539
rect 17726 11797 17786 17171
rect 18104 16352 18424 17376
rect 18643 17100 18709 17101
rect 18643 17036 18644 17100
rect 18708 17036 18709 17100
rect 18643 17035 18709 17036
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 17723 11796 17789 11797
rect 17723 11732 17724 11796
rect 17788 11732 17789 11796
rect 17723 11731 17789 11732
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 15147 10028 15213 10029
rect 15147 9964 15148 10028
rect 15212 9964 15213 10028
rect 15147 9963 15213 9964
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 9824 18424 10848
rect 18646 10029 18706 17035
rect 18643 10028 18709 10029
rect 18643 9964 18644 10028
rect 18708 9964 18709 10028
rect 18643 9963 18709 9964
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1605641404
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1605641404
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1605641404
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1605641404
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1605641404
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1605641404
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1605641404
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1605641404
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1605641404
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1605641404
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1605641404
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1605641404
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1605641404
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1605641404
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1605641404
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1605641404
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1605641404
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10672 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_101
timestamp 1605641404
transform 1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_120
timestamp 1605641404
transform 1 0 12144 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_132
timestamp 1605641404
transform 1 0 13248 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1605641404
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1605641404
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1605641404
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1605641404
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1605641404
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1605641404
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1605641404
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1605641404
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1605641404
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1605641404
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1605641404
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1605641404
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1605641404
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1605641404
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1605641404
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1605641404
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1605641404
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1605641404
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1605641404
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1605641404
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1605641404
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1605641404
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1605641404
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1605641404
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1605641404
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1605641404
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1605641404
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1605641404
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1605641404
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1605641404
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _029_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_110
timestamp 1605641404
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1605641404
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_126
timestamp 1605641404
transform 1 0 12696 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_138
timestamp 1605641404
transform 1 0 13800 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_150
timestamp 1605641404
transform 1 0 14904 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_162
timestamp 1605641404
transform 1 0 16008 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_174
timestamp 1605641404
transform 1 0 17112 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1605641404
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1605641404
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1605641404
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1605641404
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1605641404
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1605641404
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1605641404
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1605641404
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1605641404
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10304 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_93
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_99
timestamp 1605641404
transform 1 0 10212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1605641404
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_98
timestamp 1605641404
transform 1 0 10120 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11316 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10948 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1605641404
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_106
timestamp 1605641404
transform 1 0 10856 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_116
timestamp 1605641404
transform 1 0 11776 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1605641404
transform 1 0 14352 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1605641404
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1605641404
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_132
timestamp 1605641404
transform 1 0 13248 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14812 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1605641404
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp 1605641404
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 1605641404
transform 1 0 15640 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_166
timestamp 1605641404
transform 1 0 16376 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16468 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1605641404
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_176
timestamp 1605641404
transform 1 0 17296 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1605641404
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1605641404
transform 1 0 20056 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1605641404
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1605641404
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1605641404
transform 1 0 19136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1605641404
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1605641404
transform 1 0 20884 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1605641404
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1605641404
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1605641404
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1605641404
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1605641404
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_105
timestamp 1605641404
transform 1 0 10764 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_118
timestamp 1605641404
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_140
timestamp 1605641404
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1605641404
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1605641404
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 17664 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_174
timestamp 1605641404
transform 1 0 17112 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_189
timestamp 1605641404
transform 1 0 18492 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1605641404
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1605641404
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 3956 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1605641404
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1605641404
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1605641404
transform 1 0 4968 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_45
timestamp 1605641404
transform 1 0 5244 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1605641404
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1605641404
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10304 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1605641404
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_98
timestamp 1605641404
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1605641404
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14076 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1605641404
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16192 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_157
timestamp 1605641404
transform 1 0 15548 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_163
timestamp 1605641404
transform 1 0 16100 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1605641404
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_173
timestamp 1605641404
transform 1 0 17020 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_177
timestamp 1605641404
transform 1 0 17388 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1605641404
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19044 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1605641404
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_211
timestamp 1605641404
transform 1 0 20516 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1605641404
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2576 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_15
timestamp 1605641404
transform 1 0 2484 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4140 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1605641404
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5796 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_49
timestamp 1605641404
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_60
timestamp 1605641404
transform 1 0 6624 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_72
timestamp 1605641404
transform 1 0 7728 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9844 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1605641404
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1605641404
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10856 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12512 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1605641404
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14076 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_133
timestamp 1605641404
transform 1 0 13340 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16008 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1605641404
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 17664 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1605641404
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18952 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_189
timestamp 1605641404
transform 1 0 18492 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_193
timestamp 1605641404
transform 1 0 18860 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1605641404
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1605641404
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1656 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_22
timestamp 1605641404
transform 1 0 3128 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1605641404
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1605641404
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1605641404
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1605641404
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1605641404
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10580 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 9568 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_86
timestamp 1605641404
transform 1 0 9016 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1605641404
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_112
timestamp 1605641404
transform 1 0 11408 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1605641404
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_123
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12972 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_145
timestamp 1605641404
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14628 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_163
timestamp 1605641404
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1605641404
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1605641404
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_184
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18768 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_208
timestamp 1605641404
transform 1 0 20240 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _093_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 20516 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1605641404
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1605641404
transform 1 0 21252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2208 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1472 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1605641404
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1605641404
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1605641404
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1605641404
transform 1 0 6808 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5520 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1605641404
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1605641404
transform 1 0 6348 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 1605641404
transform 1 0 6716 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7268 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1605641404
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1605641404
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1605641404
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12236 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11960 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_109
timestamp 1605641404
transform 1 0 11132 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_117
timestamp 1605641404
transform 1 0 11868 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1605641404
transform 1 0 13248 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14260 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_130
timestamp 1605641404
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1605641404
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 16100 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1605641404
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_162
timestamp 1605641404
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 17848 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_179
timestamp 1605641404
transform 1 0 17572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18860 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20056 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_191
timestamp 1605641404
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1605641404
transform 1 0 19688 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1605641404
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1605641404
transform 1 0 1656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1605641404
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_10
timestamp 1605641404
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1605641404
transform 1 0 2208 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1605641404
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1605641404
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_27
timestamp 1605641404
transform 1 0 3588 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_21
timestamp 1605641404
transform 1 0 3036 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1605641404
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1605641404
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4692 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4508 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_55
timestamp 1605641404
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_53
timestamp 1605641404
transform 1 0 5980 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1605641404
transform 1 0 6716 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7820 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1605641404
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_82
timestamp 1605641404
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1605641404
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1605641404
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 8832 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1605641404
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1605641404
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1605641404
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1605641404
transform 1 0 11500 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1605641404
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1605641404
transform 1 0 11132 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1605641404
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1605641404
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1605641404
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 13984 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1605641404
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1605641404
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 1605641404
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1605641404
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16376 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15456 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 16192 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_154
timestamp 1605641404
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1605641404
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1605641404
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1605641404
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18216 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_167
timestamp 1605641404
transform 1 0 16468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_171
timestamp 1605641404
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1605641404
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_182
timestamp 1605641404
transform 1 0 17848 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 19964 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 19412 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_202
timestamp 1605641404
transform 1 0 19688 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1605641404
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_208
timestamp 1605641404
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_214
timestamp 1605641404
transform 1 0 20792 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_218
timestamp 1605641404
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1605641404
transform 1 0 1656 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2116 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1605641404
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 3864 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 1605641404
transform 1 0 3588 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_39
timestamp 1605641404
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 4968 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_45
timestamp 1605641404
transform 1 0 5244 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_49
timestamp 1605641404
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6900 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8004 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_72
timestamp 1605641404
transform 1 0 7728 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8832 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1605641404
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13800 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 13524 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_132
timestamp 1605641404
transform 1 0 13248 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14812 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_147
timestamp 1605641404
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_165
timestamp 1605641404
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1605641404
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1605641404
transform 1 0 18124 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16468 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_176
timestamp 1605641404
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1605641404
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 18492 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1605641404
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_205
timestamp 1605641404
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 20332 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1605641404
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1605641404
transform 1 0 2944 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1605641404
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1605641404
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6624 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 6348 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1605641404
transform 1 0 5520 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_56
timestamp 1605641404
transform 1 0 6256 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8280 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_76
timestamp 1605641404
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10488 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1605641404
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1605641404
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1605641404
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12328 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_138
timestamp 1605641404
transform 1 0 13800 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16284 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1605641404
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1605641404
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1605641404
transform 1 0 17296 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1605641404
transform 1 0 18308 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1605641404
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1605641404
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 19688 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_196
timestamp 1605641404
transform 1 0 19136 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1605641404
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1605641404
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_16
timestamp 1605641404
transform 1 0 2576 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4324 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 3312 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_33
timestamp 1605641404
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1605641404
transform 1 0 5980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1605641404
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1605641404
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1605641404
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1605641404
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1605641404
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9936 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8832 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_93
timestamp 1605641404
transform 1 0 9660 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_112
timestamp 1605641404
transform 1 0 11408 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_118
timestamp 1605641404
transform 1 0 11960 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1605641404
transform 1 0 13432 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1605641404
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1605641404
transform 1 0 13708 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1605641404
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14628 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16284 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1605641404
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1605641404
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_174
timestamp 1605641404
transform 1 0 17112 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1605641404
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 19136 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_193
timestamp 1605641404
transform 1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1605641404
transform 1 0 20792 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1605641404
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1605641404
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1564 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_21
timestamp 1605641404
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1605641404
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_41
timestamp 1605641404
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6164 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 5152 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1605641404
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_71
timestamp 1605641404
transform 1 0 7636 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 9016 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1605641404
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1605641404
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_102
timestamp 1605641404
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 11224 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13892 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12880 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1605641404
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1605641404
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15732 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1605641404
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1605641404
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1605641404
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17388 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1605641404
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1605641404
transform 1 0 19044 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 19504 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_193
timestamp 1605641404
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1605641404
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1605641404
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1605641404
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1748 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2852 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1605641404
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1605641404
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1605641404
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1605641404
transform 1 0 3864 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_28
timestamp 1605641404
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1605641404
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1605641404
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1605641404
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6164 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 5060 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1605641404
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_52
timestamp 1605641404
transform 1 0 5888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8648 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7268 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1605641404
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_76
timestamp 1605641404
transform 1 0 8096 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_64
timestamp 1605641404
transform 1 0 6992 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10212 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1605641404
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1605641404
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11316 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1605641404
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1605641404
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_108
timestamp 1605641404
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_119
timestamp 1605641404
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1605641404
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13432 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_19_132
timestamp 1605641404
transform 1 0 13248 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1605641404
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_131
timestamp 1605641404
transform 1 0 13156 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_143
timestamp 1605641404
transform 1 0 14260 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1605641404
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1605641404
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14996 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1605641404
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_160
timestamp 1605641404
transform 1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_164
timestamp 1605641404
transform 1 0 16192 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_160
timestamp 1605641404
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16100 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 16284 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17112 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1605641404
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_172
timestamp 1605641404
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19320 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18768 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 19780 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1605641404
transform 1 0 18860 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_197
timestamp 1605641404
transform 1 0 19228 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1605641404
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_201
timestamp 1605641404
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_214
timestamp 1605641404
transform 1 0 20792 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1605641404
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1605641404
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1605641404
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp 1605641404
transform 1 0 3772 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1605641404
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_42
timestamp 1605641404
transform 1 0 4968 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1605641404
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8556 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 8280 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1605641404
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_76
timestamp 1605641404
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10212 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1605641404
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1605641404
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1605641404
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1605641404
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13708 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 13432 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1605641404
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 14720 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 15732 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1605641404
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1605641404
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18216 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17020 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1605641404
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1605641404
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18952 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19964 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_192
timestamp 1605641404
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_203
timestamp 1605641404
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_214
timestamp 1605641404
transform 1 0 20792 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1656 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_12
timestamp 1605641404
transform 1 0 2208 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5888 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_48
timestamp 1605641404
transform 1 0 5520 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1605641404
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_80
timestamp 1605641404
transform 1 0 8464 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9844 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1605641404
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_104
timestamp 1605641404
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10856 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12604 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_122
timestamp 1605641404
transform 1 0 12328 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1605641404
transform 1 0 14076 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1605641404
transform 1 0 14628 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 15364 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1605641404
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17848 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17020 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1605641404
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_179
timestamp 1605641404
transform 1 0 17572 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19596 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_198
timestamp 1605641404
transform 1 0 19320 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1605641404
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1605641404
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1605641404
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 2392 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_11
timestamp 1605641404
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1605641404
transform 1 0 4416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 3404 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1605641404
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1605641404
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_39
timestamp 1605641404
transform 1 0 4692 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5244 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1605641404
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7820 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1605641404
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_82
timestamp 1605641404
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9936 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_23_93
timestamp 1605641404
transform 1 0 9660 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1605641404
transform 1 0 12604 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1605641404
transform 1 0 10764 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1605641404
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 13156 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1605641404
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15824 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 14812 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_147
timestamp 1605641404
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1605641404
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1605641404
transform 1 0 17480 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1605641404
transform 1 0 18308 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_176
timestamp 1605641404
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1605641404
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18860 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1605641404
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20516 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1605641404
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1605641404
transform 1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1605641404
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2300 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1605641404
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1605641404
transform 1 0 3312 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4324 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1605641404
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1605641404
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6164 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_51
timestamp 1605641404
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7820 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1605641404
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1605641404
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10120 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 8832 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_87
timestamp 1605641404
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1605641404
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1605641404
transform 1 0 10028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1605641404
transform 1 0 11776 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_114
timestamp 1605641404
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1605641404
transform 1 0 12604 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13248 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 12972 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15456 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1605641404
transform 1 0 14720 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1605641404
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_165
timestamp 1605641404
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16468 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1605641404
transform 1 0 17296 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19964 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18952 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_189
timestamp 1605641404
transform 1 0 18492 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_193
timestamp 1605641404
transform 1 0 18860 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1605641404
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1605641404
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_218
timestamp 1605641404
transform 1 0 21160 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2484 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1748 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1605641404
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4140 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_31
timestamp 1605641404
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1605641404
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_53
timestamp 1605641404
transform 1 0 5980 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8372 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6992 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_73
timestamp 1605641404
transform 1 0 7820 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10028 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1605641404
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1605641404
transform 1 0 11868 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1605641404
transform 1 0 11500 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1605641404
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13432 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14444 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1605641404
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1605641404
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1605641404
transform 1 0 15640 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16192 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1605641404
transform 1 0 15272 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1605641404
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1605641404
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1605641404
transform 1 0 18216 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_173
timestamp 1605641404
transform 1 0 17020 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1605641404
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18768 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1605641404
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_208
timestamp 1605641404
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20424 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_216
timestamp 1605641404
transform 1 0 20976 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1605641404
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1605641404
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_17
timestamp 1605641404
transform 1 0 2668 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1605641404
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1605641404
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1932 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2944 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4600 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1605641404
transform 1 0 4416 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1605641404
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1605641404
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5428 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1605641404
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1605641404
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_47
timestamp 1605641404
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1605641404
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8280 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_67
timestamp 1605641404
transform 1 0 7268 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_75
timestamp 1605641404
transform 1 0 8004 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_78
timestamp 1605641404
transform 1 0 8280 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_86
timestamp 1605641404
transform 1 0 9016 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1605641404
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1605641404
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9292 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1605641404
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_101
timestamp 1605641404
transform 1 0 10396 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10488 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11500 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1605641404
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_122
timestamp 1605641404
transform 1 0 12328 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1605641404
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1605641404
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1605641404
transform 1 0 12788 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1605641404
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13248 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13984 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_26_126
timestamp 1605641404
transform 1 0 12696 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_130
timestamp 1605641404
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1605641404
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1605641404
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 1605641404
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1605641404
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1605641404
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14996 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1605641404
transform 1 0 15456 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_157
timestamp 1605641404
transform 1 0 15548 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1605641404
transform 1 0 15824 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15824 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16008 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1605641404
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1605641404
transform 1 0 18032 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18216 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_178
timestamp 1605641404
transform 1 0 17480 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_176
timestamp 1605641404
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1605641404
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1605641404
transform 1 0 20056 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19596 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18584 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1605641404
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1605641404
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1605641404
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_202
timestamp 1605641404
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1605641404
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_218
timestamp 1605641404
transform 1 0 21160 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1605641404
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1605641404
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1605641404
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1605641404
transform 1 0 1564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1605641404
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1605641404
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4324 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1605641404
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5336 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_44
timestamp 1605641404
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_62
timestamp 1605641404
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6992 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_73
timestamp 1605641404
transform 1 0 7820 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10212 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1605641404
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_93
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1605641404
transform 1 0 11868 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_115
timestamp 1605641404
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_120
timestamp 1605641404
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_139
timestamp 1605641404
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16284 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1605641404
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1605641404
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1605641404
transform 1 0 17388 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17940 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_28_171
timestamp 1605641404
transform 1 0 16836 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_181
timestamp 1605641404
transform 1 0 17756 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19964 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_199
timestamp 1605641404
transform 1 0 19412 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1605641404
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1605641404
transform 1 0 1564 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1605641404
transform 1 0 2852 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1605641404
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1605641404
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1605641404
transform 1 0 3404 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4232 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1605641404
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_29
timestamp 1605641404
transform 1 0 3772 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_33
timestamp 1605641404
transform 1 0 4140 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_50
timestamp 1605641404
transform 1 0 5704 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1605641404
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8004 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1605641404
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1605641404
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1605641404
transform 1 0 11316 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12512 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_109
timestamp 1605641404
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1605641404
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13524 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_133
timestamp 1605641404
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1605641404
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1605641404
transform 1 0 16284 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14536 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_162
timestamp 1605641404
transform 1 0 16008 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1605641404
transform 1 0 16836 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1605641404
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1605641404
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1605641404
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1605641404
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1605641404
transform 1 0 19412 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19964 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_193
timestamp 1605641404
transform 1 0 18860 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1605641404
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1605641404
transform 1 0 20700 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_211
timestamp 1605641404
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_217
timestamp 1605641404
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1605641404
transform 1 0 2300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1605641404
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2944 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1605641404
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_17
timestamp 1605641404
transform 1 0 2668 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1605641404
transform 1 0 4784 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_26
timestamp 1605641404
transform 1 0 3496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1605641404
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_32
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5888 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_43
timestamp 1605641404
transform 1 0 5060 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_51
timestamp 1605641404
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_61
timestamp 1605641404
transform 1 0 6716 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7912 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_73
timestamp 1605641404
transform 1 0 7820 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_83
timestamp 1605641404
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9936 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1605641404
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1605641404
transform 1 0 11040 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1605641404
transform 1 0 11500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12052 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_105
timestamp 1605641404
transform 1 0 10764 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_111
timestamp 1605641404
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_117
timestamp 1605641404
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1605641404
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14168 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1605641404
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_140
timestamp 1605641404
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15916 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1605641404
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_158
timestamp 1605641404
transform 1 0 15640 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17572 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1605641404
transform 1 0 17388 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1605641404
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19228 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_195
timestamp 1605641404
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1605641404
transform 1 0 19780 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_207
timestamp 1605641404
transform 1 0 20148 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1605641404
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_218
timestamp 1605641404
transform 1 0 21160 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1605641404
transform 1 0 2576 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1605641404
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_11
timestamp 1605641404
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 1605641404
transform 1 0 2484 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_20
timestamp 1605641404
transform 1 0 2944 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1605641404
transform 1 0 4600 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1605641404
transform 1 0 3496 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1605641404
transform 1 0 4048 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_30
timestamp 1605641404
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1605641404
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_42
timestamp 1605641404
transform 1 0 4968 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_54
timestamp 1605641404
transform 1 0 6072 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1605641404
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1605641404
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10488 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1605641404
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1605641404
transform 1 0 10120 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11408 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1605641404
transform 1 0 11040 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1605641404
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13156 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_129
timestamp 1605641404
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15088 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16100 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1605641404
transform 1 0 14628 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_151
timestamp 1605641404
transform 1 0 14996 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_161
timestamp 1605641404
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1605641404
transform 1 0 16652 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1605641404
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1605641404
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19044 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1605641404
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1605641404
transform 1 0 19596 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1605641404
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1605641404
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1605641404
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1605641404
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1605641404
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1605641404
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1605641404
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1605641404
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_17
timestamp 1605641404
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1605641404
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1605641404
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1605641404
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1605641404
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1605641404
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1605641404
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1605641404
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1605641404
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1605641404
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1605641404
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1605641404
transform 1 0 13892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12696 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1605641404
transform 1 0 13524 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_143
timestamp 1605641404
transform 1 0 14260 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1605641404
transform 1 0 16192 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1605641404
transform 1 0 15640 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1605641404
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1605641404
transform 1 0 15180 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_156
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_162
timestamp 1605641404
transform 1 0 16008 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1605641404
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1605641404
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1605641404
transform 1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1605641404
transform 1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1605641404
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1605641404
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1605641404
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_193
timestamp 1605641404
transform 1 0 18860 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1605641404
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1605641404
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1605641404
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1605641404
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 11334 0 11390 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 18970 0 19026 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 22320 22448 22800 22568 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 3974 22320 4030 22800 6 chany_top_in[0]
port 82 nsew default input
rlabel metal2 s 8758 22320 8814 22800 6 chany_top_in[10]
port 83 nsew default input
rlabel metal2 s 9218 22320 9274 22800 6 chany_top_in[11]
port 84 nsew default input
rlabel metal2 s 9678 22320 9734 22800 6 chany_top_in[12]
port 85 nsew default input
rlabel metal2 s 10138 22320 10194 22800 6 chany_top_in[13]
port 86 nsew default input
rlabel metal2 s 10598 22320 10654 22800 6 chany_top_in[14]
port 87 nsew default input
rlabel metal2 s 11058 22320 11114 22800 6 chany_top_in[15]
port 88 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[16]
port 89 nsew default input
rlabel metal2 s 12070 22320 12126 22800 6 chany_top_in[17]
port 90 nsew default input
rlabel metal2 s 12530 22320 12586 22800 6 chany_top_in[18]
port 91 nsew default input
rlabel metal2 s 12990 22320 13046 22800 6 chany_top_in[19]
port 92 nsew default input
rlabel metal2 s 4434 22320 4490 22800 6 chany_top_in[1]
port 93 nsew default input
rlabel metal2 s 4894 22320 4950 22800 6 chany_top_in[2]
port 94 nsew default input
rlabel metal2 s 5354 22320 5410 22800 6 chany_top_in[3]
port 95 nsew default input
rlabel metal2 s 5906 22320 5962 22800 6 chany_top_in[4]
port 96 nsew default input
rlabel metal2 s 6366 22320 6422 22800 6 chany_top_in[5]
port 97 nsew default input
rlabel metal2 s 6826 22320 6882 22800 6 chany_top_in[6]
port 98 nsew default input
rlabel metal2 s 7286 22320 7342 22800 6 chany_top_in[7]
port 99 nsew default input
rlabel metal2 s 7746 22320 7802 22800 6 chany_top_in[8]
port 100 nsew default input
rlabel metal2 s 8206 22320 8262 22800 6 chany_top_in[9]
port 101 nsew default input
rlabel metal2 s 13450 22320 13506 22800 6 chany_top_out[0]
port 102 nsew default tristate
rlabel metal2 s 18234 22320 18290 22800 6 chany_top_out[10]
port 103 nsew default tristate
rlabel metal2 s 18694 22320 18750 22800 6 chany_top_out[11]
port 104 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 chany_top_out[12]
port 105 nsew default tristate
rlabel metal2 s 19614 22320 19670 22800 6 chany_top_out[13]
port 106 nsew default tristate
rlabel metal2 s 20166 22320 20222 22800 6 chany_top_out[14]
port 107 nsew default tristate
rlabel metal2 s 20626 22320 20682 22800 6 chany_top_out[15]
port 108 nsew default tristate
rlabel metal2 s 21086 22320 21142 22800 6 chany_top_out[16]
port 109 nsew default tristate
rlabel metal2 s 21546 22320 21602 22800 6 chany_top_out[17]
port 110 nsew default tristate
rlabel metal2 s 22006 22320 22062 22800 6 chany_top_out[18]
port 111 nsew default tristate
rlabel metal2 s 22466 22320 22522 22800 6 chany_top_out[19]
port 112 nsew default tristate
rlabel metal2 s 13910 22320 13966 22800 6 chany_top_out[1]
port 113 nsew default tristate
rlabel metal2 s 14462 22320 14518 22800 6 chany_top_out[2]
port 114 nsew default tristate
rlabel metal2 s 14922 22320 14978 22800 6 chany_top_out[3]
port 115 nsew default tristate
rlabel metal2 s 15382 22320 15438 22800 6 chany_top_out[4]
port 116 nsew default tristate
rlabel metal2 s 15842 22320 15898 22800 6 chany_top_out[5]
port 117 nsew default tristate
rlabel metal2 s 16302 22320 16358 22800 6 chany_top_out[6]
port 118 nsew default tristate
rlabel metal2 s 16762 22320 16818 22800 6 chany_top_out[7]
port 119 nsew default tristate
rlabel metal2 s 17314 22320 17370 22800 6 chany_top_out[8]
port 120 nsew default tristate
rlabel metal2 s 17774 22320 17830 22800 6 chany_top_out[9]
port 121 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_11_
port 122 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_13_
port 123 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_15_
port 124 nsew default input
rlabel metal3 s 0 3816 480 3936 6 left_bottom_grid_pin_17_
port 125 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 126 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 127 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_5_
port 128 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_7_
port 129 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_9_
port 130 nsew default input
rlabel metal2 s 3790 0 3846 480 6 prog_clk
port 131 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_11_
port 132 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_13_
port 133 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_15_
port 134 nsew default input
rlabel metal3 s 22320 3816 22800 3936 6 right_bottom_grid_pin_17_
port 135 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_1_
port 136 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_3_
port 137 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_5_
port 138 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_7_
port 139 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_9_
port 140 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 141 nsew default input
rlabel metal2 s 662 22320 718 22800 6 top_left_grid_pin_43_
port 142 nsew default input
rlabel metal2 s 1122 22320 1178 22800 6 top_left_grid_pin_44_
port 143 nsew default input
rlabel metal2 s 1582 22320 1638 22800 6 top_left_grid_pin_45_
port 144 nsew default input
rlabel metal2 s 2042 22320 2098 22800 6 top_left_grid_pin_46_
port 145 nsew default input
rlabel metal2 s 2502 22320 2558 22800 6 top_left_grid_pin_47_
port 146 nsew default input
rlabel metal2 s 3054 22320 3110 22800 6 top_left_grid_pin_48_
port 147 nsew default input
rlabel metal2 s 3514 22320 3570 22800 6 top_left_grid_pin_49_
port 148 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 149 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
