VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__3_
  CLASS BLOCK ;
  FOREIGN sb_1__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 137.320 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.400 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 53.760 140.000 54.360 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 58.520 140.000 59.120 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 63.960 140.000 64.560 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.160 140.000 74.760 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 79.600 140.000 80.200 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 85.040 140.000 85.640 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.800 140.000 90.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.240 140.000 95.840 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 12.280 140.000 12.880 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.040 140.000 17.640 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 22.480 140.000 23.080 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 27.920 140.000 28.520 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 32.680 140.000 33.280 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 43.560 140.000 44.160 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 48.320 140.000 48.920 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 2.400 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END left_top_grid_pin_11_
  PIN left_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 2.400 131.880 ;
    END
  END left_top_grid_pin_13_
  PIN left_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 2.400 137.320 ;
    END
  END left_top_grid_pin_15_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END left_top_grid_pin_1_
  PIN left_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END left_top_grid_pin_3_
  PIN left_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END left_top_grid_pin_5_
  PIN left_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END left_top_grid_pin_7_
  PIN left_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END left_top_grid_pin_9_
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.080 140.000 2.680 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END right_top_grid_pin_11_
  PIN right_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 131.280 140.000 131.880 ;
    END
  END right_top_grid_pin_13_
  PIN right_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.720 140.000 137.320 ;
    END
  END right_top_grid_pin_15_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 100.000 140.000 100.600 ;
    END
  END right_top_grid_pin_1_
  PIN right_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 105.440 140.000 106.040 ;
    END
  END right_top_grid_pin_3_
  PIN right_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 110.880 140.000 111.480 ;
    END
  END right_top_grid_pin_5_
  PIN right_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.640 140.000 116.240 ;
    END
  END right_top_grid_pin_7_
  PIN right_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.080 140.000 121.680 ;
    END
  END right_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 2.830 2.760 134.320 128.080 ;
      LAYER met2 ;
        RECT 1.930 2.680 137.450 137.205 ;
        RECT 1.930 2.195 2.110 2.680 ;
        RECT 2.950 2.195 6.710 2.680 ;
        RECT 7.550 2.195 11.310 2.680 ;
        RECT 12.150 2.195 16.370 2.680 ;
        RECT 17.210 2.195 20.970 2.680 ;
        RECT 21.810 2.195 26.030 2.680 ;
        RECT 26.870 2.195 30.630 2.680 ;
        RECT 31.470 2.195 35.690 2.680 ;
        RECT 36.530 2.195 40.290 2.680 ;
        RECT 41.130 2.195 45.350 2.680 ;
        RECT 46.190 2.195 49.950 2.680 ;
        RECT 50.790 2.195 55.010 2.680 ;
        RECT 55.850 2.195 59.610 2.680 ;
        RECT 60.450 2.195 64.670 2.680 ;
        RECT 65.510 2.195 69.270 2.680 ;
        RECT 70.110 2.195 74.330 2.680 ;
        RECT 75.170 2.195 78.930 2.680 ;
        RECT 79.770 2.195 83.990 2.680 ;
        RECT 84.830 2.195 88.590 2.680 ;
        RECT 89.430 2.195 93.650 2.680 ;
        RECT 94.490 2.195 98.250 2.680 ;
        RECT 99.090 2.195 103.310 2.680 ;
        RECT 104.150 2.195 107.910 2.680 ;
        RECT 108.750 2.195 112.970 2.680 ;
        RECT 113.810 2.195 117.570 2.680 ;
        RECT 118.410 2.195 122.630 2.680 ;
        RECT 123.470 2.195 127.230 2.680 ;
        RECT 128.070 2.195 132.290 2.680 ;
        RECT 133.130 2.195 136.890 2.680 ;
      LAYER met3 ;
        RECT 2.800 136.320 137.200 137.185 ;
        RECT 1.905 132.280 137.600 136.320 ;
        RECT 2.800 130.880 137.200 132.280 ;
        RECT 1.905 127.520 137.600 130.880 ;
        RECT 2.800 126.120 137.200 127.520 ;
        RECT 1.905 122.080 137.600 126.120 ;
        RECT 2.800 120.680 137.200 122.080 ;
        RECT 1.905 116.640 137.600 120.680 ;
        RECT 2.800 115.240 137.200 116.640 ;
        RECT 1.905 111.880 137.600 115.240 ;
        RECT 2.800 110.480 137.200 111.880 ;
        RECT 1.905 106.440 137.600 110.480 ;
        RECT 2.800 105.040 137.200 106.440 ;
        RECT 1.905 101.000 137.600 105.040 ;
        RECT 2.800 99.600 137.200 101.000 ;
        RECT 1.905 96.240 137.600 99.600 ;
        RECT 2.800 94.840 137.200 96.240 ;
        RECT 1.905 90.800 137.600 94.840 ;
        RECT 2.800 89.400 137.200 90.800 ;
        RECT 1.905 86.040 137.600 89.400 ;
        RECT 2.800 84.640 137.200 86.040 ;
        RECT 1.905 80.600 137.600 84.640 ;
        RECT 2.800 79.200 137.200 80.600 ;
        RECT 1.905 75.160 137.600 79.200 ;
        RECT 2.800 73.760 137.200 75.160 ;
        RECT 1.905 70.400 137.600 73.760 ;
        RECT 2.800 69.000 137.200 70.400 ;
        RECT 1.905 64.960 137.600 69.000 ;
        RECT 2.800 63.560 137.200 64.960 ;
        RECT 1.905 59.520 137.600 63.560 ;
        RECT 2.800 58.120 137.200 59.520 ;
        RECT 1.905 54.760 137.600 58.120 ;
        RECT 2.800 53.360 137.200 54.760 ;
        RECT 1.905 49.320 137.600 53.360 ;
        RECT 2.800 47.920 137.200 49.320 ;
        RECT 1.905 44.560 137.600 47.920 ;
        RECT 2.800 43.160 137.200 44.560 ;
        RECT 1.905 39.120 137.600 43.160 ;
        RECT 2.800 37.720 137.200 39.120 ;
        RECT 1.905 33.680 137.600 37.720 ;
        RECT 2.800 32.280 137.200 33.680 ;
        RECT 1.905 28.920 137.600 32.280 ;
        RECT 2.800 27.520 137.200 28.920 ;
        RECT 1.905 23.480 137.600 27.520 ;
        RECT 2.800 22.080 137.200 23.480 ;
        RECT 1.905 18.040 137.600 22.080 ;
        RECT 2.800 16.640 137.200 18.040 ;
        RECT 1.905 13.280 137.600 16.640 ;
        RECT 2.800 11.880 137.200 13.280 ;
        RECT 1.905 7.840 137.600 11.880 ;
        RECT 2.800 6.440 137.200 7.840 ;
        RECT 1.905 3.080 137.600 6.440 ;
        RECT 2.800 2.215 137.200 3.080 ;
      LAYER met4 ;
        RECT 22.375 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_1__3_
END LIBRARY

