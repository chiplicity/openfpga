magic
tech sky130A
magscale 1 2
timestamp 1608763374
<< checkpaint >>
rect -1260 -1260 24060 23828
<< locali >>
rect 4537 19703 4571 19941
rect 3433 18751 3467 18921
rect 5181 18683 5215 18785
rect 2881 17119 2915 17289
rect 13001 14263 13035 14365
rect 4537 12699 4571 12869
rect 9505 12631 9539 12869
rect 3801 12087 3835 12325
rect 4997 12155 5031 12257
rect 8585 11611 8619 11849
rect 9965 11679 9999 11781
rect 9873 11543 9907 11645
rect 8401 10591 8435 10761
rect 8493 10455 8527 10557
rect 14013 9911 14047 10217
rect 14749 9911 14783 10217
rect 13277 9367 13311 9469
rect 9137 8959 9171 9061
rect 9505 8891 9539 9129
rect 5457 8279 5491 8381
rect 11897 8347 11931 8585
rect 15393 8415 15427 8585
rect 5365 7735 5399 7905
rect 12909 7735 12943 7837
rect 12851 7701 12943 7735
rect 3893 7191 3927 7361
rect 18521 7327 18555 7497
rect 2881 6783 2915 6953
rect 2973 6715 3007 6953
rect 8493 6715 8527 6953
rect 9413 6715 9447 6953
rect 12817 6647 12851 6749
rect 15853 6647 15887 6817
rect 10241 6103 10275 6205
rect 18797 6103 18831 6205
rect 9505 5627 9539 5865
rect 11621 5695 11655 5797
rect 7941 5015 7975 5321
rect 8861 5015 8895 5117
rect 18245 4471 18279 4641
rect 18337 4471 18371 4709
rect 18981 4607 19015 4777
rect 21741 4199 21775 4981
rect 8677 3927 8711 4097
rect 15853 3587 15887 3689
rect 11897 3383 11931 3553
rect 16313 2975 16347 3145
rect 3801 2839 3835 2941
rect 20913 2839 20947 2941
rect 16405 2499 16439 2601
<< viali >>
rect 1961 20009 1995 20043
rect 3157 20009 3191 20043
rect 4537 19941 4571 19975
rect 1777 19873 1811 19907
rect 2421 19873 2455 19907
rect 2973 19873 3007 19907
rect 2605 19737 2639 19771
rect 4353 19737 4387 19771
rect 1685 19669 1719 19703
rect 3525 19669 3559 19703
rect 4537 19669 4571 19703
rect 4721 19669 4755 19703
rect 1961 19465 1995 19499
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 2881 19261 2915 19295
rect 3157 19261 3191 19295
rect 5089 19261 5123 19295
rect 3985 19193 4019 19227
rect 4445 19193 4479 19227
rect 5549 19193 5583 19227
rect 1593 19125 1627 19159
rect 2513 19125 2547 19159
rect 3617 19125 3651 19159
rect 4721 19125 4755 19159
rect 5917 19125 5951 19159
rect 1777 18921 1811 18955
rect 3433 18921 3467 18955
rect 2421 18853 2455 18887
rect 3157 18853 3191 18887
rect 1593 18785 1627 18819
rect 2145 18785 2179 18819
rect 2881 18785 2915 18819
rect 3433 18717 3467 18751
rect 5181 18785 5215 18819
rect 5733 18717 5767 18751
rect 4997 18649 5031 18683
rect 5181 18649 5215 18683
rect 5457 18649 5491 18683
rect 3709 18581 3743 18615
rect 4261 18581 4295 18615
rect 4721 18581 4755 18615
rect 6193 18581 6227 18615
rect 6469 18581 6503 18615
rect 9229 18581 9263 18615
rect 1961 18377 1995 18411
rect 2513 18377 2547 18411
rect 3709 18377 3743 18411
rect 5549 18377 5583 18411
rect 6193 18309 6227 18343
rect 4721 18241 4755 18275
rect 9413 18241 9447 18275
rect 11069 18241 11103 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 6561 18173 6595 18207
rect 7113 18173 7147 18207
rect 7757 18173 7791 18207
rect 9229 18173 9263 18207
rect 10885 18173 10919 18207
rect 5089 18105 5123 18139
rect 8033 18105 8067 18139
rect 1593 18037 1627 18071
rect 2881 18037 2915 18071
rect 3341 18037 3375 18071
rect 3985 18037 4019 18071
rect 4353 18037 4387 18071
rect 5917 18037 5951 18071
rect 7481 18037 7515 18071
rect 8493 18037 8527 18071
rect 10241 18037 10275 18071
rect 10609 18037 10643 18071
rect 11713 18037 11747 18071
rect 1961 17833 1995 17867
rect 6377 17833 6411 17867
rect 9873 17833 9907 17867
rect 2605 17765 2639 17799
rect 6745 17765 6779 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 5273 17697 5307 17731
rect 10241 17697 10275 17731
rect 10885 17697 10919 17731
rect 4997 17629 5031 17663
rect 10333 17629 10367 17663
rect 10517 17629 10551 17663
rect 3065 17561 3099 17595
rect 5641 17561 5675 17595
rect 7849 17561 7883 17595
rect 8309 17561 8343 17595
rect 9045 17561 9079 17595
rect 9413 17561 9447 17595
rect 11345 17561 11379 17595
rect 11805 17561 11839 17595
rect 13093 17561 13127 17595
rect 1685 17493 1719 17527
rect 3433 17493 3467 17527
rect 3801 17493 3835 17527
rect 4629 17493 4663 17527
rect 6101 17493 6135 17527
rect 7113 17493 7147 17527
rect 7481 17493 7515 17527
rect 8769 17493 8803 17527
rect 12725 17493 12759 17527
rect 1869 17289 1903 17323
rect 2881 17289 2915 17323
rect 9873 17289 9907 17323
rect 11345 17289 11379 17323
rect 11621 17289 11655 17323
rect 2421 17153 2455 17187
rect 6561 17221 6595 17255
rect 13829 17221 13863 17255
rect 1685 17085 1719 17119
rect 2237 17085 2271 17119
rect 2881 17085 2915 17119
rect 2973 17085 3007 17119
rect 3249 17085 3283 17119
rect 4261 17085 4295 17119
rect 6837 17085 6871 17119
rect 7093 17085 7127 17119
rect 9965 17085 9999 17119
rect 12449 17085 12483 17119
rect 12716 17085 12750 17119
rect 4506 17017 4540 17051
rect 10210 17017 10244 17051
rect 11989 17017 12023 17051
rect 3801 16949 3835 16983
rect 5641 16949 5675 16983
rect 6009 16949 6043 16983
rect 8217 16949 8251 16983
rect 8585 16949 8619 16983
rect 9137 16949 9171 16983
rect 9505 16949 9539 16983
rect 1961 16745 1995 16779
rect 3249 16745 3283 16779
rect 3801 16745 3835 16779
rect 5457 16745 5491 16779
rect 7113 16745 7147 16779
rect 8309 16745 8343 16779
rect 8769 16745 8803 16779
rect 11069 16745 11103 16779
rect 13001 16745 13035 16779
rect 5978 16677 6012 16711
rect 7757 16677 7791 16711
rect 1777 16609 1811 16643
rect 2329 16609 2363 16643
rect 2605 16609 2639 16643
rect 3065 16609 3099 16643
rect 4077 16609 4111 16643
rect 4333 16609 4367 16643
rect 5733 16609 5767 16643
rect 8217 16609 8251 16643
rect 8677 16609 8711 16643
rect 9956 16609 9990 16643
rect 11612 16609 11646 16643
rect 13369 16609 13403 16643
rect 13461 16609 13495 16643
rect 8953 16541 8987 16575
rect 9689 16541 9723 16575
rect 11345 16541 11379 16575
rect 13645 16541 13679 16575
rect 9413 16473 9447 16507
rect 12725 16473 12759 16507
rect 1685 16405 1719 16439
rect 7481 16405 7515 16439
rect 1777 16201 1811 16235
rect 2973 16201 3007 16235
rect 3433 16201 3467 16235
rect 4445 16201 4479 16235
rect 6837 16201 6871 16235
rect 9781 16201 9815 16235
rect 10793 16201 10827 16235
rect 12909 16201 12943 16235
rect 13461 16201 13495 16235
rect 5641 16133 5675 16167
rect 9505 16133 9539 16167
rect 12173 16133 12207 16167
rect 2329 16065 2363 16099
rect 3893 16065 3927 16099
rect 3985 16065 4019 16099
rect 4997 16065 5031 16099
rect 6101 16065 6135 16099
rect 6285 16065 6319 16099
rect 7389 16065 7423 16099
rect 8125 16065 8159 16099
rect 10425 16065 10459 16099
rect 11345 16065 11379 16099
rect 12449 16065 12483 16099
rect 13737 16065 13771 16099
rect 1593 15997 1627 16031
rect 2145 15997 2179 16031
rect 3801 15997 3835 16031
rect 6009 15997 6043 16031
rect 8392 15997 8426 16031
rect 3341 15929 3375 15963
rect 4905 15929 4939 15963
rect 5549 15929 5583 15963
rect 7205 15929 7239 15963
rect 11161 15929 11195 15963
rect 4813 15861 4847 15895
rect 7297 15861 7331 15895
rect 7849 15861 7883 15895
rect 10149 15861 10183 15895
rect 10241 15861 10275 15895
rect 11253 15861 11287 15895
rect 11897 15861 11931 15895
rect 14105 15861 14139 15895
rect 1685 15657 1719 15691
rect 5457 15657 5491 15691
rect 6009 15657 6043 15691
rect 8309 15657 8343 15691
rect 9321 15657 9355 15691
rect 11161 15657 11195 15691
rect 11529 15657 11563 15691
rect 2329 15589 2363 15623
rect 3065 15589 3099 15623
rect 4322 15589 4356 15623
rect 6193 15589 6227 15623
rect 8677 15589 8711 15623
rect 1501 15521 1535 15555
rect 2053 15521 2087 15555
rect 2789 15521 2823 15555
rect 6920 15521 6954 15555
rect 8769 15521 8803 15555
rect 10057 15521 10091 15555
rect 10149 15521 10183 15555
rect 11897 15521 11931 15555
rect 12633 15521 12667 15555
rect 4077 15453 4111 15487
rect 6653 15453 6687 15487
rect 8861 15453 8895 15487
rect 10241 15453 10275 15487
rect 11989 15453 12023 15487
rect 12173 15453 12207 15487
rect 8033 15385 8067 15419
rect 3525 15317 3559 15351
rect 9689 15317 9723 15351
rect 10701 15317 10735 15351
rect 13001 15317 13035 15351
rect 1685 15113 1719 15147
rect 5549 15113 5583 15147
rect 6009 15113 6043 15147
rect 8677 15113 8711 15147
rect 10517 15113 10551 15147
rect 12633 15113 12667 15147
rect 13369 15113 13403 15147
rect 4261 15045 4295 15079
rect 5181 15045 5215 15079
rect 7205 15045 7239 15079
rect 13001 15045 13035 15079
rect 2237 14977 2271 15011
rect 2881 14977 2915 15011
rect 6653 14977 6687 15011
rect 7849 14977 7883 15011
rect 1501 14909 1535 14943
rect 2053 14909 2087 14943
rect 3148 14909 3182 14943
rect 7021 14909 7055 14943
rect 7573 14909 7607 14943
rect 9137 14909 9171 14943
rect 9404 14909 9438 14943
rect 11161 14909 11195 14943
rect 11529 14909 11563 14943
rect 4905 14773 4939 14807
rect 7665 14773 7699 14807
rect 8217 14773 8251 14807
rect 10793 14773 10827 14807
rect 11897 14773 11931 14807
rect 1869 14569 1903 14603
rect 3157 14569 3191 14603
rect 3893 14569 3927 14603
rect 6101 14569 6135 14603
rect 9045 14569 9079 14603
rect 9689 14569 9723 14603
rect 11713 14569 11747 14603
rect 13461 14569 13495 14603
rect 6745 14501 6779 14535
rect 7288 14501 7322 14535
rect 12725 14501 12759 14535
rect 1685 14433 1719 14467
rect 2237 14433 2271 14467
rect 2513 14433 2547 14467
rect 2973 14433 3007 14467
rect 4977 14433 5011 14467
rect 10600 14433 10634 14467
rect 11989 14433 12023 14467
rect 4077 14365 4111 14399
rect 4721 14365 4755 14399
rect 7021 14365 7055 14399
rect 10333 14365 10367 14399
rect 13001 14365 13035 14399
rect 9413 14297 9447 14331
rect 13829 14297 13863 14331
rect 4629 14229 4663 14263
rect 6469 14229 6503 14263
rect 8401 14229 8435 14263
rect 8769 14229 8803 14263
rect 10149 14229 10183 14263
rect 12357 14229 12391 14263
rect 13001 14229 13035 14263
rect 13185 14229 13219 14263
rect 1961 14025 1995 14059
rect 3525 14025 3559 14059
rect 6469 14025 6503 14059
rect 7297 14025 7331 14059
rect 8309 14025 8343 14059
rect 8769 14025 8803 14059
rect 10425 14025 10459 14059
rect 14105 14025 14139 14059
rect 14473 14025 14507 14059
rect 9413 13957 9447 13991
rect 13369 13957 13403 13991
rect 2605 13889 2639 13923
rect 4169 13889 4203 13923
rect 5089 13889 5123 13923
rect 7757 13889 7791 13923
rect 7941 13889 7975 13923
rect 9873 13889 9907 13923
rect 10057 13889 10091 13923
rect 11069 13889 11103 13923
rect 12633 13889 12667 13923
rect 1777 13821 1811 13855
rect 2329 13821 2363 13855
rect 3433 13821 3467 13855
rect 3893 13821 3927 13855
rect 3985 13821 4019 13855
rect 5356 13821 5390 13855
rect 7021 13821 7055 13855
rect 8493 13821 8527 13855
rect 9781 13821 9815 13855
rect 11805 13821 11839 13855
rect 10793 13753 10827 13787
rect 12173 13753 12207 13787
rect 14933 13753 14967 13787
rect 1685 13685 1719 13719
rect 4629 13685 4663 13719
rect 7665 13685 7699 13719
rect 9137 13685 9171 13719
rect 10885 13685 10919 13719
rect 11437 13685 11471 13719
rect 13001 13685 13035 13719
rect 13829 13685 13863 13719
rect 2605 13481 2639 13515
rect 4813 13481 4847 13515
rect 5181 13481 5215 13515
rect 5825 13481 5859 13515
rect 9137 13481 9171 13515
rect 11161 13481 11195 13515
rect 12541 13481 12575 13515
rect 12909 13481 12943 13515
rect 14749 13481 14783 13515
rect 15485 13481 15519 13515
rect 1961 13413 1995 13447
rect 10048 13413 10082 13447
rect 11437 13413 11471 13447
rect 11805 13413 11839 13447
rect 13277 13413 13311 13447
rect 1685 13345 1719 13379
rect 2421 13345 2455 13379
rect 2973 13345 3007 13379
rect 3249 13345 3283 13379
rect 6193 13345 6227 13379
rect 7297 13345 7331 13379
rect 7564 13345 7598 13379
rect 5273 13277 5307 13311
rect 5365 13277 5399 13311
rect 6285 13277 6319 13311
rect 6377 13277 6411 13311
rect 9781 13277 9815 13311
rect 6837 13209 6871 13243
rect 12173 13209 12207 13243
rect 13737 13209 13771 13243
rect 3893 13141 3927 13175
rect 4353 13141 4387 13175
rect 4721 13141 4755 13175
rect 8677 13141 8711 13175
rect 8953 13141 8987 13175
rect 14105 13141 14139 13175
rect 14473 13141 14507 13175
rect 2513 12937 2547 12971
rect 4813 12937 4847 12971
rect 5549 12937 5583 12971
rect 11253 12937 11287 12971
rect 11621 12937 11655 12971
rect 11897 12937 11931 12971
rect 14473 12937 14507 12971
rect 15577 12937 15611 12971
rect 15945 12937 15979 12971
rect 4537 12869 4571 12903
rect 1685 12733 1719 12767
rect 1961 12733 1995 12767
rect 2605 12733 2639 12767
rect 9505 12869 9539 12903
rect 13369 12869 13403 12903
rect 6193 12801 6227 12835
rect 7481 12801 7515 12835
rect 8401 12801 8435 12835
rect 5457 12733 5491 12767
rect 7297 12733 7331 12767
rect 8309 12733 8343 12767
rect 2872 12665 2906 12699
rect 4537 12665 4571 12699
rect 5181 12665 5215 12699
rect 7205 12665 7239 12699
rect 8861 12665 8895 12699
rect 13737 12801 13771 12835
rect 9873 12733 9907 12767
rect 14105 12733 14139 12767
rect 9689 12665 9723 12699
rect 10140 12665 10174 12699
rect 3985 12597 4019 12631
rect 4261 12597 4295 12631
rect 5273 12597 5307 12631
rect 5917 12597 5951 12631
rect 6009 12597 6043 12631
rect 6561 12597 6595 12631
rect 6837 12597 6871 12631
rect 7849 12597 7883 12631
rect 8217 12597 8251 12631
rect 9321 12597 9355 12631
rect 9505 12597 9539 12631
rect 12633 12597 12667 12631
rect 13093 12597 13127 12631
rect 14933 12597 14967 12631
rect 15301 12597 15335 12631
rect 16405 12597 16439 12631
rect 1593 12393 1627 12427
rect 1961 12393 1995 12427
rect 3341 12393 3375 12427
rect 4445 12393 4479 12427
rect 6653 12393 6687 12427
rect 9689 12393 9723 12427
rect 10057 12393 10091 12427
rect 11437 12393 11471 12427
rect 12541 12393 12575 12427
rect 15025 12393 15059 12427
rect 16957 12393 16991 12427
rect 2421 12325 2455 12359
rect 3801 12325 3835 12359
rect 5518 12325 5552 12359
rect 7021 12325 7055 12359
rect 7472 12325 7506 12359
rect 10149 12325 10183 12359
rect 12817 12325 12851 12359
rect 1409 12257 1443 12291
rect 2329 12257 2363 12291
rect 2605 12189 2639 12223
rect 3433 12189 3467 12223
rect 3525 12189 3559 12223
rect 2973 12121 3007 12155
rect 4537 12257 4571 12291
rect 4997 12257 5031 12291
rect 10701 12257 10735 12291
rect 12173 12257 12207 12291
rect 4629 12189 4663 12223
rect 5273 12189 5307 12223
rect 7205 12189 7239 12223
rect 8861 12189 8895 12223
rect 10333 12189 10367 12223
rect 13185 12189 13219 12223
rect 4997 12121 5031 12155
rect 11897 12121 11931 12155
rect 13921 12121 13955 12155
rect 14289 12121 14323 12155
rect 15945 12121 15979 12155
rect 19073 12121 19107 12155
rect 3801 12053 3835 12087
rect 4077 12053 4111 12087
rect 5089 12053 5123 12087
rect 8585 12053 8619 12087
rect 9413 12053 9447 12087
rect 11069 12053 11103 12087
rect 11989 12053 12023 12087
rect 13553 12053 13587 12087
rect 14657 12053 14691 12087
rect 15485 12053 15519 12087
rect 16313 12053 16347 12087
rect 16589 12053 16623 12087
rect 17417 12053 17451 12087
rect 1777 11849 1811 11883
rect 2881 11849 2915 11883
rect 6469 11849 6503 11883
rect 7113 11849 7147 11883
rect 8585 11849 8619 11883
rect 9045 11849 9079 11883
rect 15577 11849 15611 11883
rect 7389 11781 7423 11815
rect 2329 11713 2363 11747
rect 8033 11713 8067 11747
rect 2145 11645 2179 11679
rect 3341 11645 3375 11679
rect 5089 11645 5123 11679
rect 7297 11645 7331 11679
rect 9965 11781 9999 11815
rect 11437 11781 11471 11815
rect 9505 11713 9539 11747
rect 9689 11713 9723 11747
rect 14473 11713 14507 11747
rect 1685 11577 1719 11611
rect 3608 11577 3642 11611
rect 5356 11577 5390 11611
rect 7849 11577 7883 11611
rect 8401 11577 8435 11611
rect 8585 11577 8619 11611
rect 9873 11645 9907 11679
rect 9965 11645 9999 11679
rect 10057 11645 10091 11679
rect 10324 11645 10358 11679
rect 12633 11645 12667 11679
rect 15209 11645 15243 11679
rect 19073 11645 19107 11679
rect 19625 11645 19659 11679
rect 20177 11645 20211 11679
rect 14841 11577 14875 11611
rect 16313 11577 16347 11611
rect 17049 11577 17083 11611
rect 17417 11577 17451 11611
rect 17785 11577 17819 11611
rect 2237 11509 2271 11543
rect 3249 11509 3283 11543
rect 4721 11509 4755 11543
rect 7757 11509 7791 11543
rect 8769 11509 8803 11543
rect 9413 11509 9447 11543
rect 9873 11509 9907 11543
rect 11713 11509 11747 11543
rect 12081 11509 12115 11543
rect 13093 11509 13127 11543
rect 13461 11509 13495 11543
rect 13737 11509 13771 11543
rect 14105 11509 14139 11543
rect 15945 11509 15979 11543
rect 16681 11509 16715 11543
rect 19257 11509 19291 11543
rect 19809 11509 19843 11543
rect 3157 11305 3191 11339
rect 4813 11305 4847 11339
rect 5181 11305 5215 11339
rect 6745 11305 6779 11339
rect 7113 11305 7147 11339
rect 9229 11305 9263 11339
rect 11345 11305 11379 11339
rect 12909 11305 12943 11339
rect 16221 11305 16255 11339
rect 17325 11305 17359 11339
rect 2044 11237 2078 11271
rect 5641 11237 5675 11271
rect 7481 11237 7515 11271
rect 9956 11237 9990 11271
rect 13645 11237 13679 11271
rect 3617 11169 3651 11203
rect 4537 11169 4571 11203
rect 5549 11169 5583 11203
rect 7573 11169 7607 11203
rect 7840 11169 7874 11203
rect 16589 11169 16623 11203
rect 16957 11169 16991 11203
rect 18521 11169 18555 11203
rect 1777 11101 1811 11135
rect 5733 11101 5767 11135
rect 6193 11101 6227 11135
rect 9689 11101 9723 11135
rect 14749 11101 14783 11135
rect 18061 11101 18095 11135
rect 8953 11033 8987 11067
rect 11069 11033 11103 11067
rect 11897 11033 11931 11067
rect 13369 11033 13403 11067
rect 14381 11033 14415 11067
rect 15945 11033 15979 11067
rect 17693 11033 17727 11067
rect 18705 11033 18739 11067
rect 1685 10965 1719 10999
rect 12265 10965 12299 10999
rect 12633 10965 12667 10999
rect 14013 10965 14047 10999
rect 15577 10965 15611 10999
rect 2881 10761 2915 10795
rect 6377 10761 6411 10795
rect 7573 10761 7607 10795
rect 8401 10761 8435 10795
rect 10241 10761 10275 10795
rect 13921 10761 13955 10795
rect 17233 10761 17267 10795
rect 19809 10761 19843 10795
rect 3157 10693 3191 10727
rect 1501 10625 1535 10659
rect 3709 10625 3743 10659
rect 4721 10625 4755 10659
rect 7113 10625 7147 10659
rect 8217 10625 8251 10659
rect 9965 10693 9999 10727
rect 14289 10693 14323 10727
rect 15025 10693 15059 10727
rect 19073 10693 19107 10727
rect 19441 10693 19475 10727
rect 10885 10625 10919 10659
rect 15761 10625 15795 10659
rect 17601 10625 17635 10659
rect 1768 10557 1802 10591
rect 8401 10557 8435 10591
rect 8493 10557 8527 10591
rect 8585 10557 8619 10591
rect 8852 10557 8886 10591
rect 11437 10557 11471 10591
rect 14657 10557 14691 10591
rect 18153 10557 18187 10591
rect 18705 10557 18739 10591
rect 3617 10489 3651 10523
rect 4988 10489 5022 10523
rect 10701 10489 10735 10523
rect 11713 10489 11747 10523
rect 16129 10489 16163 10523
rect 3525 10421 3559 10455
rect 4261 10421 4295 10455
rect 6101 10421 6135 10455
rect 7941 10421 7975 10455
rect 8033 10421 8067 10455
rect 8493 10421 8527 10455
rect 10609 10421 10643 10455
rect 11253 10421 11287 10455
rect 12081 10421 12115 10455
rect 12909 10421 12943 10455
rect 13277 10421 13311 10455
rect 13553 10421 13587 10455
rect 15393 10421 15427 10455
rect 16589 10421 16623 10455
rect 16957 10421 16991 10455
rect 18337 10421 18371 10455
rect 2145 10217 2179 10251
rect 2513 10217 2547 10251
rect 3157 10217 3191 10251
rect 3617 10217 3651 10251
rect 5733 10217 5767 10251
rect 6101 10217 6135 10251
rect 8493 10217 8527 10251
rect 13553 10217 13587 10251
rect 13829 10217 13863 10251
rect 14013 10217 14047 10251
rect 7021 10149 7055 10183
rect 1685 10081 1719 10115
rect 2053 10081 2087 10115
rect 4344 10081 4378 10115
rect 6193 10081 6227 10115
rect 6745 10081 6779 10115
rect 8677 10081 8711 10115
rect 9321 10081 9355 10115
rect 10333 10081 10367 10115
rect 12173 10081 12207 10115
rect 12440 10081 12474 10115
rect 2605 10013 2639 10047
rect 2697 10013 2731 10047
rect 4077 10013 4111 10047
rect 6285 10013 6319 10047
rect 8033 10013 8067 10047
rect 14749 10217 14783 10251
rect 15025 10217 15059 10251
rect 17325 10217 17359 10251
rect 17785 10217 17819 10251
rect 18061 10217 18095 10251
rect 19165 10217 19199 10251
rect 19533 10217 19567 10251
rect 19901 10217 19935 10251
rect 20269 10217 20303 10251
rect 14657 9945 14691 9979
rect 16957 10149 16991 10183
rect 18429 10149 18463 10183
rect 18797 10149 18831 10183
rect 15485 10013 15519 10047
rect 5457 9877 5491 9911
rect 7481 9877 7515 9911
rect 7849 9877 7883 9911
rect 8953 9877 8987 9911
rect 9137 9877 9171 9911
rect 9965 9877 9999 9911
rect 11805 9877 11839 9911
rect 14013 9877 14047 9911
rect 14197 9877 14231 9911
rect 14749 9877 14783 9911
rect 15853 9877 15887 9911
rect 16313 9877 16347 9911
rect 16589 9877 16623 9911
rect 2329 9673 2363 9707
rect 18613 9673 18647 9707
rect 18981 9673 19015 9707
rect 20453 9673 20487 9707
rect 1777 9605 1811 9639
rect 4629 9605 4663 9639
rect 5641 9605 5675 9639
rect 7021 9605 7055 9639
rect 7205 9605 7239 9639
rect 9505 9605 9539 9639
rect 18245 9605 18279 9639
rect 20821 9605 20855 9639
rect 21189 9605 21223 9639
rect 2973 9537 3007 9571
rect 5181 9537 5215 9571
rect 6193 9537 6227 9571
rect 7757 9537 7791 9571
rect 8217 9537 8251 9571
rect 9045 9537 9079 9571
rect 10149 9537 10183 9571
rect 11897 9537 11931 9571
rect 13001 9537 13035 9571
rect 17049 9537 17083 9571
rect 2789 9469 2823 9503
rect 3433 9469 3467 9503
rect 3801 9469 3835 9503
rect 8861 9469 8895 9503
rect 11069 9469 11103 9503
rect 11713 9469 11747 9503
rect 13277 9469 13311 9503
rect 13921 9469 13955 9503
rect 14188 9469 14222 9503
rect 15945 9469 15979 9503
rect 16681 9469 16715 9503
rect 4537 9401 4571 9435
rect 6101 9401 6135 9435
rect 7665 9401 7699 9435
rect 9965 9401 9999 9435
rect 10517 9401 10551 9435
rect 12817 9401 12851 9435
rect 13461 9401 13495 9435
rect 17417 9401 17451 9435
rect 19441 9401 19475 9435
rect 19809 9401 19843 9435
rect 2145 9333 2179 9367
rect 2697 9333 2731 9367
rect 4077 9333 4111 9367
rect 4997 9333 5031 9367
rect 5089 9333 5123 9367
rect 6009 9333 6043 9367
rect 7573 9333 7607 9367
rect 8493 9333 8527 9367
rect 8953 9333 8987 9367
rect 9873 9333 9907 9367
rect 11253 9333 11287 9367
rect 11621 9333 11655 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 13277 9333 13311 9367
rect 15301 9333 15335 9367
rect 15669 9333 15703 9367
rect 16405 9333 16439 9367
rect 17785 9333 17819 9367
rect 20085 9333 20119 9367
rect 1685 9129 1719 9163
rect 4261 9129 4295 9163
rect 4905 9129 4939 9163
rect 7941 9129 7975 9163
rect 8677 9129 8711 9163
rect 9321 9129 9355 9163
rect 9505 9129 9539 9163
rect 14933 9129 14967 9163
rect 19441 9129 19475 9163
rect 2044 9061 2078 9095
rect 6806 9061 6840 9095
rect 8769 9061 8803 9095
rect 9137 9061 9171 9095
rect 1777 8993 1811 9027
rect 4813 8993 4847 9027
rect 5457 8993 5491 9027
rect 6561 8993 6595 9027
rect 3433 8925 3467 8959
rect 5089 8925 5123 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9956 9061 9990 9095
rect 12164 9061 12198 9095
rect 17601 9061 17635 9095
rect 19809 9061 19843 9095
rect 20177 9061 20211 9095
rect 11897 8993 11931 9027
rect 13553 8993 13587 9027
rect 13820 8993 13854 9027
rect 17233 8993 17267 9027
rect 9689 8925 9723 8959
rect 15301 8925 15335 8959
rect 16129 8925 16163 8959
rect 3801 8857 3835 8891
rect 6377 8857 6411 8891
rect 8309 8857 8343 8891
rect 9505 8857 9539 8891
rect 11713 8857 11747 8891
rect 16865 8857 16899 8891
rect 18061 8857 18095 8891
rect 3157 8789 3191 8823
rect 4445 8789 4479 8823
rect 6009 8789 6043 8823
rect 11069 8789 11103 8823
rect 13277 8789 13311 8823
rect 15761 8789 15795 8823
rect 16589 8789 16623 8823
rect 18429 8789 18463 8823
rect 18705 8789 18739 8823
rect 19073 8789 19107 8823
rect 20637 8789 20671 8823
rect 21189 8789 21223 8823
rect 1869 8585 1903 8619
rect 2145 8585 2179 8619
rect 2513 8585 2547 8619
rect 5273 8585 5307 8619
rect 8493 8585 8527 8619
rect 11621 8585 11655 8619
rect 11897 8585 11931 8619
rect 13369 8585 13403 8619
rect 13553 8585 13587 8619
rect 15393 8585 15427 8619
rect 15577 8585 15611 8619
rect 19717 8585 19751 8619
rect 20545 8585 20579 8619
rect 20821 8585 20855 8619
rect 21189 8585 21223 8619
rect 2697 8517 2731 8551
rect 6561 8517 6595 8551
rect 8217 8517 8251 8551
rect 9689 8517 9723 8551
rect 3157 8449 3191 8483
rect 3249 8449 3283 8483
rect 6009 8449 6043 8483
rect 6193 8449 6227 8483
rect 9137 8449 9171 8483
rect 9505 8449 9539 8483
rect 10241 8449 10275 8483
rect 11529 8449 11563 8483
rect 3893 8381 3927 8415
rect 4160 8381 4194 8415
rect 5457 8381 5491 8415
rect 6837 8381 6871 8415
rect 7104 8381 7138 8415
rect 8861 8381 8895 8415
rect 10149 8381 10183 8415
rect 10701 8381 10735 8415
rect 11805 8381 11839 8415
rect 3801 8313 3835 8347
rect 13093 8517 13127 8551
rect 12449 8449 12483 8483
rect 14197 8449 14231 8483
rect 15117 8449 15151 8483
rect 18981 8517 19015 8551
rect 20085 8517 20119 8551
rect 17417 8449 17451 8483
rect 18613 8449 18647 8483
rect 12081 8381 12115 8415
rect 13921 8381 13955 8415
rect 14933 8381 14967 8415
rect 15393 8381 15427 8415
rect 16405 8381 16439 8415
rect 17141 8381 17175 8415
rect 10057 8313 10091 8347
rect 11069 8313 11103 8347
rect 11897 8313 11931 8347
rect 16681 8313 16715 8347
rect 19349 8313 19383 8347
rect 3065 8245 3099 8279
rect 5457 8245 5491 8279
rect 5549 8245 5583 8279
rect 5917 8245 5951 8279
rect 8953 8245 8987 8279
rect 14013 8245 14047 8279
rect 14565 8245 14599 8279
rect 15025 8245 15059 8279
rect 16037 8245 16071 8279
rect 18337 8245 18371 8279
rect 3065 8041 3099 8075
rect 4353 8041 4387 8075
rect 4813 8041 4847 8075
rect 7113 8041 7147 8075
rect 8861 8041 8895 8075
rect 15025 8041 15059 8075
rect 17325 8041 17359 8075
rect 21097 8041 21131 8075
rect 5724 7973 5758 8007
rect 17969 7973 18003 8007
rect 1952 7905 1986 7939
rect 5365 7905 5399 7939
rect 5457 7905 5491 7939
rect 7297 7905 7331 7939
rect 11152 7905 11186 7939
rect 16201 7905 16235 7939
rect 20545 7905 20579 7939
rect 1685 7837 1719 7871
rect 4905 7837 4939 7871
rect 5089 7837 5123 7871
rect 10885 7837 10919 7871
rect 12541 7837 12575 7871
rect 12909 7837 12943 7871
rect 15945 7837 15979 7871
rect 19073 7837 19107 7871
rect 8585 7769 8619 7803
rect 9229 7769 9263 7803
rect 10057 7769 10091 7803
rect 13369 7769 13403 7803
rect 14013 7769 14047 7803
rect 18337 7769 18371 7803
rect 3525 7701 3559 7735
rect 3801 7701 3835 7735
rect 4445 7701 4479 7735
rect 5365 7701 5399 7735
rect 6837 7701 6871 7735
rect 7573 7701 7607 7735
rect 7941 7701 7975 7735
rect 10793 7701 10827 7735
rect 12265 7701 12299 7735
rect 12817 7701 12851 7735
rect 13001 7701 13035 7735
rect 14565 7701 14599 7735
rect 15853 7701 15887 7735
rect 17601 7701 17635 7735
rect 18705 7701 18739 7735
rect 19533 7701 19567 7735
rect 19809 7701 19843 7735
rect 20177 7701 20211 7735
rect 3065 7497 3099 7531
rect 4077 7497 4111 7531
rect 5089 7497 5123 7531
rect 9045 7497 9079 7531
rect 15577 7497 15611 7531
rect 16313 7497 16347 7531
rect 18521 7497 18555 7531
rect 18613 7497 18647 7531
rect 19349 7497 19383 7531
rect 2053 7429 2087 7463
rect 6469 7429 6503 7463
rect 12449 7429 12483 7463
rect 2513 7361 2547 7395
rect 2697 7361 2731 7395
rect 3617 7361 3651 7395
rect 3893 7361 3927 7395
rect 4537 7361 4571 7395
rect 4721 7361 4755 7395
rect 5641 7361 5675 7395
rect 7665 7361 7699 7395
rect 9321 7361 9355 7395
rect 11621 7361 11655 7395
rect 13093 7361 13127 7395
rect 16957 7361 16991 7395
rect 2421 7225 2455 7259
rect 3525 7225 3559 7259
rect 20821 7429 20855 7463
rect 20453 7361 20487 7395
rect 5549 7293 5583 7327
rect 6101 7293 6135 7327
rect 12817 7293 12851 7327
rect 13461 7293 13495 7327
rect 14197 7293 14231 7327
rect 16129 7293 16163 7327
rect 16773 7293 16807 7327
rect 18521 7293 18555 7327
rect 18981 7293 19015 7327
rect 4445 7225 4479 7259
rect 7932 7225 7966 7259
rect 9577 7225 9611 7259
rect 14464 7225 14498 7259
rect 16681 7225 16715 7259
rect 21189 7225 21223 7259
rect 1869 7157 1903 7191
rect 3433 7157 3467 7191
rect 3893 7157 3927 7191
rect 5457 7157 5491 7191
rect 7205 7157 7239 7191
rect 10701 7157 10735 7191
rect 10977 7157 11011 7191
rect 11345 7157 11379 7191
rect 11437 7157 11471 7191
rect 11989 7157 12023 7191
rect 12909 7157 12943 7191
rect 14013 7157 14047 7191
rect 17325 7157 17359 7191
rect 17785 7157 17819 7191
rect 18245 7157 18279 7191
rect 19717 7157 19751 7191
rect 20085 7157 20119 7191
rect 2789 6953 2823 6987
rect 2881 6953 2915 6987
rect 1676 6885 1710 6919
rect 1409 6749 1443 6783
rect 2881 6749 2915 6783
rect 2973 6953 3007 6987
rect 3157 6953 3191 6987
rect 6653 6953 6687 6987
rect 7573 6953 7607 6987
rect 8493 6953 8527 6987
rect 9045 6953 9079 6987
rect 9413 6953 9447 6987
rect 10517 6953 10551 6987
rect 17785 6953 17819 6987
rect 18153 6953 18187 6987
rect 3433 6817 3467 6851
rect 3893 6817 3927 6851
rect 4445 6817 4479 6851
rect 4537 6817 4571 6851
rect 5273 6817 5307 6851
rect 6193 6817 6227 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 4721 6749 4755 6783
rect 5549 6749 5583 6783
rect 7757 6749 7791 6783
rect 8953 6817 8987 6851
rect 9137 6749 9171 6783
rect 2973 6681 3007 6715
rect 4077 6681 4111 6715
rect 5089 6681 5123 6715
rect 7205 6681 7239 6715
rect 8493 6681 8527 6715
rect 11161 6885 11195 6919
rect 9689 6817 9723 6851
rect 10701 6817 10735 6851
rect 11612 6817 11646 6851
rect 13185 6817 13219 6851
rect 13461 6817 13495 6851
rect 13728 6817 13762 6851
rect 15301 6817 15335 6851
rect 15853 6817 15887 6851
rect 16304 6817 16338 6851
rect 18797 6817 18831 6851
rect 20269 6817 20303 6851
rect 11345 6749 11379 6783
rect 12817 6749 12851 6783
rect 15485 6749 15519 6783
rect 9413 6681 9447 6715
rect 16037 6749 16071 6783
rect 18429 6749 18463 6783
rect 20729 6749 20763 6783
rect 19901 6681 19935 6715
rect 6009 6613 6043 6647
rect 7021 6613 7055 6647
rect 8585 6613 8619 6647
rect 10149 6613 10183 6647
rect 12725 6613 12759 6647
rect 12817 6613 12851 6647
rect 13001 6613 13035 6647
rect 14841 6613 14875 6647
rect 15853 6613 15887 6647
rect 17417 6613 17451 6647
rect 19165 6613 19199 6647
rect 19533 6613 19567 6647
rect 21097 6613 21131 6647
rect 1685 6409 1719 6443
rect 3617 6409 3651 6443
rect 19349 6409 19383 6443
rect 5549 6341 5583 6375
rect 10057 6341 10091 6375
rect 11713 6341 11747 6375
rect 13829 6341 13863 6375
rect 16221 6341 16255 6375
rect 20821 6341 20855 6375
rect 1777 6273 1811 6307
rect 6193 6273 6227 6307
rect 7389 6273 7423 6307
rect 10333 6273 10367 6307
rect 12449 6273 12483 6307
rect 14749 6273 14783 6307
rect 15669 6273 15703 6307
rect 15853 6273 15887 6307
rect 16865 6273 16899 6307
rect 18245 6273 18279 6307
rect 19717 6273 19751 6307
rect 2237 6205 2271 6239
rect 4169 6205 4203 6239
rect 4436 6205 4470 6239
rect 6285 6205 6319 6239
rect 7205 6205 7239 6239
rect 8309 6205 8343 6239
rect 10241 6205 10275 6239
rect 15577 6205 15611 6239
rect 16589 6205 16623 6239
rect 18797 6205 18831 6239
rect 20085 6205 20119 6239
rect 2504 6137 2538 6171
rect 7297 6137 7331 6171
rect 8576 6137 8610 6171
rect 10578 6137 10612 6171
rect 12716 6137 12750 6171
rect 14473 6137 14507 6171
rect 20453 6137 20487 6171
rect 3985 6069 4019 6103
rect 6837 6069 6871 6103
rect 7849 6069 7883 6103
rect 9689 6069 9723 6103
rect 10241 6069 10275 6103
rect 12081 6069 12115 6103
rect 14105 6069 14139 6103
rect 14565 6069 14599 6103
rect 15209 6069 15243 6103
rect 16681 6069 16715 6103
rect 17325 6069 17359 6103
rect 17693 6069 17727 6103
rect 18613 6069 18647 6103
rect 18797 6069 18831 6103
rect 18981 6069 19015 6103
rect 21189 6069 21223 6103
rect 1961 5865 1995 5899
rect 2421 5865 2455 5899
rect 3525 5865 3559 5899
rect 6929 5865 6963 5899
rect 8953 5865 8987 5899
rect 9505 5865 9539 5899
rect 11069 5865 11103 5899
rect 13001 5865 13035 5899
rect 14105 5865 14139 5899
rect 19441 5865 19475 5899
rect 5457 5797 5491 5831
rect 2789 5729 2823 5763
rect 4445 5729 4479 5763
rect 5549 5729 5583 5763
rect 5816 5729 5850 5763
rect 7461 5729 7495 5763
rect 2881 5661 2915 5695
rect 2973 5661 3007 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 7205 5661 7239 5695
rect 10057 5797 10091 5831
rect 11621 5797 11655 5831
rect 11805 5797 11839 5831
rect 12357 5797 12391 5831
rect 16313 5797 16347 5831
rect 18337 5797 18371 5831
rect 18705 5797 18739 5831
rect 19073 5797 19107 5831
rect 11161 5729 11195 5763
rect 13369 5729 13403 5763
rect 14473 5729 14507 5763
rect 15669 5729 15703 5763
rect 15945 5729 15979 5763
rect 16681 5729 16715 5763
rect 16948 5729 16982 5763
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 11253 5661 11287 5695
rect 11621 5661 11655 5695
rect 12449 5661 12483 5695
rect 12633 5661 12667 5695
rect 13645 5661 13679 5695
rect 14565 5661 14599 5695
rect 14657 5661 14691 5695
rect 20545 5661 20579 5695
rect 9505 5593 9539 5627
rect 10701 5593 10735 5627
rect 18061 5593 18095 5627
rect 20177 5593 20211 5627
rect 2329 5525 2363 5559
rect 3801 5525 3835 5559
rect 4077 5525 4111 5559
rect 8585 5525 8619 5559
rect 9321 5525 9355 5559
rect 9689 5525 9723 5559
rect 11989 5525 12023 5559
rect 15485 5525 15519 5559
rect 19809 5525 19843 5559
rect 21097 5525 21131 5559
rect 3801 5321 3835 5355
rect 5181 5321 5215 5355
rect 7941 5321 7975 5355
rect 13921 5321 13955 5355
rect 15209 5321 15243 5355
rect 17417 5321 17451 5355
rect 18245 5321 18279 5355
rect 18981 5321 19015 5355
rect 19349 5321 19383 5355
rect 4813 5253 4847 5287
rect 7021 5253 7055 5287
rect 4445 5185 4479 5219
rect 6193 5185 6227 5219
rect 6285 5185 6319 5219
rect 7573 5185 7607 5219
rect 6101 5117 6135 5151
rect 1869 5049 1903 5083
rect 3617 5049 3651 5083
rect 4169 5049 4203 5083
rect 7389 5049 7423 5083
rect 10885 5253 10919 5287
rect 19717 5253 19751 5287
rect 8493 5185 8527 5219
rect 8585 5185 8619 5219
rect 11621 5185 11655 5219
rect 11805 5185 11839 5219
rect 12909 5185 12943 5219
rect 14749 5185 14783 5219
rect 15577 5185 15611 5219
rect 8861 5117 8895 5151
rect 9505 5117 9539 5151
rect 9772 5117 9806 5151
rect 12449 5117 12483 5151
rect 14013 5117 14047 5151
rect 16037 5117 16071 5151
rect 20453 5117 20487 5151
rect 9045 5049 9079 5083
rect 11529 5049 11563 5083
rect 13277 5049 13311 5083
rect 14289 5049 14323 5083
rect 16304 5049 16338 5083
rect 20821 5049 20855 5083
rect 2237 4981 2271 5015
rect 2789 4981 2823 5015
rect 3157 4981 3191 5015
rect 4261 4981 4295 5015
rect 5549 4981 5583 5015
rect 5733 4981 5767 5015
rect 7481 4981 7515 5015
rect 7941 4981 7975 5015
rect 8033 4981 8067 5015
rect 8401 4981 8435 5015
rect 8861 4981 8895 5015
rect 11161 4981 11195 5015
rect 12173 4981 12207 5015
rect 17785 4981 17819 5015
rect 18613 4981 18647 5015
rect 20085 4981 20119 5015
rect 21281 4981 21315 5015
rect 21741 4981 21775 5015
rect 1777 4777 1811 4811
rect 2237 4777 2271 4811
rect 3157 4777 3191 4811
rect 3801 4777 3835 4811
rect 5181 4777 5215 4811
rect 6377 4777 6411 4811
rect 6745 4777 6779 4811
rect 7389 4777 7423 4811
rect 10057 4777 10091 4811
rect 10241 4777 10275 4811
rect 14473 4777 14507 4811
rect 14933 4777 14967 4811
rect 17417 4777 17451 4811
rect 18981 4777 19015 4811
rect 20545 4777 20579 4811
rect 10968 4709 11002 4743
rect 12624 4709 12658 4743
rect 18337 4709 18371 4743
rect 1685 4641 1719 4675
rect 2145 4641 2179 4675
rect 3249 4641 3283 4675
rect 4905 4641 4939 4675
rect 5733 4641 5767 4675
rect 7757 4641 7791 4675
rect 10701 4641 10735 4675
rect 12357 4641 12391 4675
rect 15301 4641 15335 4675
rect 15568 4641 15602 4675
rect 17325 4641 17359 4675
rect 17969 4641 18003 4675
rect 18245 4641 18279 4675
rect 2421 4573 2455 4607
rect 3433 4573 3467 4607
rect 5825 4573 5859 4607
rect 5917 4573 5951 4607
rect 6837 4573 6871 4607
rect 6929 4573 6963 4607
rect 7849 4573 7883 4607
rect 7941 4573 7975 4607
rect 14013 4573 14047 4607
rect 17509 4573 17543 4607
rect 2789 4505 2823 4539
rect 8769 4505 8803 4539
rect 12081 4505 12115 4539
rect 16681 4505 16715 4539
rect 4261 4437 4295 4471
rect 5365 4437 5399 4471
rect 8493 4437 8527 4471
rect 9137 4437 9171 4471
rect 13737 4437 13771 4471
rect 16957 4437 16991 4471
rect 18245 4437 18279 4471
rect 18521 4641 18555 4675
rect 19432 4709 19466 4743
rect 18797 4573 18831 4607
rect 18981 4573 19015 4607
rect 19165 4573 19199 4607
rect 18337 4437 18371 4471
rect 21097 4437 21131 4471
rect 3341 4233 3375 4267
rect 4997 4233 5031 4267
rect 8217 4233 8251 4267
rect 16313 4233 16347 4267
rect 18705 4233 18739 4267
rect 18981 4233 19015 4267
rect 19441 4233 19475 4267
rect 11253 4165 11287 4199
rect 16037 4165 16071 4199
rect 21741 4165 21775 4199
rect 1501 4097 1535 4131
rect 1961 4097 1995 4131
rect 5825 4097 5859 4131
rect 6837 4097 6871 4131
rect 8677 4097 8711 4131
rect 9229 4097 9263 4131
rect 9413 4097 9447 4131
rect 10425 4097 10459 4131
rect 11069 4097 11103 4131
rect 11897 4097 11931 4131
rect 13001 4097 13035 4131
rect 14657 4097 14691 4131
rect 16865 4097 16899 4131
rect 20177 4097 20211 4131
rect 3617 4029 3651 4063
rect 5641 4029 5675 4063
rect 8493 4029 8527 4063
rect 2228 3961 2262 3995
rect 3862 3961 3896 3995
rect 7082 3961 7116 3995
rect 9137 4029 9171 4063
rect 12633 4029 12667 4063
rect 13268 4029 13302 4063
rect 16773 4029 16807 4063
rect 17325 4029 17359 4063
rect 10149 3961 10183 3995
rect 14924 3961 14958 3995
rect 16681 3961 16715 3995
rect 17693 3961 17727 3995
rect 19809 3961 19843 3995
rect 5273 3893 5307 3927
rect 5733 3893 5767 3927
rect 6285 3893 6319 3927
rect 8677 3893 8711 3927
rect 8769 3893 8803 3927
rect 9781 3893 9815 3927
rect 10241 3893 10275 3927
rect 11621 3893 11655 3927
rect 11713 3893 11747 3927
rect 14381 3893 14415 3927
rect 18245 3893 18279 3927
rect 20545 3893 20579 3927
rect 20913 3893 20947 3927
rect 4077 3689 4111 3723
rect 4445 3689 4479 3723
rect 6837 3689 6871 3723
rect 9321 3689 9355 3723
rect 10425 3689 10459 3723
rect 13001 3689 13035 3723
rect 15853 3689 15887 3723
rect 17417 3689 17451 3723
rect 18153 3689 18187 3723
rect 18889 3689 18923 3723
rect 5724 3621 5758 3655
rect 8186 3621 8220 3655
rect 11621 3621 11655 3655
rect 12449 3621 12483 3655
rect 13369 3621 13403 3655
rect 17877 3621 17911 3655
rect 18521 3621 18555 3655
rect 1501 3553 1535 3587
rect 1768 3553 1802 3587
rect 3249 3553 3283 3587
rect 4537 3553 4571 3587
rect 5457 3553 5491 3587
rect 7941 3553 7975 3587
rect 10333 3553 10367 3587
rect 11897 3553 11931 3587
rect 12173 3553 12207 3587
rect 13461 3553 13495 3587
rect 14381 3553 14415 3587
rect 15025 3553 15059 3587
rect 15301 3553 15335 3587
rect 15577 3553 15611 3587
rect 15853 3553 15887 3587
rect 16681 3553 16715 3587
rect 21097 3553 21131 3587
rect 3525 3485 3559 3519
rect 4629 3485 4663 3519
rect 10517 3485 10551 3519
rect 2881 3417 2915 3451
rect 12081 3485 12115 3519
rect 13645 3485 13679 3519
rect 14473 3485 14507 3519
rect 14657 3485 14691 3519
rect 16037 3485 16071 3519
rect 16497 3485 16531 3519
rect 16865 3485 16899 3519
rect 20361 3485 20395 3519
rect 19993 3417 20027 3451
rect 5273 3349 5307 3383
rect 7481 3349 7515 3383
rect 7849 3349 7883 3383
rect 9965 3349 9999 3383
rect 10977 3349 11011 3383
rect 11897 3349 11931 3383
rect 14013 3349 14047 3383
rect 19257 3349 19291 3383
rect 19625 3349 19659 3383
rect 10149 3145 10183 3179
rect 14013 3145 14047 3179
rect 14381 3145 14415 3179
rect 15393 3145 15427 3179
rect 16313 3145 16347 3179
rect 1685 3077 1719 3111
rect 2053 3077 2087 3111
rect 2421 3077 2455 3111
rect 2881 3077 2915 3111
rect 3525 3009 3559 3043
rect 4537 3009 4571 3043
rect 6193 3009 6227 3043
rect 7665 3009 7699 3043
rect 8309 3009 8343 3043
rect 11069 3009 11103 3043
rect 16037 3009 16071 3043
rect 19165 3077 19199 3111
rect 20177 3077 20211 3111
rect 2697 2941 2731 2975
rect 3249 2941 3283 2975
rect 3801 2941 3835 2975
rect 3893 2941 3927 2975
rect 4804 2941 4838 2975
rect 7389 2941 7423 2975
rect 8033 2941 8067 2975
rect 8769 2941 8803 2975
rect 11529 2941 11563 2975
rect 12449 2941 12483 2975
rect 13185 2941 13219 2975
rect 14565 2941 14599 2975
rect 14841 2941 14875 2975
rect 15761 2941 15795 2975
rect 16313 2941 16347 2975
rect 16405 2941 16439 2975
rect 17141 2941 17175 2975
rect 17417 2941 17451 2975
rect 18067 2941 18101 2975
rect 18613 2941 18647 2975
rect 19993 2941 20027 2975
rect 20545 2941 20579 2975
rect 20913 2941 20947 2975
rect 9014 2873 9048 2907
rect 11805 2873 11839 2907
rect 12725 2873 12759 2907
rect 13461 2873 13495 2907
rect 15853 2873 15887 2907
rect 16681 2873 16715 2907
rect 19533 2873 19567 2907
rect 3341 2805 3375 2839
rect 3801 2805 3835 2839
rect 4445 2805 4479 2839
rect 5917 2805 5951 2839
rect 7021 2805 7055 2839
rect 7481 2805 7515 2839
rect 10517 2805 10551 2839
rect 10885 2805 10919 2839
rect 10977 2805 11011 2839
rect 18245 2805 18279 2839
rect 18797 2805 18831 2839
rect 20729 2805 20763 2839
rect 20913 2805 20947 2839
rect 21189 2805 21223 2839
rect 1685 2601 1719 2635
rect 2789 2601 2823 2635
rect 3341 2601 3375 2635
rect 5825 2601 5859 2635
rect 6285 2601 6319 2635
rect 9045 2601 9079 2635
rect 10241 2601 10275 2635
rect 11529 2601 11563 2635
rect 16405 2601 16439 2635
rect 2053 2533 2087 2567
rect 4344 2533 4378 2567
rect 10149 2533 10183 2567
rect 3249 2465 3283 2499
rect 4077 2465 4111 2499
rect 6193 2465 6227 2499
rect 7297 2465 7331 2499
rect 7389 2465 7423 2499
rect 7941 2465 7975 2499
rect 10793 2465 10827 2499
rect 11922 2465 11956 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16405 2465 16439 2499
rect 16589 2465 16623 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19717 2465 19751 2499
rect 19993 2465 20027 2499
rect 3525 2397 3559 2431
rect 6377 2397 6411 2431
rect 7573 2397 7607 2431
rect 9137 2397 9171 2431
rect 9229 2397 9263 2431
rect 10333 2397 10367 2431
rect 11253 2397 11287 2431
rect 20177 2397 20211 2431
rect 2881 2329 2915 2363
rect 9781 2329 9815 2363
rect 16221 2329 16255 2363
rect 17325 2329 17359 2363
rect 18521 2329 18555 2363
rect 2421 2261 2455 2295
rect 5457 2261 5491 2295
rect 6929 2261 6963 2295
rect 8309 2261 8343 2295
rect 8677 2261 8711 2295
rect 12081 2261 12115 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 13921 2261 13955 2295
rect 14473 2261 14507 2295
rect 15025 2261 15059 2295
rect 15669 2261 15703 2295
rect 16773 2261 16807 2295
rect 17877 2261 17911 2295
rect 19073 2261 19107 2295
<< metal1 >>
rect 4062 20680 4068 20732
rect 4120 20720 4126 20732
rect 5166 20720 5172 20732
rect 4120 20692 5172 20720
rect 4120 20680 4126 20692
rect 5166 20680 5172 20692
rect 5224 20680 5230 20732
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2774 20040 2780 20052
rect 1995 20012 2780 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 3142 20040 3148 20052
rect 3103 20012 3148 20040
rect 3142 20000 3148 20012
rect 3200 20000 3206 20052
rect 4525 19975 4583 19981
rect 4525 19972 4537 19975
rect 1780 19944 4537 19972
rect 1780 19913 1808 19944
rect 4525 19941 4537 19944
rect 4571 19941 4583 19975
rect 4525 19935 4583 19941
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 1765 19867 1823 19873
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 2961 19907 3019 19913
rect 2961 19873 2973 19907
rect 3007 19904 3019 19907
rect 5534 19904 5540 19916
rect 3007 19876 5540 19904
rect 3007 19873 3019 19876
rect 2961 19867 3019 19873
rect 2424 19836 2452 19867
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 3142 19836 3148 19848
rect 2424 19808 3148 19836
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 2593 19771 2651 19777
rect 2593 19737 2605 19771
rect 2639 19768 2651 19771
rect 2866 19768 2872 19780
rect 2639 19740 2872 19768
rect 2639 19737 2651 19740
rect 2593 19731 2651 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19768 4399 19771
rect 4982 19768 4988 19780
rect 4387 19740 4988 19768
rect 4387 19737 4399 19740
rect 4341 19731 4399 19737
rect 4982 19728 4988 19740
rect 5040 19728 5046 19780
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 3050 19660 3056 19712
rect 3108 19700 3114 19712
rect 3513 19703 3571 19709
rect 3513 19700 3525 19703
rect 3108 19672 3525 19700
rect 3108 19660 3114 19672
rect 3513 19669 3525 19672
rect 3559 19669 3571 19703
rect 3513 19663 3571 19669
rect 4525 19703 4583 19709
rect 4525 19669 4537 19703
rect 4571 19700 4583 19703
rect 4709 19703 4767 19709
rect 4709 19700 4721 19703
rect 4571 19672 4721 19700
rect 4571 19669 4583 19672
rect 4525 19663 4583 19669
rect 4709 19669 4721 19672
rect 4755 19700 4767 19703
rect 5626 19700 5632 19712
rect 4755 19672 5632 19700
rect 4755 19669 4767 19672
rect 4709 19663 4767 19669
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 4982 19360 4988 19372
rect 2976 19332 4988 19360
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 1854 19292 1860 19304
rect 1811 19264 1860 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 2976 19292 3004 19332
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 3142 19292 3148 19304
rect 2915 19264 3004 19292
rect 3055 19264 3148 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 3142 19252 3148 19264
rect 3200 19292 3206 19304
rect 5077 19295 5135 19301
rect 5077 19292 5089 19295
rect 3200 19264 5089 19292
rect 3200 19252 3206 19264
rect 5077 19261 5089 19264
rect 5123 19261 5135 19295
rect 9030 19292 9036 19304
rect 5077 19255 5135 19261
rect 5184 19264 9036 19292
rect 3973 19227 4031 19233
rect 3973 19224 3985 19227
rect 3160 19196 3985 19224
rect 3160 19168 3188 19196
rect 3973 19193 3985 19196
rect 4019 19193 4031 19227
rect 3973 19187 4031 19193
rect 4062 19184 4068 19236
rect 4120 19224 4126 19236
rect 4433 19227 4491 19233
rect 4433 19224 4445 19227
rect 4120 19196 4445 19224
rect 4120 19184 4126 19196
rect 4433 19193 4445 19196
rect 4479 19224 4491 19227
rect 5184 19224 5212 19264
rect 9030 19252 9036 19264
rect 9088 19252 9094 19304
rect 5534 19224 5540 19236
rect 4479 19196 5212 19224
rect 5447 19196 5540 19224
rect 4479 19193 4491 19196
rect 4433 19187 4491 19193
rect 5534 19184 5540 19196
rect 5592 19224 5598 19236
rect 6270 19224 6276 19236
rect 5592 19196 6276 19224
rect 5592 19184 5598 19196
rect 6270 19184 6276 19196
rect 6328 19184 6334 19236
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2958 19156 2964 19168
rect 2547 19128 2964 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3142 19116 3148 19168
rect 3200 19116 3206 19168
rect 3510 19116 3516 19168
rect 3568 19156 3574 19168
rect 3605 19159 3663 19165
rect 3605 19156 3617 19159
rect 3568 19128 3617 19156
rect 3568 19116 3574 19128
rect 3605 19125 3617 19128
rect 3651 19125 3663 19159
rect 4706 19156 4712 19168
rect 4667 19128 4712 19156
rect 3605 19119 3663 19125
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5902 19156 5908 19168
rect 5863 19128 5908 19156
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1765 18955 1823 18961
rect 1765 18921 1777 18955
rect 1811 18952 1823 18955
rect 3234 18952 3240 18964
rect 1811 18924 3240 18952
rect 1811 18921 1823 18924
rect 1765 18915 1823 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 4062 18952 4068 18964
rect 3467 18924 4068 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 1854 18844 1860 18896
rect 1912 18884 1918 18896
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 1912 18856 2421 18884
rect 1912 18844 1918 18856
rect 2409 18853 2421 18856
rect 2455 18884 2467 18887
rect 3050 18884 3056 18896
rect 2455 18856 3056 18884
rect 2455 18853 2467 18856
rect 2409 18847 2467 18853
rect 3050 18844 3056 18856
rect 3108 18844 3114 18896
rect 3145 18887 3203 18893
rect 3145 18853 3157 18887
rect 3191 18884 3203 18887
rect 3326 18884 3332 18896
rect 3191 18856 3332 18884
rect 3191 18853 3203 18856
rect 3145 18847 3203 18853
rect 3326 18844 3332 18856
rect 3384 18884 3390 18896
rect 4706 18884 4712 18896
rect 3384 18856 4712 18884
rect 3384 18844 3390 18856
rect 4706 18844 4712 18856
rect 4764 18844 4770 18896
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18785 1639 18819
rect 1581 18779 1639 18785
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18785 2191 18819
rect 2133 18779 2191 18785
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 5169 18819 5227 18825
rect 5169 18816 5181 18819
rect 2915 18788 5181 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 5169 18785 5181 18788
rect 5215 18785 5227 18819
rect 5169 18779 5227 18785
rect 1596 18612 1624 18779
rect 2148 18748 2176 18779
rect 3421 18751 3479 18757
rect 3421 18748 3433 18751
rect 2148 18720 3433 18748
rect 3421 18717 3433 18720
rect 3467 18717 3479 18751
rect 3602 18748 3608 18760
rect 3421 18711 3479 18717
rect 3528 18720 3608 18748
rect 2314 18640 2320 18692
rect 2372 18680 2378 18692
rect 3528 18680 3556 18720
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 3804 18720 5733 18748
rect 3804 18680 3832 18720
rect 5721 18717 5733 18720
rect 5767 18748 5779 18751
rect 9398 18748 9404 18760
rect 5767 18720 9404 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 2372 18652 3556 18680
rect 3620 18652 3832 18680
rect 2372 18640 2378 18652
rect 3620 18612 3648 18652
rect 3878 18640 3884 18692
rect 3936 18680 3942 18692
rect 4985 18683 5043 18689
rect 4985 18680 4997 18683
rect 3936 18652 4997 18680
rect 3936 18640 3942 18652
rect 4985 18649 4997 18652
rect 5031 18649 5043 18683
rect 4985 18643 5043 18649
rect 5169 18683 5227 18689
rect 5169 18649 5181 18683
rect 5215 18680 5227 18683
rect 5445 18683 5503 18689
rect 5445 18680 5457 18683
rect 5215 18652 5457 18680
rect 5215 18649 5227 18652
rect 5169 18643 5227 18649
rect 5445 18649 5457 18652
rect 5491 18680 5503 18683
rect 8938 18680 8944 18692
rect 5491 18652 8944 18680
rect 5491 18649 5503 18652
rect 5445 18643 5503 18649
rect 8938 18640 8944 18652
rect 8996 18640 9002 18692
rect 1596 18584 3648 18612
rect 3697 18615 3755 18621
rect 3697 18581 3709 18615
rect 3743 18612 3755 18615
rect 3786 18612 3792 18624
rect 3743 18584 3792 18612
rect 3743 18581 3755 18584
rect 3697 18575 3755 18581
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 4709 18615 4767 18621
rect 4709 18581 4721 18615
rect 4755 18612 4767 18615
rect 4798 18612 4804 18624
rect 4755 18584 4804 18612
rect 4755 18581 4767 18584
rect 4709 18575 4767 18581
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 6181 18615 6239 18621
rect 6181 18612 6193 18615
rect 5960 18584 6193 18612
rect 5960 18572 5966 18584
rect 6181 18581 6193 18584
rect 6227 18612 6239 18615
rect 6457 18615 6515 18621
rect 6457 18612 6469 18615
rect 6227 18584 6469 18612
rect 6227 18581 6239 18584
rect 6181 18575 6239 18581
rect 6457 18581 6469 18584
rect 6503 18612 6515 18615
rect 7466 18612 7472 18624
rect 6503 18584 7472 18612
rect 6503 18581 6515 18584
rect 6457 18575 6515 18581
rect 7466 18572 7472 18584
rect 7524 18572 7530 18624
rect 9214 18612 9220 18624
rect 9175 18584 9220 18612
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2774 18408 2780 18420
rect 2547 18380 2780 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3697 18411 3755 18417
rect 3697 18377 3709 18411
rect 3743 18408 3755 18411
rect 5074 18408 5080 18420
rect 3743 18380 5080 18408
rect 3743 18377 3755 18380
rect 3697 18371 3755 18377
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5537 18411 5595 18417
rect 5537 18377 5549 18411
rect 5583 18408 5595 18411
rect 6546 18408 6552 18420
rect 5583 18380 6552 18408
rect 5583 18377 5595 18380
rect 5537 18371 5595 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 2130 18300 2136 18352
rect 2188 18340 2194 18352
rect 6181 18343 6239 18349
rect 6181 18340 6193 18343
rect 2188 18312 6193 18340
rect 2188 18300 2194 18312
rect 6181 18309 6193 18312
rect 6227 18309 6239 18343
rect 6181 18303 6239 18309
rect 6270 18300 6276 18352
rect 6328 18340 6334 18352
rect 6328 18312 11100 18340
rect 6328 18300 6334 18312
rect 2958 18272 2964 18284
rect 1780 18244 2964 18272
rect 1780 18213 1808 18244
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3050 18232 3056 18284
rect 3108 18272 3114 18284
rect 4709 18275 4767 18281
rect 4709 18272 4721 18275
rect 3108 18244 4721 18272
rect 3108 18232 3114 18244
rect 4709 18241 4721 18244
rect 4755 18241 4767 18275
rect 9398 18272 9404 18284
rect 9359 18244 9404 18272
rect 4709 18235 4767 18241
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 11072 18281 11100 18312
rect 11057 18275 11115 18281
rect 11057 18241 11069 18275
rect 11103 18241 11115 18275
rect 11057 18235 11115 18241
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 1765 18167 1823 18173
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2406 18164 2412 18216
rect 2464 18204 2470 18216
rect 6549 18207 6607 18213
rect 6549 18204 6561 18207
rect 2464 18176 6561 18204
rect 2464 18164 2470 18176
rect 6549 18173 6561 18176
rect 6595 18173 6607 18207
rect 6549 18167 6607 18173
rect 7101 18207 7159 18213
rect 7101 18173 7113 18207
rect 7147 18204 7159 18207
rect 7466 18204 7472 18216
rect 7147 18176 7472 18204
rect 7147 18173 7159 18176
rect 7101 18167 7159 18173
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18204 7803 18207
rect 9214 18204 9220 18216
rect 7791 18176 8340 18204
rect 9175 18176 9220 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 3418 18096 3424 18148
rect 3476 18136 3482 18148
rect 3476 18108 4108 18136
rect 3476 18096 3482 18108
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 1452 18040 1593 18068
rect 1452 18028 1458 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 2682 18028 2688 18080
rect 2740 18068 2746 18080
rect 2869 18071 2927 18077
rect 2869 18068 2881 18071
rect 2740 18040 2881 18068
rect 2740 18028 2746 18040
rect 2869 18037 2881 18040
rect 2915 18037 2927 18071
rect 3326 18068 3332 18080
rect 3287 18040 3332 18068
rect 2869 18031 2927 18037
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 3970 18068 3976 18080
rect 3931 18040 3976 18068
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 4080 18068 4108 18108
rect 4154 18096 4160 18148
rect 4212 18136 4218 18148
rect 5077 18139 5135 18145
rect 5077 18136 5089 18139
rect 4212 18108 5089 18136
rect 4212 18096 4218 18108
rect 5077 18105 5089 18108
rect 5123 18105 5135 18139
rect 5077 18099 5135 18105
rect 5626 18096 5632 18148
rect 5684 18136 5690 18148
rect 8021 18139 8079 18145
rect 8021 18136 8033 18139
rect 5684 18108 8033 18136
rect 5684 18096 5690 18108
rect 8021 18105 8033 18108
rect 8067 18105 8079 18139
rect 8021 18099 8079 18105
rect 8312 18080 8340 18176
rect 9214 18164 9220 18176
rect 9272 18204 9278 18216
rect 9858 18204 9864 18216
rect 9272 18176 9864 18204
rect 9272 18164 9278 18176
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 10919 18176 11744 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 11716 18080 11744 18176
rect 4341 18071 4399 18077
rect 4341 18068 4353 18071
rect 4080 18040 4353 18068
rect 4341 18037 4353 18040
rect 4387 18037 4399 18071
rect 4341 18031 4399 18037
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 6270 18068 6276 18080
rect 5951 18040 6276 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 7469 18071 7527 18077
rect 7469 18037 7481 18071
rect 7515 18068 7527 18071
rect 8202 18068 8208 18080
rect 7515 18040 8208 18068
rect 7515 18037 7527 18040
rect 7469 18031 7527 18037
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 8481 18071 8539 18077
rect 8481 18068 8493 18071
rect 8352 18040 8493 18068
rect 8352 18028 8358 18040
rect 8481 18037 8493 18040
rect 8527 18037 8539 18071
rect 8481 18031 8539 18037
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10229 18071 10287 18077
rect 10229 18068 10241 18071
rect 10192 18040 10241 18068
rect 10192 18028 10198 18040
rect 10229 18037 10241 18040
rect 10275 18037 10287 18071
rect 10229 18031 10287 18037
rect 10318 18028 10324 18080
rect 10376 18068 10382 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10376 18040 10609 18068
rect 10376 18028 10382 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 11698 18068 11704 18080
rect 11659 18040 11704 18068
rect 10597 18031 10655 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 2314 17824 2320 17876
rect 2372 17824 2378 17876
rect 2498 17824 2504 17876
rect 2556 17864 2562 17876
rect 6365 17867 6423 17873
rect 6365 17864 6377 17867
rect 2556 17836 6377 17864
rect 2556 17824 2562 17836
rect 6365 17833 6377 17836
rect 6411 17833 6423 17867
rect 9858 17864 9864 17876
rect 9819 17836 9864 17864
rect 6365 17827 6423 17833
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 2332 17796 2360 17824
rect 2593 17799 2651 17805
rect 2593 17796 2605 17799
rect 2332 17768 2605 17796
rect 2593 17765 2605 17768
rect 2639 17765 2651 17799
rect 2593 17759 2651 17765
rect 3878 17756 3884 17808
rect 3936 17796 3942 17808
rect 6733 17799 6791 17805
rect 6733 17796 6745 17799
rect 3936 17768 6745 17796
rect 3936 17756 3942 17768
rect 6733 17765 6745 17768
rect 6779 17765 6791 17799
rect 11790 17796 11796 17808
rect 6733 17759 6791 17765
rect 7852 17768 11796 17796
rect 1762 17728 1768 17740
rect 1723 17700 1768 17728
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 2314 17728 2320 17740
rect 2275 17700 2320 17728
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 2866 17688 2872 17740
rect 2924 17728 2930 17740
rect 5261 17731 5319 17737
rect 5261 17728 5273 17731
rect 2924 17700 5273 17728
rect 2924 17688 2930 17700
rect 5261 17697 5273 17700
rect 5307 17697 5319 17731
rect 5261 17691 5319 17697
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17660 5043 17663
rect 5534 17660 5540 17672
rect 5031 17632 5540 17660
rect 5031 17629 5043 17632
rect 4985 17623 5043 17629
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 2590 17552 2596 17604
rect 2648 17592 2654 17604
rect 3053 17595 3111 17601
rect 3053 17592 3065 17595
rect 2648 17564 3065 17592
rect 2648 17552 2654 17564
rect 3053 17561 3065 17564
rect 3099 17561 3111 17595
rect 3053 17555 3111 17561
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 7852 17601 7880 17768
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 10226 17728 10232 17740
rect 10187 17700 10232 17728
rect 10226 17688 10232 17700
rect 10284 17728 10290 17740
rect 10873 17731 10931 17737
rect 10873 17728 10885 17731
rect 10284 17700 10885 17728
rect 10284 17688 10290 17700
rect 10873 17697 10885 17700
rect 10919 17697 10931 17731
rect 10873 17691 10931 17697
rect 10318 17660 10324 17672
rect 10279 17632 10324 17660
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17660 10563 17663
rect 11146 17660 11152 17672
rect 10551 17632 11152 17660
rect 10551 17629 10563 17632
rect 10505 17623 10563 17629
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 13262 17660 13268 17672
rect 11348 17632 13268 17660
rect 5629 17595 5687 17601
rect 5629 17592 5641 17595
rect 3568 17564 5641 17592
rect 3568 17552 3574 17564
rect 5629 17561 5641 17564
rect 5675 17561 5687 17595
rect 7837 17595 7895 17601
rect 7837 17592 7849 17595
rect 5629 17555 5687 17561
rect 7484 17564 7849 17592
rect 7484 17536 7512 17564
rect 7837 17561 7849 17564
rect 7883 17561 7895 17595
rect 7837 17555 7895 17561
rect 8202 17552 8208 17604
rect 8260 17592 8266 17604
rect 8297 17595 8355 17601
rect 8297 17592 8309 17595
rect 8260 17564 8309 17592
rect 8260 17552 8266 17564
rect 8297 17561 8309 17564
rect 8343 17592 8355 17595
rect 9033 17595 9091 17601
rect 9033 17592 9045 17595
rect 8343 17564 9045 17592
rect 8343 17561 8355 17564
rect 8297 17555 8355 17561
rect 9033 17561 9045 17564
rect 9079 17592 9091 17595
rect 9122 17592 9128 17604
rect 9079 17564 9128 17592
rect 9079 17561 9091 17564
rect 9033 17555 9091 17561
rect 9122 17552 9128 17564
rect 9180 17592 9186 17604
rect 11348 17601 11376 17632
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 9180 17564 9413 17592
rect 9180 17552 9186 17564
rect 9401 17561 9413 17564
rect 9447 17592 9459 17595
rect 11333 17595 11391 17601
rect 11333 17592 11345 17595
rect 9447 17564 11345 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 11333 17561 11345 17564
rect 11379 17561 11391 17595
rect 11333 17555 11391 17561
rect 11793 17595 11851 17601
rect 11793 17561 11805 17595
rect 11839 17592 11851 17595
rect 12434 17592 12440 17604
rect 11839 17564 12440 17592
rect 11839 17561 11851 17564
rect 11793 17555 11851 17561
rect 12434 17552 12440 17564
rect 12492 17592 12498 17604
rect 13081 17595 13139 17601
rect 13081 17592 13093 17595
rect 12492 17564 13093 17592
rect 12492 17552 12498 17564
rect 13081 17561 13093 17564
rect 13127 17561 13139 17595
rect 13081 17555 13139 17561
rect 1673 17527 1731 17533
rect 1673 17493 1685 17527
rect 1719 17524 1731 17527
rect 2222 17524 2228 17536
rect 1719 17496 2228 17524
rect 1719 17493 1731 17496
rect 1673 17487 1731 17493
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 2682 17484 2688 17536
rect 2740 17524 2746 17536
rect 3421 17527 3479 17533
rect 3421 17524 3433 17527
rect 2740 17496 3433 17524
rect 2740 17484 2746 17496
rect 3421 17493 3433 17496
rect 3467 17493 3479 17527
rect 3421 17487 3479 17493
rect 3602 17484 3608 17536
rect 3660 17524 3666 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3660 17496 3801 17524
rect 3660 17484 3666 17496
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 3789 17487 3847 17493
rect 4617 17527 4675 17533
rect 4617 17493 4629 17527
rect 4663 17524 4675 17527
rect 4706 17524 4712 17536
rect 4663 17496 4712 17524
rect 4663 17493 4675 17496
rect 4617 17487 4675 17493
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 6086 17524 6092 17536
rect 6047 17496 6092 17524
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 6880 17496 7113 17524
rect 6880 17484 6886 17496
rect 7101 17493 7113 17496
rect 7147 17493 7159 17527
rect 7466 17524 7472 17536
rect 7427 17496 7472 17524
rect 7101 17487 7159 17493
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 8754 17524 8760 17536
rect 8715 17496 8760 17524
rect 8754 17484 8760 17496
rect 8812 17484 8818 17536
rect 12710 17524 12716 17536
rect 12671 17496 12716 17524
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1854 17320 1860 17332
rect 1815 17292 1860 17320
rect 1854 17280 1860 17292
rect 1912 17280 1918 17332
rect 2869 17323 2927 17329
rect 2869 17289 2881 17323
rect 2915 17320 2927 17323
rect 6454 17320 6460 17332
rect 2915 17292 6460 17320
rect 2915 17289 2927 17292
rect 2869 17283 2927 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17320 9919 17323
rect 10226 17320 10232 17332
rect 9907 17292 10232 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11333 17323 11391 17329
rect 11333 17320 11345 17323
rect 11204 17292 11345 17320
rect 11204 17280 11210 17292
rect 11333 17289 11345 17292
rect 11379 17320 11391 17323
rect 11606 17320 11612 17332
rect 11379 17292 11612 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 2314 17212 2320 17264
rect 2372 17252 2378 17264
rect 6549 17255 6607 17261
rect 2372 17224 4292 17252
rect 2372 17212 2378 17224
rect 1762 17144 1768 17196
rect 1820 17184 1826 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 1820 17156 2421 17184
rect 1820 17144 1826 17156
rect 2409 17153 2421 17156
rect 2455 17184 2467 17187
rect 4154 17184 4160 17196
rect 2455 17156 4160 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4264 17184 4292 17224
rect 6549 17221 6561 17255
rect 6595 17252 6607 17255
rect 6822 17252 6828 17264
rect 6595 17224 6828 17252
rect 6595 17221 6607 17224
rect 6549 17215 6607 17221
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 13814 17252 13820 17264
rect 13727 17224 13820 17252
rect 13814 17212 13820 17224
rect 13872 17252 13878 17264
rect 17954 17252 17960 17264
rect 13872 17224 17960 17252
rect 13872 17212 13878 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 6840 17184 6868 17212
rect 4264 17156 4384 17184
rect 6840 17156 6960 17184
rect 1670 17116 1676 17128
rect 1631 17088 1676 17116
rect 1670 17076 1676 17088
rect 1728 17116 1734 17128
rect 2038 17116 2044 17128
rect 1728 17088 2044 17116
rect 1728 17076 1734 17088
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17085 2283 17119
rect 2225 17079 2283 17085
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 2961 17119 3019 17125
rect 2961 17116 2973 17119
rect 2915 17088 2973 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 2961 17085 2973 17088
rect 3007 17085 3019 17119
rect 2961 17079 3019 17085
rect 2240 17048 2268 17079
rect 3142 17076 3148 17128
rect 3200 17116 3206 17128
rect 3237 17119 3295 17125
rect 3237 17116 3249 17119
rect 3200 17088 3249 17116
rect 3200 17076 3206 17088
rect 3237 17085 3249 17088
rect 3283 17085 3295 17119
rect 3237 17079 3295 17085
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4249 17119 4307 17125
rect 4249 17116 4261 17119
rect 4120 17088 4261 17116
rect 4120 17076 4126 17088
rect 4249 17085 4261 17088
rect 4295 17085 4307 17119
rect 4356 17116 4384 17156
rect 6270 17116 6276 17128
rect 4356 17088 6276 17116
rect 4249 17079 4307 17085
rect 6270 17076 6276 17088
rect 6328 17076 6334 17128
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6696 17088 6837 17116
rect 6696 17076 6702 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6932 17116 6960 17156
rect 7081 17119 7139 17125
rect 7081 17116 7093 17119
rect 6932 17088 7093 17116
rect 6825 17079 6883 17085
rect 7081 17085 7093 17088
rect 7127 17085 7139 17119
rect 7081 17079 7139 17085
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9732 17088 9965 17116
rect 9732 17076 9738 17088
rect 9953 17085 9965 17088
rect 9999 17085 10011 17119
rect 12434 17116 12440 17128
rect 12395 17088 12440 17116
rect 9953 17079 10011 17085
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 12710 17125 12716 17128
rect 12704 17116 12716 17125
rect 12671 17088 12716 17116
rect 12704 17079 12716 17088
rect 12710 17076 12716 17079
rect 12768 17076 12774 17128
rect 3694 17048 3700 17060
rect 2240 17020 3700 17048
rect 3694 17008 3700 17020
rect 3752 17008 3758 17060
rect 4154 17008 4160 17060
rect 4212 17048 4218 17060
rect 4494 17051 4552 17057
rect 4494 17048 4506 17051
rect 4212 17020 4506 17048
rect 4212 17008 4218 17020
rect 4494 17017 4506 17020
rect 4540 17048 4552 17051
rect 4706 17048 4712 17060
rect 4540 17020 4712 17048
rect 4540 17017 4552 17020
rect 4494 17011 4552 17017
rect 4706 17008 4712 17020
rect 4764 17008 4770 17060
rect 10134 17008 10140 17060
rect 10192 17057 10198 17060
rect 10192 17051 10256 17057
rect 10192 17017 10210 17051
rect 10244 17048 10256 17051
rect 11977 17051 12035 17057
rect 11977 17048 11989 17051
rect 10244 17020 11989 17048
rect 10244 17017 10256 17020
rect 10192 17011 10256 17017
rect 11977 17017 11989 17020
rect 12023 17017 12035 17051
rect 11977 17011 12035 17017
rect 10192 17008 10198 17011
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3510 16980 3516 16992
rect 3016 16952 3516 16980
rect 3016 16940 3022 16952
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 3786 16980 3792 16992
rect 3747 16952 3792 16980
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 5626 16980 5632 16992
rect 5587 16952 5632 16980
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 5994 16980 6000 16992
rect 5955 16952 6000 16980
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 8202 16980 8208 16992
rect 8163 16952 8208 16980
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 8570 16980 8576 16992
rect 8531 16952 8576 16980
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9493 16983 9551 16989
rect 9493 16980 9505 16983
rect 9171 16952 9505 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9493 16949 9505 16952
rect 9539 16980 9551 16983
rect 9582 16980 9588 16992
rect 9539 16952 9588 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2958 16776 2964 16788
rect 2332 16748 2964 16776
rect 2332 16649 2360 16748
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3234 16776 3240 16788
rect 3195 16748 3240 16776
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 3786 16776 3792 16788
rect 3747 16748 3792 16776
rect 3786 16736 3792 16748
rect 3844 16736 3850 16788
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 4764 16748 5457 16776
rect 4764 16736 4770 16748
rect 5445 16745 5457 16748
rect 5491 16745 5503 16779
rect 5445 16739 5503 16745
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 7101 16779 7159 16785
rect 7101 16776 7113 16779
rect 6880 16748 7113 16776
rect 6880 16736 6886 16748
rect 7101 16745 7113 16748
rect 7147 16745 7159 16779
rect 8294 16776 8300 16788
rect 8255 16748 8300 16776
rect 7101 16739 7159 16745
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 8754 16776 8760 16788
rect 8715 16748 8760 16776
rect 8754 16736 8760 16748
rect 8812 16776 8818 16788
rect 9766 16776 9772 16788
rect 8812 16748 9772 16776
rect 8812 16736 8818 16748
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 11054 16776 11060 16788
rect 10192 16748 11060 16776
rect 10192 16736 10198 16748
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11698 16736 11704 16788
rect 11756 16776 11762 16788
rect 12989 16779 13047 16785
rect 12989 16776 13001 16779
rect 11756 16748 13001 16776
rect 11756 16736 11762 16748
rect 12989 16745 13001 16748
rect 13035 16745 13047 16779
rect 12989 16739 13047 16745
rect 3418 16708 3424 16720
rect 2424 16680 3424 16708
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 2317 16643 2375 16649
rect 1811 16612 2268 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 2240 16572 2268 16612
rect 2317 16609 2329 16643
rect 2363 16609 2375 16643
rect 2317 16603 2375 16609
rect 2424 16572 2452 16680
rect 3418 16668 3424 16680
rect 3476 16668 3482 16720
rect 4080 16680 5120 16708
rect 4080 16652 4108 16680
rect 2593 16643 2651 16649
rect 2593 16609 2605 16643
rect 2639 16640 2651 16643
rect 3050 16640 3056 16652
rect 2639 16612 3056 16640
rect 2639 16609 2651 16612
rect 2593 16603 2651 16609
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 4062 16640 4068 16652
rect 4023 16612 4068 16640
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4321 16643 4379 16649
rect 4321 16640 4333 16643
rect 4172 16612 4333 16640
rect 2240 16544 2452 16572
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 4172 16572 4200 16612
rect 4321 16609 4333 16612
rect 4367 16640 4379 16643
rect 4890 16640 4896 16652
rect 4367 16612 4896 16640
rect 4367 16609 4379 16612
rect 4321 16603 4379 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 5092 16640 5120 16680
rect 5626 16668 5632 16720
rect 5684 16708 5690 16720
rect 5966 16711 6024 16717
rect 5966 16708 5978 16711
rect 5684 16680 5978 16708
rect 5684 16668 5690 16680
rect 5966 16677 5978 16680
rect 6012 16708 6024 16711
rect 7374 16708 7380 16720
rect 6012 16680 7380 16708
rect 6012 16677 6024 16680
rect 5966 16671 6024 16677
rect 7374 16668 7380 16680
rect 7432 16708 7438 16720
rect 7745 16711 7803 16717
rect 7745 16708 7757 16711
rect 7432 16680 7757 16708
rect 7432 16668 7438 16680
rect 7745 16677 7757 16680
rect 7791 16677 7803 16711
rect 7745 16671 7803 16677
rect 9122 16668 9128 16720
rect 9180 16708 9186 16720
rect 9674 16708 9680 16720
rect 9180 16680 9680 16708
rect 9180 16668 9186 16680
rect 9674 16668 9680 16680
rect 9732 16668 9738 16720
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 5092 16612 5733 16640
rect 5721 16609 5733 16612
rect 5767 16640 5779 16643
rect 7466 16640 7472 16652
rect 5767 16612 7472 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 7466 16600 7472 16612
rect 7524 16600 7530 16652
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8251 16612 8524 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 3016 16544 4200 16572
rect 8496 16572 8524 16612
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 8665 16643 8723 16649
rect 8665 16640 8677 16643
rect 8628 16612 8677 16640
rect 8628 16600 8634 16612
rect 8665 16609 8677 16612
rect 8711 16640 8723 16643
rect 9306 16640 9312 16652
rect 8711 16612 9312 16640
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 9950 16649 9956 16652
rect 9944 16640 9956 16649
rect 9911 16612 9956 16640
rect 9944 16603 9956 16612
rect 9950 16600 9956 16603
rect 10008 16600 10014 16652
rect 11606 16649 11612 16652
rect 11600 16640 11612 16649
rect 11567 16612 11612 16640
rect 11600 16603 11612 16612
rect 11606 16600 11612 16603
rect 11664 16600 11670 16652
rect 13354 16640 13360 16652
rect 13315 16612 13360 16640
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16640 13507 16643
rect 13722 16640 13728 16652
rect 13495 16612 13728 16640
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 8496 16544 8953 16572
rect 3016 16532 3022 16544
rect 8941 16541 8953 16544
rect 8987 16572 8999 16575
rect 8987 16544 9628 16572
rect 8987 16541 8999 16544
rect 8941 16535 8999 16541
rect 9398 16504 9404 16516
rect 6932 16476 9404 16504
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 6932 16436 6960 16476
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 7466 16436 7472 16448
rect 4856 16408 6960 16436
rect 7427 16408 7472 16436
rect 4856 16396 4862 16408
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 9600 16436 9628 16544
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 11333 16575 11391 16581
rect 9732 16544 9777 16572
rect 9732 16532 9738 16544
rect 11333 16541 11345 16575
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16572 13691 16575
rect 13814 16572 13820 16584
rect 13679 16544 13820 16572
rect 13679 16541 13691 16544
rect 13633 16535 13691 16541
rect 9950 16436 9956 16448
rect 9600 16408 9956 16436
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 11348 16436 11376 16535
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 12710 16504 12716 16516
rect 12671 16476 12716 16504
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 12434 16436 12440 16448
rect 11348 16408 12440 16436
rect 12434 16396 12440 16408
rect 12492 16436 12498 16448
rect 13078 16436 13084 16448
rect 12492 16408 13084 16436
rect 12492 16396 12498 16408
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1762 16232 1768 16244
rect 1723 16204 1768 16232
rect 1762 16192 1768 16204
rect 1820 16192 1826 16244
rect 2958 16232 2964 16244
rect 2919 16204 2964 16232
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3421 16235 3479 16241
rect 3421 16201 3433 16235
rect 3467 16232 3479 16235
rect 3510 16232 3516 16244
rect 3467 16204 3516 16232
rect 3467 16201 3479 16204
rect 3421 16195 3479 16201
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 4246 16232 4252 16244
rect 3620 16204 4252 16232
rect 2038 16056 2044 16108
rect 2096 16096 2102 16108
rect 2317 16099 2375 16105
rect 2317 16096 2329 16099
rect 2096 16068 2329 16096
rect 2096 16056 2102 16068
rect 2317 16065 2329 16068
rect 2363 16065 2375 16099
rect 3620 16096 3648 16204
rect 4246 16192 4252 16204
rect 4304 16232 4310 16244
rect 4433 16235 4491 16241
rect 4433 16232 4445 16235
rect 4304 16204 4445 16232
rect 4304 16192 4310 16204
rect 4433 16201 4445 16204
rect 4479 16201 4491 16235
rect 4433 16195 4491 16201
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6144 16204 6837 16232
rect 6144 16192 6150 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 9122 16232 9128 16244
rect 6825 16195 6883 16201
rect 8128 16204 9128 16232
rect 3694 16124 3700 16176
rect 3752 16164 3758 16176
rect 5629 16167 5687 16173
rect 5629 16164 5641 16167
rect 3752 16136 5641 16164
rect 3752 16124 3758 16136
rect 5629 16133 5641 16136
rect 5675 16133 5687 16167
rect 5629 16127 5687 16133
rect 3881 16099 3939 16105
rect 3881 16096 3893 16099
rect 3620 16068 3893 16096
rect 2317 16059 2375 16065
rect 3881 16065 3893 16068
rect 3927 16065 3939 16099
rect 3881 16059 3939 16065
rect 3973 16099 4031 16105
rect 3973 16065 3985 16099
rect 4019 16096 4031 16099
rect 4154 16096 4160 16108
rect 4019 16068 4160 16096
rect 4019 16065 4031 16068
rect 3973 16059 4031 16065
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 15997 1639 16031
rect 1581 15991 1639 15997
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 3786 16028 3792 16040
rect 2179 16000 2636 16028
rect 3747 16000 3792 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 1596 15960 1624 15991
rect 2314 15960 2320 15972
rect 1596 15932 2320 15960
rect 2314 15920 2320 15932
rect 2372 15920 2378 15972
rect 2608 15892 2636 16000
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 3329 15963 3387 15969
rect 3329 15929 3341 15963
rect 3375 15960 3387 15963
rect 3988 15960 4016 16059
rect 4154 16056 4160 16068
rect 4212 16056 4218 16108
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 4985 16099 5043 16105
rect 4985 16096 4997 16099
rect 4948 16068 4997 16096
rect 4948 16056 4954 16068
rect 4985 16065 4997 16068
rect 5031 16065 5043 16099
rect 6086 16096 6092 16108
rect 6047 16068 6092 16096
rect 4985 16059 5043 16065
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 6273 16099 6331 16105
rect 6273 16065 6285 16099
rect 6319 16096 6331 16099
rect 6822 16096 6828 16108
rect 6319 16068 6828 16096
rect 6319 16065 6331 16068
rect 6273 16059 6331 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 8128 16105 8156 16204
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 9766 16232 9772 16244
rect 9727 16204 9772 16232
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 10376 16204 10793 16232
rect 10376 16192 10382 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 10781 16195 10839 16201
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 12897 16235 12955 16241
rect 12897 16232 12909 16235
rect 11664 16204 12909 16232
rect 11664 16192 11670 16204
rect 12897 16201 12909 16204
rect 12943 16201 12955 16235
rect 12897 16195 12955 16201
rect 13449 16235 13507 16241
rect 13449 16201 13461 16235
rect 13495 16232 13507 16235
rect 13814 16232 13820 16244
rect 13495 16204 13820 16232
rect 13495 16201 13507 16204
rect 13449 16195 13507 16201
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 9493 16167 9551 16173
rect 9493 16133 9505 16167
rect 9539 16164 9551 16167
rect 9950 16164 9956 16176
rect 9539 16136 9956 16164
rect 9539 16133 9551 16136
rect 9493 16127 9551 16133
rect 9950 16124 9956 16136
rect 10008 16164 10014 16176
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 10008 16136 12173 16164
rect 10008 16124 10014 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12161 16127 12219 16133
rect 8113 16099 8171 16105
rect 8113 16065 8125 16099
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 9640 16068 10425 16096
rect 9640 16056 9646 16068
rect 10413 16065 10425 16068
rect 10459 16096 10471 16099
rect 10502 16096 10508 16108
rect 10459 16068 10508 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11333 16099 11391 16105
rect 11333 16096 11345 16099
rect 11112 16068 11345 16096
rect 11112 16056 11118 16068
rect 11333 16065 11345 16068
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16096 12495 16099
rect 13354 16096 13360 16108
rect 12483 16068 13360 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 13354 16056 13360 16068
rect 13412 16096 13418 16108
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13412 16068 13737 16096
rect 13412 16056 13418 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 5994 16028 6000 16040
rect 5955 16000 6000 16028
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 8380 16031 8438 16037
rect 8380 15997 8392 16031
rect 8426 16028 8438 16031
rect 9600 16028 9628 16056
rect 8426 16000 9628 16028
rect 8426 15997 8438 16000
rect 8380 15991 8438 15997
rect 3375 15932 4016 15960
rect 4893 15963 4951 15969
rect 3375 15929 3387 15932
rect 3329 15923 3387 15929
rect 4893 15929 4905 15963
rect 4939 15960 4951 15963
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 4939 15932 5549 15960
rect 4939 15929 4951 15932
rect 4893 15923 4951 15929
rect 5537 15929 5549 15932
rect 5583 15960 5595 15963
rect 5718 15960 5724 15972
rect 5583 15932 5724 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 5718 15920 5724 15932
rect 5776 15920 5782 15972
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 7466 15960 7472 15972
rect 7239 15932 7472 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 7466 15920 7472 15932
rect 7524 15960 7530 15972
rect 11146 15960 11152 15972
rect 7524 15932 11152 15960
rect 7524 15920 7530 15932
rect 11146 15920 11152 15932
rect 11204 15920 11210 15972
rect 4430 15892 4436 15904
rect 2608 15864 4436 15892
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7558 15892 7564 15904
rect 7331 15864 7564 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7558 15852 7564 15864
rect 7616 15892 7622 15904
rect 7837 15895 7895 15901
rect 7837 15892 7849 15895
rect 7616 15864 7849 15892
rect 7616 15852 7622 15864
rect 7837 15861 7849 15864
rect 7883 15861 7895 15895
rect 7837 15855 7895 15861
rect 9398 15852 9404 15904
rect 9456 15892 9462 15904
rect 10137 15895 10195 15901
rect 10137 15892 10149 15895
rect 9456 15864 10149 15892
rect 9456 15852 9462 15864
rect 10137 15861 10149 15864
rect 10183 15861 10195 15895
rect 10137 15855 10195 15861
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15892 10287 15895
rect 10686 15892 10692 15904
rect 10275 15864 10692 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 11241 15895 11299 15901
rect 11241 15861 11253 15895
rect 11287 15892 11299 15895
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11287 15864 11897 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 11885 15861 11897 15864
rect 11931 15892 11943 15895
rect 12342 15892 12348 15904
rect 11931 15864 12348 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14093 15895 14151 15901
rect 14093 15892 14105 15895
rect 13780 15864 14105 15892
rect 13780 15852 13786 15864
rect 14093 15861 14105 15864
rect 14139 15861 14151 15895
rect 14093 15855 14151 15861
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 3142 15688 3148 15700
rect 2056 15660 3148 15688
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 1578 15552 1584 15564
rect 1535 15524 1584 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 2056 15561 2084 15660
rect 3142 15648 3148 15660
rect 3200 15688 3206 15700
rect 3694 15688 3700 15700
rect 3200 15660 3700 15688
rect 3200 15648 3206 15660
rect 3694 15648 3700 15660
rect 3752 15648 3758 15700
rect 4890 15648 4896 15700
rect 4948 15688 4954 15700
rect 5442 15688 5448 15700
rect 4948 15660 5448 15688
rect 4948 15648 4954 15660
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5994 15688 6000 15700
rect 5955 15660 6000 15688
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 6104 15660 8309 15688
rect 2314 15620 2320 15632
rect 2275 15592 2320 15620
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 2866 15620 2872 15632
rect 2792 15592 2872 15620
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 2332 15484 2360 15580
rect 2792 15561 2820 15592
rect 2866 15580 2872 15592
rect 2924 15580 2930 15632
rect 3053 15623 3111 15629
rect 3053 15589 3065 15623
rect 3099 15620 3111 15623
rect 3418 15620 3424 15632
rect 3099 15592 3424 15620
rect 3099 15589 3111 15592
rect 3053 15583 3111 15589
rect 3418 15580 3424 15592
rect 3476 15580 3482 15632
rect 4246 15580 4252 15632
rect 4304 15629 4310 15632
rect 4304 15623 4368 15629
rect 4304 15589 4322 15623
rect 4356 15589 4368 15623
rect 4304 15583 4368 15589
rect 4304 15580 4310 15583
rect 4430 15580 4436 15632
rect 4488 15620 4494 15632
rect 4706 15620 4712 15632
rect 4488 15592 4712 15620
rect 4488 15580 4494 15592
rect 4706 15580 4712 15592
rect 4764 15620 4770 15632
rect 6104 15620 6132 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 9306 15688 9312 15700
rect 9267 15660 9312 15688
rect 8297 15651 8355 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 11146 15688 11152 15700
rect 11107 15660 11152 15688
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11517 15691 11575 15697
rect 11517 15657 11529 15691
rect 11563 15688 11575 15691
rect 13722 15688 13728 15700
rect 11563 15660 13728 15688
rect 11563 15657 11575 15660
rect 11517 15651 11575 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 4764 15592 6132 15620
rect 6181 15623 6239 15629
rect 4764 15580 4770 15592
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 8662 15620 8668 15632
rect 6227 15592 8668 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 8662 15580 8668 15592
rect 8720 15580 8726 15632
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15521 2835 15555
rect 3970 15552 3976 15564
rect 2777 15515 2835 15521
rect 2884 15524 3976 15552
rect 2884 15484 2912 15524
rect 3970 15512 3976 15524
rect 4028 15512 4034 15564
rect 6914 15561 6920 15564
rect 6908 15552 6920 15561
rect 6875 15524 6920 15552
rect 6908 15515 6920 15524
rect 6914 15512 6920 15515
rect 6972 15512 6978 15564
rect 8754 15552 8760 15564
rect 8715 15524 8760 15552
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 10042 15552 10048 15564
rect 10003 15524 10048 15552
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10410 15552 10416 15564
rect 10183 15524 10416 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10410 15512 10416 15524
rect 10468 15512 10474 15564
rect 11882 15552 11888 15564
rect 11843 15524 11888 15552
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 12621 15555 12679 15561
rect 12621 15521 12633 15555
rect 12667 15552 12679 15555
rect 12710 15552 12716 15564
rect 12667 15524 12716 15552
rect 12667 15521 12679 15524
rect 12621 15515 12679 15521
rect 4062 15484 4068 15496
rect 2332 15456 2912 15484
rect 4023 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 6638 15484 6644 15496
rect 6599 15456 6644 15484
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 8846 15484 8852 15496
rect 8807 15456 8852 15484
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 10008 15456 10241 15484
rect 10008 15444 10014 15456
rect 10229 15453 10241 15456
rect 10275 15484 10287 15487
rect 10962 15484 10968 15496
rect 10275 15456 10968 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11974 15484 11980 15496
rect 11935 15456 11980 15484
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15484 12219 15487
rect 12636 15484 12664 15515
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12207 15456 12664 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 8021 15419 8079 15425
rect 8021 15385 8033 15419
rect 8067 15416 8079 15419
rect 8864 15416 8892 15444
rect 8067 15388 8892 15416
rect 8067 15385 8079 15388
rect 8021 15379 8079 15385
rect 3510 15348 3516 15360
rect 3471 15320 3516 15348
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 4982 15308 4988 15360
rect 5040 15348 5046 15360
rect 9677 15351 9735 15357
rect 9677 15348 9689 15351
rect 5040 15320 9689 15348
rect 5040 15308 5046 15320
rect 9677 15317 9689 15320
rect 9723 15317 9735 15351
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 9677 15311 9735 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 12989 15351 13047 15357
rect 12989 15317 13001 15351
rect 13035 15348 13047 15351
rect 13078 15348 13084 15360
rect 13035 15320 13084 15348
rect 13035 15317 13047 15320
rect 12989 15311 13047 15317
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 1670 15144 1676 15156
rect 1631 15116 1676 15144
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 4062 15144 4068 15156
rect 2884 15116 4068 15144
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 2884 15017 2912 15116
rect 4062 15104 4068 15116
rect 4120 15144 4126 15156
rect 4706 15144 4712 15156
rect 4120 15116 4712 15144
rect 4120 15104 4126 15116
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 5500 15116 5549 15144
rect 5500 15104 5506 15116
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 5537 15107 5595 15113
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5684 15116 6009 15144
rect 5684 15104 5690 15116
rect 5997 15113 6009 15116
rect 6043 15113 6055 15147
rect 8662 15144 8668 15156
rect 8623 15116 8668 15144
rect 5997 15107 6055 15113
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 10502 15144 10508 15156
rect 8812 15116 10088 15144
rect 10463 15116 10508 15144
rect 8812 15104 8818 15116
rect 4246 15076 4252 15088
rect 4159 15048 4252 15076
rect 4246 15036 4252 15048
rect 4304 15076 4310 15088
rect 5169 15079 5227 15085
rect 5169 15076 5181 15079
rect 4304 15048 5181 15076
rect 4304 15036 4310 15048
rect 5169 15045 5181 15048
rect 5215 15045 5227 15079
rect 5169 15039 5227 15045
rect 7193 15079 7251 15085
rect 7193 15045 7205 15079
rect 7239 15076 7251 15079
rect 8772 15076 8800 15104
rect 7239 15048 8800 15076
rect 10060 15076 10088 15116
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 11882 15144 11888 15156
rect 10652 15116 11888 15144
rect 10652 15104 10658 15116
rect 11882 15104 11888 15116
rect 11940 15144 11946 15156
rect 12621 15147 12679 15153
rect 12621 15144 12633 15147
rect 11940 15116 12633 15144
rect 11940 15104 11946 15116
rect 12621 15113 12633 15116
rect 12667 15113 12679 15147
rect 12621 15107 12679 15113
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 13320 15116 13369 15144
rect 13320 15104 13326 15116
rect 13357 15113 13369 15116
rect 13403 15113 13415 15147
rect 13357 15107 13415 15113
rect 12989 15079 13047 15085
rect 12989 15076 13001 15079
rect 10060 15048 13001 15076
rect 7239 15045 7251 15048
rect 7193 15039 7251 15045
rect 12989 15045 13001 15048
rect 13035 15045 13047 15079
rect 12989 15039 13047 15045
rect 2225 15011 2283 15017
rect 2225 15008 2237 15011
rect 1636 14980 2237 15008
rect 1636 14968 1642 14980
rect 2225 14977 2237 14980
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 3970 14968 3976 15020
rect 4028 15008 4034 15020
rect 6641 15011 6699 15017
rect 4028 14980 6592 15008
rect 4028 14968 4034 14980
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14909 1547 14943
rect 1489 14903 1547 14909
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 3136 14943 3194 14949
rect 2087 14912 2452 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 1504 14872 1532 14903
rect 2424 14872 2452 14912
rect 3136 14909 3148 14943
rect 3182 14940 3194 14943
rect 3510 14940 3516 14952
rect 3182 14912 3516 14940
rect 3182 14909 3194 14912
rect 3136 14903 3194 14909
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 6564 14940 6592 14980
rect 6641 14977 6653 15011
rect 6687 15008 6699 15011
rect 6914 15008 6920 15020
rect 6687 14980 6920 15008
rect 6687 14977 6699 14980
rect 6641 14971 6699 14977
rect 6914 14968 6920 14980
rect 6972 15008 6978 15020
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 6972 14980 7849 15008
rect 6972 14968 6978 14980
rect 7837 14977 7849 14980
rect 7883 15008 7895 15011
rect 8202 15008 8208 15020
rect 7883 14980 8208 15008
rect 7883 14977 7895 14980
rect 7837 14971 7895 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 10502 15008 10508 15020
rect 10244 14980 10508 15008
rect 7009 14943 7067 14949
rect 7009 14940 7021 14943
rect 6564 14912 7021 14940
rect 7009 14909 7021 14912
rect 7055 14940 7067 14943
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7055 14912 7573 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 7561 14909 7573 14912
rect 7607 14909 7619 14943
rect 7561 14903 7619 14909
rect 5074 14872 5080 14884
rect 1504 14844 2176 14872
rect 2424 14844 5080 14872
rect 2148 14804 2176 14844
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 7576 14872 7604 14903
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 9122 14940 9128 14952
rect 8352 14912 9128 14940
rect 8352 14900 8358 14912
rect 9122 14900 9128 14912
rect 9180 14900 9186 14952
rect 9392 14943 9450 14949
rect 9392 14909 9404 14943
rect 9438 14940 9450 14943
rect 9950 14940 9956 14952
rect 9438 14912 9956 14940
rect 9438 14909 9450 14912
rect 9392 14903 9450 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 10244 14872 10272 14980
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 10962 14900 10968 14952
rect 11020 14940 11026 14952
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 11020 14912 11161 14940
rect 11020 14900 11026 14912
rect 11149 14909 11161 14912
rect 11195 14940 11207 14943
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11195 14912 11529 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 7576 14844 10272 14872
rect 2866 14804 2872 14816
rect 2148 14776 2872 14804
rect 2866 14764 2872 14776
rect 2924 14804 2930 14816
rect 3326 14804 3332 14816
rect 2924 14776 3332 14804
rect 2924 14764 2930 14776
rect 3326 14764 3332 14776
rect 3384 14764 3390 14816
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4856 14776 4905 14804
rect 4856 14764 4862 14776
rect 4893 14773 4905 14776
rect 4939 14804 4951 14807
rect 5350 14804 5356 14816
rect 4939 14776 5356 14804
rect 4939 14773 4951 14776
rect 4893 14767 4951 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 7650 14804 7656 14816
rect 7611 14776 7656 14804
rect 7650 14764 7656 14776
rect 7708 14804 7714 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 7708 14776 8217 14804
rect 7708 14764 7714 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 10594 14804 10600 14816
rect 8536 14776 10600 14804
rect 8536 14764 8542 14776
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11882 14804 11888 14816
rect 11843 14776 11888 14804
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 3142 14600 3148 14612
rect 3103 14572 3148 14600
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4246 14600 4252 14612
rect 3927 14572 4252 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5166 14600 5172 14612
rect 5040 14572 5172 14600
rect 5040 14560 5046 14572
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14569 6147 14603
rect 6089 14563 6147 14569
rect 2130 14532 2136 14544
rect 1688 14504 2136 14532
rect 1688 14473 1716 14504
rect 2130 14492 2136 14504
rect 2188 14492 2194 14544
rect 3510 14492 3516 14544
rect 3568 14532 3574 14544
rect 6104 14532 6132 14563
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 8260 14572 9045 14600
rect 8260 14560 8266 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9033 14563 9091 14569
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 10042 14600 10048 14612
rect 9723 14572 10048 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 10042 14560 10048 14572
rect 10100 14600 10106 14612
rect 10778 14600 10784 14612
rect 10100 14572 10784 14600
rect 10100 14560 10106 14572
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 11020 14572 11713 14600
rect 11020 14560 11026 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 11701 14563 11759 14569
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 13320 14572 13461 14600
rect 13320 14560 13326 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 13449 14563 13507 14569
rect 6362 14532 6368 14544
rect 3568 14504 6368 14532
rect 3568 14492 3574 14504
rect 6362 14492 6368 14504
rect 6420 14532 6426 14544
rect 6733 14535 6791 14541
rect 6733 14532 6745 14535
rect 6420 14504 6745 14532
rect 6420 14492 6426 14504
rect 6733 14501 6745 14504
rect 6779 14501 6791 14535
rect 6733 14495 6791 14501
rect 7276 14535 7334 14541
rect 7276 14501 7288 14535
rect 7322 14532 7334 14535
rect 8754 14532 8760 14544
rect 7322 14504 8760 14532
rect 7322 14501 7334 14504
rect 7276 14495 7334 14501
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 10410 14492 10416 14544
rect 10468 14532 10474 14544
rect 12713 14535 12771 14541
rect 12713 14532 12725 14535
rect 10468 14504 12725 14532
rect 10468 14492 10474 14504
rect 12713 14501 12725 14504
rect 12759 14501 12771 14535
rect 12713 14495 12771 14501
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14433 1731 14467
rect 2222 14464 2228 14476
rect 2135 14436 2228 14464
rect 1673 14427 1731 14433
rect 2222 14424 2228 14436
rect 2280 14464 2286 14476
rect 2406 14464 2412 14476
rect 2280 14436 2412 14464
rect 2280 14424 2286 14436
rect 2406 14424 2412 14436
rect 2464 14424 2470 14476
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14464 2559 14467
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2547 14436 2973 14464
rect 2547 14433 2559 14436
rect 2501 14427 2559 14433
rect 2961 14433 2973 14436
rect 3007 14464 3019 14467
rect 3786 14464 3792 14476
rect 3007 14436 3792 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 4965 14467 5023 14473
rect 4965 14464 4977 14467
rect 4632 14436 4977 14464
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 3936 14368 4077 14396
rect 3936 14356 3942 14368
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4632 14269 4660 14436
rect 4965 14433 4977 14436
rect 5011 14433 5023 14467
rect 4965 14427 5023 14433
rect 10588 14467 10646 14473
rect 10588 14433 10600 14467
rect 10634 14464 10646 14467
rect 11054 14464 11060 14476
rect 10634 14436 11060 14464
rect 10634 14433 10646 14436
rect 10588 14427 10646 14433
rect 11054 14424 11060 14436
rect 11112 14464 11118 14476
rect 11974 14464 11980 14476
rect 11112 14436 11980 14464
rect 11112 14424 11118 14436
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 4764 14368 4809 14396
rect 4764 14356 4770 14368
rect 6638 14356 6644 14408
rect 6696 14396 6702 14408
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6696 14368 7021 14396
rect 6696 14356 6702 14368
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 10318 14396 10324 14408
rect 10279 14368 10324 14396
rect 7009 14359 7067 14365
rect 4617 14263 4675 14269
rect 4617 14229 4629 14263
rect 4663 14260 4675 14263
rect 4706 14260 4712 14272
rect 4663 14232 4712 14260
rect 4663 14229 4675 14232
rect 4617 14223 4675 14229
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 6457 14263 6515 14269
rect 6457 14229 6469 14263
rect 6503 14260 6515 14263
rect 6638 14260 6644 14272
rect 6503 14232 6644 14260
rect 6503 14229 6515 14232
rect 6457 14223 6515 14229
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 7024 14260 7052 14359
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 11848 14368 13001 14396
rect 11848 14356 11854 14368
rect 12989 14365 13001 14368
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 9401 14331 9459 14337
rect 9401 14328 9413 14331
rect 8404 14300 9413 14328
rect 8404 14272 8432 14300
rect 9401 14297 9413 14300
rect 9447 14297 9459 14331
rect 9401 14291 9459 14297
rect 11330 14288 11336 14340
rect 11388 14328 11394 14340
rect 13817 14331 13875 14337
rect 13817 14328 13829 14331
rect 11388 14300 13829 14328
rect 11388 14288 11394 14300
rect 13817 14297 13829 14300
rect 13863 14328 13875 14331
rect 14458 14328 14464 14340
rect 13863 14300 14464 14328
rect 13863 14297 13875 14300
rect 13817 14291 13875 14297
rect 14458 14288 14464 14300
rect 14516 14288 14522 14340
rect 7374 14260 7380 14272
rect 7024 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8386 14260 8392 14272
rect 8347 14232 8392 14260
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 8754 14260 8760 14272
rect 8715 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 10134 14260 10140 14272
rect 10095 14232 10140 14260
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 12345 14263 12403 14269
rect 12345 14260 12357 14263
rect 10284 14232 12357 14260
rect 10284 14220 10290 14232
rect 12345 14229 12357 14232
rect 12391 14229 12403 14263
rect 12345 14223 12403 14229
rect 12989 14263 13047 14269
rect 12989 14229 13001 14263
rect 13035 14260 13047 14263
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 13035 14232 13185 14260
rect 13035 14229 13047 14232
rect 12989 14223 13047 14229
rect 13173 14229 13185 14232
rect 13219 14260 13231 14263
rect 13722 14260 13728 14272
rect 13219 14232 13728 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 3513 14059 3571 14065
rect 3513 14056 3525 14059
rect 3016 14028 3525 14056
rect 3016 14016 3022 14028
rect 3513 14025 3525 14028
rect 3559 14025 3571 14059
rect 3513 14019 3571 14025
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 6457 14059 6515 14065
rect 6457 14056 6469 14059
rect 4764 14028 6469 14056
rect 4764 14016 4770 14028
rect 6457 14025 6469 14028
rect 6503 14025 6515 14059
rect 6457 14019 6515 14025
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 7285 14059 7343 14065
rect 7285 14056 7297 14059
rect 6604 14028 7297 14056
rect 6604 14016 6610 14028
rect 7285 14025 7297 14028
rect 7331 14025 7343 14059
rect 7285 14019 7343 14025
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 8294 14056 8300 14068
rect 7432 14028 8300 14056
rect 7432 14016 7438 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8754 14056 8760 14068
rect 8715 14028 8760 14056
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 10413 14059 10471 14065
rect 8864 14028 10364 14056
rect 8864 13988 8892 14028
rect 7760 13960 8892 13988
rect 1946 13920 1952 13932
rect 1780 13892 1952 13920
rect 1780 13861 1808 13892
rect 1946 13880 1952 13892
rect 2004 13920 2010 13932
rect 2498 13920 2504 13932
rect 2004 13892 2504 13920
rect 2004 13880 2010 13892
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2866 13920 2872 13932
rect 2639 13892 2872 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 3602 13920 3608 13932
rect 3160 13892 3608 13920
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 3160 13852 3188 13892
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4246 13920 4252 13932
rect 4203 13892 4252 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4890 13880 4896 13932
rect 4948 13920 4954 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4948 13892 5089 13920
rect 4948 13880 4954 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 7282 13880 7288 13932
rect 7340 13920 7346 13932
rect 7760 13929 7788 13960
rect 8938 13948 8944 14000
rect 8996 13988 9002 14000
rect 9401 13991 9459 13997
rect 9401 13988 9413 13991
rect 8996 13960 9413 13988
rect 8996 13948 9002 13960
rect 9401 13957 9413 13960
rect 9447 13957 9459 13991
rect 9401 13951 9459 13957
rect 9490 13948 9496 14000
rect 9548 13988 9554 14000
rect 10226 13988 10232 14000
rect 9548 13960 9628 13988
rect 9548 13948 9554 13960
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7340 13892 7757 13920
rect 7340 13880 7346 13892
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13920 7987 13923
rect 8294 13920 8300 13932
rect 7975 13892 8300 13920
rect 7975 13889 7987 13892
rect 7929 13883 7987 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 8570 13880 8576 13932
rect 8628 13920 8634 13932
rect 8628 13892 9536 13920
rect 8628 13880 8634 13892
rect 2363 13824 3188 13852
rect 3421 13855 3479 13861
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2884 13796 2912 13824
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 3878 13852 3884 13864
rect 3467 13824 3884 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13852 4031 13855
rect 5344 13855 5402 13861
rect 4019 13824 5028 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 2866 13744 2872 13796
rect 2924 13744 2930 13796
rect 5000 13784 5028 13824
rect 5344 13821 5356 13855
rect 5390 13852 5402 13855
rect 6638 13852 6644 13864
rect 5390 13824 6644 13852
rect 5390 13821 5402 13824
rect 5344 13815 5402 13821
rect 6638 13812 6644 13824
rect 6696 13852 6702 13864
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 6696 13824 7021 13852
rect 6696 13812 6702 13824
rect 7009 13821 7021 13824
rect 7055 13821 7067 13855
rect 7009 13815 7067 13821
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 8478 13852 8484 13864
rect 7156 13824 8484 13852
rect 7156 13812 7162 13824
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 5534 13784 5540 13796
rect 5000 13756 5540 13784
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 8294 13744 8300 13796
rect 8352 13784 8358 13796
rect 9508 13784 9536 13892
rect 9600 13852 9628 13960
rect 9876 13960 10232 13988
rect 9876 13932 9904 13960
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 10336 13988 10364 14028
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 10502 14056 10508 14068
rect 10459 14028 10508 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 13262 14016 13268 14068
rect 13320 14056 13326 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13320 14028 14105 14056
rect 13320 14016 13326 14028
rect 14093 14025 14105 14028
rect 14139 14056 14151 14059
rect 14274 14056 14280 14068
rect 14139 14028 14280 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14458 14056 14464 14068
rect 14419 14028 14464 14056
rect 14458 14016 14464 14028
rect 14516 14056 14522 14068
rect 15470 14056 15476 14068
rect 14516 14028 15476 14056
rect 14516 14016 14522 14028
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 13354 13988 13360 14000
rect 10336 13960 11192 13988
rect 13315 13960 13360 13988
rect 9858 13920 9864 13932
rect 9771 13892 9864 13920
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 10042 13920 10048 13932
rect 10003 13892 10048 13920
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 11054 13920 11060 13932
rect 11015 13892 11060 13920
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 11164 13920 11192 13960
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 11164 13892 12633 13920
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 9769 13855 9827 13861
rect 9600 13824 9720 13852
rect 9692 13784 9720 13824
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10134 13852 10140 13864
rect 9815 13824 10140 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11532 13824 11805 13852
rect 9950 13784 9956 13796
rect 8352 13756 8708 13784
rect 9508 13756 9628 13784
rect 9692 13756 9956 13784
rect 8352 13744 8358 13756
rect 8680 13728 8708 13756
rect 1673 13719 1731 13725
rect 1673 13685 1685 13719
rect 1719 13716 1731 13719
rect 4062 13716 4068 13728
rect 1719 13688 4068 13716
rect 1719 13685 1731 13688
rect 1673 13679 1731 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4617 13719 4675 13725
rect 4617 13685 4629 13719
rect 4663 13716 4675 13719
rect 5166 13716 5172 13728
rect 4663 13688 5172 13716
rect 4663 13685 4675 13688
rect 4617 13679 4675 13685
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 7653 13719 7711 13725
rect 7653 13716 7665 13719
rect 6880 13688 7665 13716
rect 6880 13676 6886 13688
rect 7653 13685 7665 13688
rect 7699 13716 7711 13719
rect 8478 13716 8484 13728
rect 7699 13688 8484 13716
rect 7699 13685 7711 13688
rect 7653 13679 7711 13685
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 9125 13719 9183 13725
rect 9125 13716 9137 13719
rect 8720 13688 9137 13716
rect 8720 13676 8726 13688
rect 9125 13685 9137 13688
rect 9171 13685 9183 13719
rect 9600 13716 9628 13756
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10781 13787 10839 13793
rect 10781 13784 10793 13787
rect 10376 13756 10793 13784
rect 10376 13744 10382 13756
rect 10781 13753 10793 13756
rect 10827 13784 10839 13787
rect 11532 13784 11560 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 10827 13756 11560 13784
rect 10827 13753 10839 13756
rect 10781 13747 10839 13753
rect 11974 13744 11980 13796
rect 12032 13784 12038 13796
rect 12161 13787 12219 13793
rect 12161 13784 12173 13787
rect 12032 13756 12173 13784
rect 12032 13744 12038 13756
rect 12161 13753 12173 13756
rect 12207 13753 12219 13787
rect 12161 13747 12219 13753
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 13078 13784 13084 13796
rect 12492 13756 13084 13784
rect 12492 13744 12498 13756
rect 13078 13744 13084 13756
rect 13136 13784 13142 13796
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 13136 13756 14933 13784
rect 13136 13744 13142 13756
rect 14921 13753 14933 13756
rect 14967 13784 14979 13787
rect 16390 13784 16396 13796
rect 14967 13756 16396 13784
rect 14967 13753 14979 13756
rect 14921 13747 14979 13753
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 9766 13716 9772 13728
rect 9600 13688 9772 13716
rect 9125 13679 9183 13685
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10468 13688 10885 13716
rect 10468 13676 10474 13688
rect 10873 13685 10885 13688
rect 10919 13716 10931 13719
rect 11425 13719 11483 13725
rect 11425 13716 11437 13719
rect 10919 13688 11437 13716
rect 10919 13685 10931 13688
rect 10873 13679 10931 13685
rect 11425 13685 11437 13688
rect 11471 13685 11483 13719
rect 12986 13716 12992 13728
rect 12947 13688 12992 13716
rect 11425 13679 11483 13685
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 13780 13688 13829 13716
rect 13780 13676 13786 13688
rect 13817 13685 13829 13688
rect 13863 13716 13875 13719
rect 15194 13716 15200 13728
rect 13863 13688 15200 13716
rect 13863 13685 13875 13688
rect 13817 13679 13875 13685
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2593 13515 2651 13521
rect 2593 13481 2605 13515
rect 2639 13512 2651 13515
rect 2774 13512 2780 13524
rect 2639 13484 2780 13512
rect 2639 13481 2651 13484
rect 2593 13475 2651 13481
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 3694 13472 3700 13524
rect 3752 13512 3758 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 3752 13484 4813 13512
rect 3752 13472 3758 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 5166 13512 5172 13524
rect 5127 13484 5172 13512
rect 4801 13475 4859 13481
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5592 13484 5825 13512
rect 5592 13472 5598 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 5813 13475 5871 13481
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 8570 13512 8576 13524
rect 5960 13484 8576 13512
rect 5960 13472 5966 13484
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 9125 13515 9183 13521
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 10134 13512 10140 13524
rect 9171 13484 10140 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 11149 13515 11207 13521
rect 11149 13512 11161 13515
rect 11112 13484 11161 13512
rect 11112 13472 11118 13484
rect 11149 13481 11161 13484
rect 11195 13481 11207 13515
rect 12526 13512 12532 13524
rect 12487 13484 12532 13512
rect 11149 13475 11207 13481
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12894 13512 12900 13524
rect 12855 13484 12900 13512
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14332 13484 14749 13512
rect 14332 13472 14338 13484
rect 14737 13481 14749 13484
rect 14783 13512 14795 13515
rect 15286 13512 15292 13524
rect 14783 13484 15292 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 15470 13512 15476 13524
rect 15431 13484 15476 13512
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 1949 13447 2007 13453
rect 1949 13413 1961 13447
rect 1995 13444 2007 13447
rect 2130 13444 2136 13456
rect 1995 13416 2136 13444
rect 1995 13413 2007 13416
rect 1949 13407 2007 13413
rect 2130 13404 2136 13416
rect 2188 13404 2194 13456
rect 3142 13444 3148 13456
rect 2976 13416 3148 13444
rect 1670 13376 1676 13388
rect 1631 13348 1676 13376
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 2976 13385 3004 13416
rect 3142 13404 3148 13416
rect 3200 13444 3206 13456
rect 9398 13444 9404 13456
rect 3200 13416 9404 13444
rect 3200 13404 3206 13416
rect 9398 13404 9404 13416
rect 9456 13404 9462 13456
rect 10042 13453 10048 13456
rect 10036 13444 10048 13453
rect 10003 13416 10048 13444
rect 10036 13407 10048 13416
rect 10100 13444 10106 13456
rect 10962 13444 10968 13456
rect 10100 13416 10968 13444
rect 10042 13404 10048 13407
rect 10100 13404 10106 13416
rect 10962 13404 10968 13416
rect 11020 13444 11026 13456
rect 11425 13447 11483 13453
rect 11425 13444 11437 13447
rect 11020 13416 11437 13444
rect 11020 13404 11026 13416
rect 11425 13413 11437 13416
rect 11471 13444 11483 13447
rect 11793 13447 11851 13453
rect 11793 13444 11805 13447
rect 11471 13416 11805 13444
rect 11471 13413 11483 13416
rect 11425 13407 11483 13413
rect 11793 13413 11805 13416
rect 11839 13413 11851 13447
rect 11793 13407 11851 13413
rect 11974 13404 11980 13456
rect 12032 13444 12038 13456
rect 13265 13447 13323 13453
rect 13265 13444 13277 13447
rect 12032 13416 13277 13444
rect 12032 13404 12038 13416
rect 13265 13413 13277 13416
rect 13311 13413 13323 13447
rect 13265 13407 13323 13413
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13345 2467 13379
rect 2409 13339 2467 13345
rect 2961 13379 3019 13385
rect 2961 13345 2973 13379
rect 3007 13345 3019 13379
rect 2961 13339 3019 13345
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13376 3295 13379
rect 5902 13376 5908 13388
rect 3283 13348 5908 13376
rect 3283 13345 3295 13348
rect 3237 13339 3295 13345
rect 2424 13308 2452 13339
rect 3252 13308 3280 13339
rect 5902 13336 5908 13348
rect 5960 13336 5966 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 7006 13376 7012 13388
rect 6227 13348 7012 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7285 13379 7343 13385
rect 7285 13345 7297 13379
rect 7331 13376 7343 13379
rect 7374 13376 7380 13388
rect 7331 13348 7380 13376
rect 7331 13345 7343 13348
rect 7285 13339 7343 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7552 13379 7610 13385
rect 7552 13345 7564 13379
rect 7598 13376 7610 13379
rect 7598 13348 8432 13376
rect 7598 13345 7610 13348
rect 7552 13339 7610 13345
rect 2424 13280 3280 13308
rect 4706 13268 4712 13320
rect 4764 13268 4770 13320
rect 5258 13308 5264 13320
rect 5219 13280 5264 13308
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 4246 13200 4252 13252
rect 4304 13240 4310 13252
rect 4724 13240 4752 13268
rect 5368 13240 5396 13271
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 5868 13280 6285 13308
rect 5868 13268 5874 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 4304 13212 5396 13240
rect 6288 13240 6316 13271
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 6420 13280 6465 13308
rect 6420 13268 6426 13280
rect 8404 13252 8432 13348
rect 8478 13336 8484 13388
rect 8536 13376 8542 13388
rect 12986 13376 12992 13388
rect 8536 13348 12992 13376
rect 8536 13336 8542 13348
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 9766 13308 9772 13320
rect 9727 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 6825 13243 6883 13249
rect 6825 13240 6837 13243
rect 6288 13212 6837 13240
rect 4304 13200 4310 13212
rect 6825 13209 6837 13212
rect 6871 13209 6883 13243
rect 6825 13203 6883 13209
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 8444 13212 9076 13240
rect 8444 13200 8450 13212
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4154 13172 4160 13184
rect 3927 13144 4160 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 4341 13175 4399 13181
rect 4341 13141 4353 13175
rect 4387 13172 4399 13175
rect 4706 13172 4712 13184
rect 4387 13144 4712 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4798 13132 4804 13184
rect 4856 13172 4862 13184
rect 8478 13172 8484 13184
rect 4856 13144 8484 13172
rect 4856 13132 4862 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 8662 13172 8668 13184
rect 8623 13144 8668 13172
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 8938 13172 8944 13184
rect 8899 13144 8944 13172
rect 8938 13132 8944 13144
rect 8996 13132 9002 13184
rect 9048 13172 9076 13212
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 12161 13243 12219 13249
rect 12161 13240 12173 13243
rect 10836 13212 12173 13240
rect 10836 13200 10842 13212
rect 12161 13209 12173 13212
rect 12207 13209 12219 13243
rect 12161 13203 12219 13209
rect 12250 13200 12256 13252
rect 12308 13240 12314 13252
rect 13725 13243 13783 13249
rect 13725 13240 13737 13243
rect 12308 13212 13737 13240
rect 12308 13200 12314 13212
rect 13725 13209 13737 13212
rect 13771 13240 13783 13243
rect 17310 13240 17316 13252
rect 13771 13212 17316 13240
rect 13771 13209 13783 13212
rect 13725 13203 13783 13209
rect 17310 13200 17316 13212
rect 17368 13200 17374 13252
rect 11606 13172 11612 13184
rect 9048 13144 11612 13172
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 14093 13175 14151 13181
rect 14093 13141 14105 13175
rect 14139 13172 14151 13175
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14139 13144 14473 13172
rect 14139 13141 14151 13144
rect 14093 13135 14151 13141
rect 14461 13141 14473 13144
rect 14507 13172 14519 13175
rect 15194 13172 15200 13184
rect 14507 13144 15200 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 4246 12968 4252 12980
rect 2547 12940 4252 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4801 12971 4859 12977
rect 4801 12937 4813 12971
rect 4847 12968 4859 12971
rect 5166 12968 5172 12980
rect 4847 12940 5172 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5537 12971 5595 12977
rect 5537 12968 5549 12971
rect 5316 12940 5549 12968
rect 5316 12928 5322 12940
rect 5537 12937 5549 12940
rect 5583 12968 5595 12971
rect 5583 12940 10824 12968
rect 5583 12937 5595 12940
rect 5537 12931 5595 12937
rect 4525 12903 4583 12909
rect 4525 12869 4537 12903
rect 4571 12900 4583 12903
rect 4571 12872 8524 12900
rect 4571 12869 4583 12872
rect 4525 12863 4583 12869
rect 1688 12804 2728 12832
rect 1688 12773 1716 12804
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12733 1731 12767
rect 1946 12764 1952 12776
rect 1907 12736 1952 12764
rect 1673 12727 1731 12733
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 2498 12724 2504 12776
rect 2556 12764 2562 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2556 12736 2605 12764
rect 2556 12724 2562 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2700 12764 2728 12804
rect 3602 12792 3608 12844
rect 3660 12832 3666 12844
rect 6181 12835 6239 12841
rect 3660 12804 5580 12832
rect 3660 12792 3666 12804
rect 3878 12764 3884 12776
rect 2700 12736 3884 12764
rect 2593 12727 2651 12733
rect 3878 12724 3884 12736
rect 3936 12764 3942 12776
rect 4798 12764 4804 12776
rect 3936 12736 4804 12764
rect 3936 12724 3942 12736
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5552 12764 5580 12804
rect 6181 12801 6193 12835
rect 6227 12832 6239 12835
rect 6638 12832 6644 12844
rect 6227 12804 6644 12832
rect 6227 12801 6239 12804
rect 6181 12795 6239 12801
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 8386 12832 8392 12844
rect 7515 12804 8392 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 8496 12832 8524 12872
rect 8570 12860 8576 12912
rect 8628 12900 8634 12912
rect 9493 12903 9551 12909
rect 9493 12900 9505 12903
rect 8628 12872 9505 12900
rect 8628 12860 8634 12872
rect 9493 12869 9505 12872
rect 9539 12869 9551 12903
rect 10796 12900 10824 12940
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 11020 12940 11253 12968
rect 11020 12928 11026 12940
rect 11241 12937 11253 12940
rect 11287 12937 11299 12971
rect 11606 12968 11612 12980
rect 11519 12940 11612 12968
rect 11241 12931 11299 12937
rect 11606 12928 11612 12940
rect 11664 12968 11670 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11664 12940 11897 12968
rect 11664 12928 11670 12940
rect 11885 12937 11897 12940
rect 11931 12937 11943 12971
rect 11885 12931 11943 12937
rect 13446 12928 13452 12980
rect 13504 12968 13510 12980
rect 14461 12971 14519 12977
rect 14461 12968 14473 12971
rect 13504 12940 14473 12968
rect 13504 12928 13510 12940
rect 14461 12937 14473 12940
rect 14507 12937 14519 12971
rect 14461 12931 14519 12937
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 15344 12940 15577 12968
rect 15344 12928 15350 12940
rect 15565 12937 15577 12940
rect 15611 12968 15623 12971
rect 15933 12971 15991 12977
rect 15933 12968 15945 12971
rect 15611 12940 15945 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 15933 12937 15945 12940
rect 15979 12937 15991 12971
rect 15933 12931 15991 12937
rect 13357 12903 13415 12909
rect 13357 12900 13369 12903
rect 10796 12872 13369 12900
rect 9493 12863 9551 12869
rect 13357 12869 13369 12872
rect 13403 12869 13415 12903
rect 13357 12863 13415 12869
rect 8496 12804 9996 12832
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 5552 12736 7297 12764
rect 7285 12733 7297 12736
rect 7331 12764 7343 12767
rect 8202 12764 8208 12776
rect 7331 12736 8208 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 8478 12764 8484 12776
rect 8343 12736 8484 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 8478 12724 8484 12736
rect 8536 12764 8542 12776
rect 8938 12764 8944 12776
rect 8536 12736 8944 12764
rect 8536 12724 8542 12736
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 9861 12767 9919 12773
rect 9861 12764 9873 12767
rect 9824 12736 9873 12764
rect 9824 12724 9830 12736
rect 9861 12733 9873 12736
rect 9907 12733 9919 12767
rect 9968 12764 9996 12804
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 10928 12804 13737 12832
rect 10928 12792 10934 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 9968 12736 14105 12764
rect 9861 12727 9919 12733
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 2682 12656 2688 12708
rect 2740 12696 2746 12708
rect 2860 12699 2918 12705
rect 2860 12696 2872 12699
rect 2740 12668 2872 12696
rect 2740 12656 2746 12668
rect 2860 12665 2872 12668
rect 2906 12696 2918 12699
rect 3050 12696 3056 12708
rect 2906 12668 3056 12696
rect 2906 12665 2918 12668
rect 2860 12659 2918 12665
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 4525 12699 4583 12705
rect 4525 12696 4537 12699
rect 3528 12668 4537 12696
rect 1762 12588 1768 12640
rect 1820 12628 1826 12640
rect 3528 12628 3556 12668
rect 4525 12665 4537 12668
rect 4571 12665 4583 12699
rect 4525 12659 4583 12665
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5169 12699 5227 12705
rect 4948 12668 5120 12696
rect 4948 12656 4954 12668
rect 1820 12600 3556 12628
rect 1820 12588 1826 12600
rect 3602 12588 3608 12640
rect 3660 12628 3666 12640
rect 3973 12631 4031 12637
rect 3973 12628 3985 12631
rect 3660 12600 3985 12628
rect 3660 12588 3666 12600
rect 3973 12597 3985 12600
rect 4019 12597 4031 12631
rect 4246 12628 4252 12640
rect 4207 12600 4252 12628
rect 3973 12591 4031 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4430 12588 4436 12640
rect 4488 12628 4494 12640
rect 4982 12628 4988 12640
rect 4488 12600 4988 12628
rect 4488 12588 4494 12600
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5092 12628 5120 12668
rect 5169 12665 5181 12699
rect 5215 12696 5227 12699
rect 7193 12699 7251 12705
rect 5215 12668 5948 12696
rect 5215 12665 5227 12668
rect 5169 12659 5227 12665
rect 5920 12640 5948 12668
rect 7193 12665 7205 12699
rect 7239 12696 7251 12699
rect 8849 12699 8907 12705
rect 8849 12696 8861 12699
rect 7239 12668 8861 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 8849 12665 8861 12668
rect 8895 12696 8907 12699
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 8895 12668 9689 12696
rect 8895 12665 8907 12668
rect 8849 12659 8907 12665
rect 9677 12665 9689 12668
rect 9723 12665 9735 12699
rect 9677 12659 9735 12665
rect 10128 12699 10186 12705
rect 10128 12665 10140 12699
rect 10174 12696 10186 12699
rect 10502 12696 10508 12708
rect 10174 12668 10508 12696
rect 10174 12665 10186 12668
rect 10128 12659 10186 12665
rect 10502 12656 10508 12668
rect 10560 12656 10566 12708
rect 5258 12628 5264 12640
rect 5092 12600 5264 12628
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5902 12628 5908 12640
rect 5863 12600 5908 12628
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 5997 12631 6055 12637
rect 5997 12597 6009 12631
rect 6043 12628 6055 12631
rect 6086 12628 6092 12640
rect 6043 12600 6092 12628
rect 6043 12597 6055 12600
rect 5997 12591 6055 12597
rect 6086 12588 6092 12600
rect 6144 12628 6150 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6144 12600 6561 12628
rect 6144 12588 6150 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6549 12591 6607 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7837 12631 7895 12637
rect 7837 12628 7849 12631
rect 7340 12600 7849 12628
rect 7340 12588 7346 12600
rect 7837 12597 7849 12600
rect 7883 12597 7895 12631
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 7837 12591 7895 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 9306 12628 9312 12640
rect 8352 12600 9312 12628
rect 8352 12588 8358 12600
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9493 12631 9551 12637
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 11974 12628 11980 12640
rect 9539 12600 11980 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12618 12628 12624 12640
rect 12579 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 13081 12631 13139 12637
rect 13081 12597 13093 12631
rect 13127 12628 13139 12631
rect 13170 12628 13176 12640
rect 13127 12600 13176 12628
rect 13127 12597 13139 12600
rect 13081 12591 13139 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 14921 12631 14979 12637
rect 14921 12597 14933 12631
rect 14967 12628 14979 12631
rect 15194 12628 15200 12640
rect 14967 12600 15200 12628
rect 14967 12597 14979 12600
rect 14921 12591 14979 12597
rect 15194 12588 15200 12600
rect 15252 12628 15258 12640
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15252 12600 15301 12628
rect 15252 12588 15258 12600
rect 15289 12597 15301 12600
rect 15335 12628 15347 12631
rect 15838 12628 15844 12640
rect 15335 12600 15844 12628
rect 15335 12597 15347 12600
rect 15289 12591 15347 12597
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 16390 12628 16396 12640
rect 16303 12600 16396 12628
rect 16390 12588 16396 12600
rect 16448 12628 16454 12640
rect 17402 12628 17408 12640
rect 16448 12600 17408 12628
rect 16448 12588 16454 12600
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2222 12424 2228 12436
rect 1995 12396 2228 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2222 12384 2228 12396
rect 2280 12384 2286 12436
rect 3329 12427 3387 12433
rect 3329 12393 3341 12427
rect 3375 12424 3387 12427
rect 4246 12424 4252 12436
rect 3375 12396 4252 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4430 12424 4436 12436
rect 4391 12396 4436 12424
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 6638 12424 6644 12436
rect 4672 12396 5672 12424
rect 6599 12396 6644 12424
rect 4672 12384 4678 12396
rect 2409 12359 2467 12365
rect 2409 12325 2421 12359
rect 2455 12356 2467 12359
rect 3789 12359 3847 12365
rect 3789 12356 3801 12359
rect 2455 12328 3801 12356
rect 2455 12325 2467 12328
rect 2409 12319 2467 12325
rect 3789 12325 3801 12328
rect 3835 12325 3847 12359
rect 3789 12319 3847 12325
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 5442 12356 5448 12368
rect 4764 12328 5448 12356
rect 4764 12316 4770 12328
rect 5442 12316 5448 12328
rect 5500 12365 5506 12368
rect 5500 12359 5564 12365
rect 5500 12325 5518 12359
rect 5552 12325 5564 12359
rect 5644 12356 5672 12396
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 9677 12427 9735 12433
rect 6748 12396 8800 12424
rect 6748 12356 6776 12396
rect 7006 12356 7012 12368
rect 5644 12328 6776 12356
rect 6967 12328 7012 12356
rect 5500 12319 5564 12325
rect 5500 12316 5506 12319
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 7460 12359 7518 12365
rect 7460 12325 7472 12359
rect 7506 12356 7518 12359
rect 8662 12356 8668 12368
rect 7506 12328 8668 12356
rect 7506 12325 7518 12328
rect 7460 12319 7518 12325
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 8772 12356 8800 12396
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9858 12424 9864 12436
rect 9723 12396 9864 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10870 12424 10876 12436
rect 10100 12396 10876 12424
rect 10100 12384 10106 12396
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11425 12427 11483 12433
rect 11425 12424 11437 12427
rect 11112 12396 11437 12424
rect 11112 12384 11118 12396
rect 11425 12393 11437 12396
rect 11471 12393 11483 12427
rect 11425 12387 11483 12393
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12618 12424 12624 12436
rect 12575 12396 12624 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 12710 12384 12716 12436
rect 12768 12424 12774 12436
rect 15013 12427 15071 12433
rect 15013 12424 15025 12427
rect 12768 12396 15025 12424
rect 12768 12384 12774 12396
rect 15013 12393 15025 12396
rect 15059 12393 15071 12427
rect 15013 12387 15071 12393
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 16945 12427 17003 12433
rect 16945 12424 16957 12427
rect 15528 12396 16957 12424
rect 15528 12384 15534 12396
rect 16945 12393 16957 12396
rect 16991 12424 17003 12427
rect 20806 12424 20812 12436
rect 16991 12396 20812 12424
rect 16991 12393 17003 12396
rect 16945 12387 17003 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 9950 12356 9956 12368
rect 8772 12328 9956 12356
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 10137 12359 10195 12365
rect 10137 12325 10149 12359
rect 10183 12325 10195 12359
rect 10137 12319 10195 12325
rect 1394 12288 1400 12300
rect 1307 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12288 1458 12300
rect 1946 12288 1952 12300
rect 1452 12260 1952 12288
rect 1452 12248 1458 12260
rect 1946 12248 1952 12260
rect 2004 12248 2010 12300
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 3602 12288 3608 12300
rect 2363 12260 2544 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2516 12152 2544 12260
rect 2608 12260 3608 12288
rect 2608 12229 2636 12260
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 4890 12288 4896 12300
rect 4571 12260 4896 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12288 5043 12291
rect 8294 12288 8300 12300
rect 5031 12260 8300 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 9858 12288 9864 12300
rect 8864 12260 9864 12288
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 3418 12220 3424 12232
rect 3379 12192 3424 12220
rect 2593 12183 2651 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3510 12180 3516 12232
rect 3568 12220 3574 12232
rect 4614 12220 4620 12232
rect 3568 12192 4620 12220
rect 3568 12180 3574 12192
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 4764 12192 5212 12220
rect 4764 12180 4770 12192
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2516 12124 2973 12152
rect 2961 12121 2973 12124
rect 3007 12152 3019 12155
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 3007 12124 4997 12152
rect 3007 12121 3019 12124
rect 2961 12115 3019 12121
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 5184 12152 5212 12192
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 5316 12192 5361 12220
rect 5316 12180 5322 12192
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6880 12192 7205 12220
rect 6880 12180 6886 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 8864 12229 8892 12260
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 10152 12288 10180 12319
rect 10226 12316 10232 12368
rect 10284 12356 10290 12368
rect 12805 12359 12863 12365
rect 12805 12356 12817 12359
rect 10284 12328 12817 12356
rect 10284 12316 10290 12328
rect 12805 12325 12817 12328
rect 12851 12325 12863 12359
rect 12805 12319 12863 12325
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 10152 12260 10701 12288
rect 10152 12232 10180 12260
rect 10689 12257 10701 12260
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 11146 12248 11152 12300
rect 11204 12288 11210 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11204 12260 12173 12288
rect 11204 12248 11210 12260
rect 12161 12257 12173 12260
rect 12207 12288 12219 12291
rect 15562 12288 15568 12300
rect 12207 12260 15568 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 8849 12223 8907 12229
rect 8849 12220 8861 12223
rect 8260 12192 8861 12220
rect 8260 12180 8266 12192
rect 8849 12189 8861 12192
rect 8895 12189 8907 12223
rect 8849 12183 8907 12189
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 10042 12220 10048 12232
rect 9180 12192 10048 12220
rect 9180 12180 9186 12192
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10134 12180 10140 12232
rect 10192 12180 10198 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10502 12220 10508 12232
rect 10367 12192 10508 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10502 12180 10508 12192
rect 10560 12220 10566 12232
rect 11698 12220 11704 12232
rect 10560 12192 11704 12220
rect 10560 12180 10566 12192
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 12860 12192 13185 12220
rect 12860 12180 12866 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 11606 12152 11612 12164
rect 5184 12124 5304 12152
rect 4985 12115 5043 12121
rect 3050 12044 3056 12096
rect 3108 12084 3114 12096
rect 3510 12084 3516 12096
rect 3108 12056 3516 12084
rect 3108 12044 3114 12056
rect 3510 12044 3516 12056
rect 3568 12044 3574 12096
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3835 12056 4077 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 4065 12053 4077 12056
rect 4111 12084 4123 12087
rect 4706 12084 4712 12096
rect 4111 12056 4712 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4948 12056 5089 12084
rect 4948 12044 4954 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5276 12084 5304 12124
rect 6196 12124 7052 12152
rect 6196 12084 6224 12124
rect 5276 12056 6224 12084
rect 7024 12084 7052 12124
rect 8128 12124 11612 12152
rect 8128 12084 8156 12124
rect 11606 12112 11612 12124
rect 11664 12112 11670 12164
rect 11885 12155 11943 12161
rect 11885 12121 11897 12155
rect 11931 12152 11943 12155
rect 12066 12152 12072 12164
rect 11931 12124 12072 12152
rect 11931 12121 11943 12124
rect 11885 12115 11943 12121
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 13909 12155 13967 12161
rect 13909 12152 13921 12155
rect 12912 12124 13921 12152
rect 7024 12056 8156 12084
rect 5077 12047 5135 12053
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8260 12056 8585 12084
rect 8260 12044 8266 12056
rect 8573 12053 8585 12056
rect 8619 12053 8631 12087
rect 9398 12084 9404 12096
rect 9359 12056 9404 12084
rect 8573 12047 8631 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 10962 12084 10968 12096
rect 9824 12056 10968 12084
rect 9824 12044 9830 12056
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11112 12056 11157 12084
rect 11112 12044 11118 12056
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11848 12056 11989 12084
rect 11848 12044 11854 12056
rect 11977 12053 11989 12056
rect 12023 12084 12035 12087
rect 12434 12084 12440 12096
rect 12023 12056 12440 12084
rect 12023 12053 12035 12056
rect 11977 12047 12035 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12912 12084 12940 12124
rect 13909 12121 13921 12124
rect 13955 12121 13967 12155
rect 14274 12152 14280 12164
rect 14235 12124 14280 12152
rect 13909 12115 13967 12121
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 15838 12112 15844 12164
rect 15896 12152 15902 12164
rect 15933 12155 15991 12161
rect 15933 12152 15945 12155
rect 15896 12124 15945 12152
rect 15896 12112 15902 12124
rect 15933 12121 15945 12124
rect 15979 12152 15991 12155
rect 16482 12152 16488 12164
rect 15979 12124 16488 12152
rect 15979 12121 15991 12124
rect 15933 12115 15991 12121
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 19058 12152 19064 12164
rect 19019 12124 19064 12152
rect 19058 12112 19064 12124
rect 19116 12112 19122 12164
rect 13538 12084 13544 12096
rect 12584 12056 12940 12084
rect 13499 12056 13544 12084
rect 12584 12044 12590 12056
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 13872 12056 14657 12084
rect 13872 12044 13878 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 15436 12056 15485 12084
rect 15436 12044 15442 12056
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 15473 12047 15531 12053
rect 16301 12087 16359 12093
rect 16301 12053 16313 12087
rect 16347 12084 16359 12087
rect 16390 12084 16396 12096
rect 16347 12056 16396 12084
rect 16347 12053 16359 12056
rect 16301 12047 16359 12053
rect 16390 12044 16396 12056
rect 16448 12084 16454 12096
rect 16577 12087 16635 12093
rect 16577 12084 16589 12087
rect 16448 12056 16589 12084
rect 16448 12044 16454 12056
rect 16577 12053 16589 12056
rect 16623 12053 16635 12087
rect 17402 12084 17408 12096
rect 17363 12056 17408 12084
rect 16577 12047 16635 12053
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1762 11880 1768 11892
rect 1723 11852 1768 11880
rect 1762 11840 1768 11852
rect 1820 11840 1826 11892
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 4246 11880 4252 11892
rect 2915 11852 4252 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5500 11852 6469 11880
rect 5500 11840 5506 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 7098 11880 7104 11892
rect 7059 11852 7104 11880
rect 6457 11843 6515 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 7892 11852 8585 11880
rect 7892 11840 7898 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 9030 11880 9036 11892
rect 8991 11852 9036 11880
rect 8573 11843 8631 11849
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 10226 11880 10232 11892
rect 9508 11852 10232 11880
rect 6270 11772 6276 11824
rect 6328 11812 6334 11824
rect 7377 11815 7435 11821
rect 7377 11812 7389 11815
rect 6328 11784 7389 11812
rect 6328 11772 6334 11784
rect 7377 11781 7389 11784
rect 7423 11781 7435 11815
rect 7377 11775 7435 11781
rect 2314 11744 2320 11756
rect 2275 11716 2320 11744
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 9122 11744 9128 11756
rect 8067 11716 9128 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9508 11753 9536 11852
rect 10226 11840 10232 11852
rect 10284 11880 10290 11892
rect 13538 11880 13544 11892
rect 10284 11852 11100 11880
rect 10284 11840 10290 11852
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 9953 11815 10011 11821
rect 9953 11812 9965 11815
rect 9824 11784 9965 11812
rect 9824 11772 9830 11784
rect 9953 11781 9965 11784
rect 9999 11781 10011 11815
rect 9953 11775 10011 11781
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 11072 11744 11100 11852
rect 11256 11852 13544 11880
rect 11256 11824 11284 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 15562 11880 15568 11892
rect 15523 11852 15568 11880
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 11238 11772 11244 11824
rect 11296 11772 11302 11824
rect 11425 11815 11483 11821
rect 11425 11781 11437 11815
rect 11471 11812 11483 11815
rect 11698 11812 11704 11824
rect 11471 11784 11704 11812
rect 11471 11781 11483 11784
rect 11425 11775 11483 11781
rect 11698 11772 11704 11784
rect 11756 11812 11762 11824
rect 12618 11812 12624 11824
rect 11756 11784 12624 11812
rect 11756 11772 11762 11784
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 9723 11716 10180 11744
rect 11072 11716 14473 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2958 11676 2964 11688
rect 2179 11648 2964 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3292 11648 3341 11676
rect 3292 11636 3298 11648
rect 3329 11645 3341 11648
rect 3375 11676 3387 11679
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 3375 11648 5089 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 5077 11645 5089 11648
rect 5123 11676 5135 11679
rect 5166 11676 5172 11688
rect 5123 11648 5172 11676
rect 5123 11645 5135 11648
rect 5077 11639 5135 11645
rect 5166 11636 5172 11648
rect 5224 11676 5230 11688
rect 6822 11676 6828 11688
rect 5224 11648 6828 11676
rect 5224 11636 5230 11648
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7282 11676 7288 11688
rect 7243 11648 7288 11676
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 9861 11679 9919 11685
rect 9861 11676 9873 11679
rect 7984 11648 9873 11676
rect 7984 11636 7990 11648
rect 9861 11645 9873 11648
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 9999 11648 10057 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10045 11645 10057 11648
rect 10091 11645 10103 11679
rect 10152 11676 10180 11716
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 10312 11679 10370 11685
rect 10312 11676 10324 11679
rect 10152 11648 10324 11676
rect 10045 11639 10103 11645
rect 10312 11645 10324 11648
rect 10358 11676 10370 11679
rect 11054 11676 11060 11688
rect 10358 11648 11060 11676
rect 10358 11645 10370 11648
rect 10312 11639 10370 11645
rect 11054 11636 11060 11648
rect 11112 11676 11118 11688
rect 12066 11676 12072 11688
rect 11112 11648 12072 11676
rect 11112 11636 11118 11648
rect 12066 11636 12072 11648
rect 12124 11676 12130 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12124 11648 12633 11676
rect 12124 11636 12130 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 13780 11648 15209 11676
rect 13780 11636 13786 11648
rect 15197 11645 15209 11648
rect 15243 11645 15255 11679
rect 19058 11676 19064 11688
rect 19019 11648 19064 11676
rect 15197 11639 15255 11645
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 19610 11676 19616 11688
rect 19571 11648 19616 11676
rect 19610 11636 19616 11648
rect 19668 11676 19674 11688
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 19668 11648 20177 11676
rect 19668 11636 19674 11648
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 3602 11617 3608 11620
rect 1673 11611 1731 11617
rect 1673 11577 1685 11611
rect 1719 11608 1731 11611
rect 3596 11608 3608 11617
rect 1719 11580 3608 11608
rect 1719 11577 1731 11580
rect 1673 11571 1731 11577
rect 3596 11571 3608 11580
rect 3602 11568 3608 11571
rect 3660 11568 3666 11620
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 4246 11608 4252 11620
rect 4120 11580 4252 11608
rect 4120 11568 4126 11580
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 5350 11617 5356 11620
rect 5344 11608 5356 11617
rect 5311 11580 5356 11608
rect 5344 11571 5356 11580
rect 5350 11568 5356 11571
rect 5408 11568 5414 11620
rect 7834 11608 7840 11620
rect 7795 11580 7840 11608
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 8386 11608 8392 11620
rect 8036 11580 8392 11608
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 2188 11512 2237 11540
rect 2188 11500 2194 11512
rect 2225 11509 2237 11512
rect 2271 11540 2283 11543
rect 2406 11540 2412 11552
rect 2271 11512 2412 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3237 11543 3295 11549
rect 3237 11540 3249 11543
rect 2832 11512 3249 11540
rect 2832 11500 2838 11512
rect 3237 11509 3249 11512
rect 3283 11540 3295 11543
rect 3418 11540 3424 11552
rect 3283 11512 3424 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 7745 11543 7803 11549
rect 7745 11509 7757 11543
rect 7791 11540 7803 11543
rect 8036 11540 8064 11580
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 8573 11611 8631 11617
rect 8573 11577 8585 11611
rect 8619 11608 8631 11611
rect 12342 11608 12348 11620
rect 8619 11580 12348 11608
rect 8619 11577 8631 11580
rect 8573 11571 8631 11577
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 13630 11568 13636 11620
rect 13688 11608 13694 11620
rect 14829 11611 14887 11617
rect 14829 11608 14841 11611
rect 13688 11580 14841 11608
rect 13688 11568 13694 11580
rect 14829 11577 14841 11580
rect 14875 11577 14887 11611
rect 14829 11571 14887 11577
rect 15378 11568 15384 11620
rect 15436 11608 15442 11620
rect 16301 11611 16359 11617
rect 16301 11608 16313 11611
rect 15436 11580 16313 11608
rect 15436 11568 15442 11580
rect 16301 11577 16313 11580
rect 16347 11577 16359 11611
rect 16301 11571 16359 11577
rect 16390 11568 16396 11620
rect 16448 11608 16454 11620
rect 17037 11611 17095 11617
rect 17037 11608 17049 11611
rect 16448 11580 17049 11608
rect 16448 11568 16454 11580
rect 17037 11577 17049 11580
rect 17083 11608 17095 11611
rect 17405 11611 17463 11617
rect 17405 11608 17417 11611
rect 17083 11580 17417 11608
rect 17083 11577 17095 11580
rect 17037 11571 17095 11577
rect 17405 11577 17417 11580
rect 17451 11608 17463 11611
rect 17773 11611 17831 11617
rect 17773 11608 17785 11611
rect 17451 11580 17785 11608
rect 17451 11577 17463 11580
rect 17405 11571 17463 11577
rect 17773 11577 17785 11580
rect 17819 11577 17831 11611
rect 17773 11571 17831 11577
rect 7791 11512 8064 11540
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 9398 11540 9404 11552
rect 8812 11512 8857 11540
rect 9359 11512 9404 11540
rect 8812 11500 8818 11512
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10778 11540 10784 11552
rect 9907 11512 10784 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 10928 11512 11713 11540
rect 10928 11500 10934 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 12066 11540 12072 11552
rect 12027 11512 12072 11540
rect 11701 11503 11759 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13446 11540 13452 11552
rect 13407 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13722 11540 13728 11552
rect 13683 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 14090 11540 14096 11552
rect 14051 11512 14096 11540
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15933 11543 15991 11549
rect 15933 11540 15945 11543
rect 15252 11512 15945 11540
rect 15252 11500 15258 11512
rect 15933 11509 15945 11512
rect 15979 11540 15991 11543
rect 16206 11540 16212 11552
rect 15979 11512 16212 11540
rect 15979 11509 15991 11512
rect 15933 11503 15991 11509
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16482 11500 16488 11552
rect 16540 11540 16546 11552
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16540 11512 16681 11540
rect 16540 11500 16546 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 19242 11540 19248 11552
rect 19203 11512 19248 11540
rect 16669 11503 16727 11509
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 20346 11540 20352 11552
rect 19843 11512 20352 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2498 11296 2504 11348
rect 2556 11296 2562 11348
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3145 11339 3203 11345
rect 3145 11336 3157 11339
rect 3108 11308 3157 11336
rect 3108 11296 3114 11308
rect 3145 11305 3157 11308
rect 3191 11305 3203 11339
rect 3145 11299 3203 11305
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 4801 11339 4859 11345
rect 4801 11336 4813 11339
rect 3660 11308 4813 11336
rect 3660 11296 3666 11308
rect 4801 11305 4813 11308
rect 4847 11305 4859 11339
rect 4801 11299 4859 11305
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5132 11308 5181 11336
rect 5132 11296 5138 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 5169 11299 5227 11305
rect 6733 11339 6791 11345
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 7006 11336 7012 11348
rect 6779 11308 7012 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 7006 11296 7012 11308
rect 7064 11336 7070 11348
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 7064 11308 7113 11336
rect 7064 11296 7070 11308
rect 7101 11305 7113 11308
rect 7147 11336 7159 11339
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 7147 11308 9229 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 9456 11308 11345 11336
rect 9456 11296 9462 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12124 11308 12909 11336
rect 12124 11296 12130 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 15620 11308 16221 11336
rect 15620 11296 15626 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16209 11299 16267 11305
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 16540 11308 17325 11336
rect 16540 11296 16546 11308
rect 17313 11305 17325 11308
rect 17359 11305 17371 11339
rect 17313 11299 17371 11305
rect 2032 11271 2090 11277
rect 2032 11237 2044 11271
rect 2078 11268 2090 11271
rect 2314 11268 2320 11280
rect 2078 11240 2320 11268
rect 2078 11237 2090 11240
rect 2032 11231 2090 11237
rect 2314 11228 2320 11240
rect 2372 11228 2378 11280
rect 2516 11200 2544 11296
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 5350 11268 5356 11280
rect 4212 11240 5356 11268
rect 4212 11228 4218 11240
rect 5350 11228 5356 11240
rect 5408 11228 5414 11280
rect 5626 11268 5632 11280
rect 5539 11240 5632 11268
rect 5626 11228 5632 11240
rect 5684 11268 5690 11280
rect 6822 11268 6828 11280
rect 5684 11240 6828 11268
rect 5684 11228 5690 11240
rect 6822 11228 6828 11240
rect 6880 11228 6886 11280
rect 7469 11271 7527 11277
rect 7469 11237 7481 11271
rect 7515 11268 7527 11271
rect 8110 11268 8116 11280
rect 7515 11240 8116 11268
rect 7515 11237 7527 11240
rect 7469 11231 7527 11237
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 9674 11268 9680 11280
rect 9180 11240 9680 11268
rect 9180 11228 9186 11240
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 9950 11277 9956 11280
rect 9944 11268 9956 11277
rect 9911 11240 9956 11268
rect 9944 11231 9956 11240
rect 9950 11228 9956 11231
rect 10008 11228 10014 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 12268 11240 13645 11268
rect 3234 11200 3240 11212
rect 1780 11172 3240 11200
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 1780 11141 1808 11172
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 3605 11203 3663 11209
rect 3605 11169 3617 11203
rect 3651 11200 3663 11203
rect 3786 11200 3792 11212
rect 3651 11172 3792 11200
rect 3651 11169 3663 11172
rect 3605 11163 3663 11169
rect 3786 11160 3792 11172
rect 3844 11160 3850 11212
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4172 11172 4537 11200
rect 4172 11144 4200 11172
rect 4525 11169 4537 11172
rect 4571 11200 4583 11203
rect 4982 11200 4988 11212
rect 4571 11172 4988 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 5537 11203 5595 11209
rect 5537 11169 5549 11203
rect 5583 11200 5595 11203
rect 5583 11172 6224 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 6196 11144 6224 11172
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7432 11172 7573 11200
rect 7432 11160 7438 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 7828 11203 7886 11209
rect 7828 11169 7840 11203
rect 7874 11200 7886 11203
rect 8202 11200 8208 11212
rect 7874 11172 8208 11200
rect 7874 11169 7886 11172
rect 7828 11163 7886 11169
rect 8202 11160 8208 11172
rect 8260 11200 8266 11212
rect 8260 11172 10732 11200
rect 8260 11160 8266 11172
rect 1765 11135 1823 11141
rect 1765 11132 1777 11135
rect 1544 11104 1777 11132
rect 1544 11092 1550 11104
rect 1765 11101 1777 11104
rect 1811 11101 1823 11135
rect 1765 11095 1823 11101
rect 4154 11092 4160 11144
rect 4212 11092 4218 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 6178 11132 6184 11144
rect 6139 11104 6184 11132
rect 5721 11095 5779 11101
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 5736 11064 5764 11095
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 9122 11132 9128 11144
rect 8956 11104 9128 11132
rect 8956 11073 8984 11104
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 10704 11132 10732 11172
rect 10778 11160 10784 11212
rect 10836 11200 10842 11212
rect 12268 11200 12296 11240
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 10836 11172 12296 11200
rect 10836 11160 10842 11172
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 13722 11200 13728 11212
rect 12400 11172 13728 11200
rect 12400 11160 12406 11172
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 15436 11172 16589 11200
rect 15436 11160 15442 11172
rect 16577 11169 16589 11172
rect 16623 11200 16635 11203
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 16623 11172 16957 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 16945 11169 16957 11172
rect 16991 11200 17003 11203
rect 17586 11200 17592 11212
rect 16991 11172 17592 11200
rect 16991 11169 17003 11172
rect 16945 11163 17003 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 18506 11200 18512 11212
rect 18467 11172 18512 11200
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 10704 11104 13400 11132
rect 13372 11076 13400 11104
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 13964 11104 14749 11132
rect 13964 11092 13970 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 16390 11132 16396 11144
rect 15344 11104 16396 11132
rect 15344 11092 15350 11104
rect 16390 11092 16396 11104
rect 16448 11132 16454 11144
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 16448 11104 18061 11132
rect 16448 11092 16454 11104
rect 18049 11101 18061 11104
rect 18095 11132 18107 11135
rect 19426 11132 19432 11144
rect 18095 11104 19432 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 5500 11036 5764 11064
rect 8941 11067 8999 11073
rect 5500 11024 5506 11036
rect 8941 11033 8953 11067
rect 8987 11033 8999 11067
rect 11054 11064 11060 11076
rect 11015 11036 11060 11064
rect 8941 11027 8999 11033
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11885 11067 11943 11073
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 12434 11064 12440 11076
rect 11931 11036 12440 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 13354 11064 13360 11076
rect 13315 11036 13360 11064
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 14366 11064 14372 11076
rect 14327 11036 14372 11064
rect 14366 11024 14372 11036
rect 14424 11024 14430 11076
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 16022 11064 16028 11076
rect 15979 11036 16028 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 16022 11024 16028 11036
rect 16080 11024 16086 11076
rect 16574 11024 16580 11076
rect 16632 11064 16638 11076
rect 17681 11067 17739 11073
rect 17681 11064 17693 11067
rect 16632 11036 17693 11064
rect 16632 11024 16638 11036
rect 17681 11033 17693 11036
rect 17727 11064 17739 11067
rect 18598 11064 18604 11076
rect 17727 11036 18604 11064
rect 17727 11033 17739 11036
rect 17681 11027 17739 11033
rect 18598 11024 18604 11036
rect 18656 11024 18662 11076
rect 18693 11067 18751 11073
rect 18693 11033 18705 11067
rect 18739 11064 18751 11067
rect 19058 11064 19064 11076
rect 18739 11036 19064 11064
rect 18739 11033 18751 11036
rect 18693 11027 18751 11033
rect 19058 11024 19064 11036
rect 19116 11024 19122 11076
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 1762 10996 1768 11008
rect 1719 10968 1768 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 1762 10956 1768 10968
rect 1820 10956 1826 11008
rect 1946 10956 1952 11008
rect 2004 10996 2010 11008
rect 3050 10996 3056 11008
rect 2004 10968 3056 10996
rect 2004 10956 2010 10968
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 9582 10996 9588 11008
rect 3752 10968 9588 10996
rect 3752 10956 3758 10968
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10778 10996 10784 11008
rect 9732 10968 10784 10996
rect 9732 10956 9738 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 12253 10999 12311 11005
rect 12253 10965 12265 10999
rect 12299 10996 12311 10999
rect 12621 10999 12679 11005
rect 12621 10996 12633 10999
rect 12299 10968 12633 10996
rect 12299 10965 12311 10968
rect 12253 10959 12311 10965
rect 12621 10965 12633 10968
rect 12667 10996 12679 10999
rect 13538 10996 13544 11008
rect 12667 10968 13544 10996
rect 12667 10965 12679 10968
rect 12621 10959 12679 10965
rect 13538 10956 13544 10968
rect 13596 10956 13602 11008
rect 13998 10996 14004 11008
rect 13959 10968 14004 10996
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 15565 10999 15623 11005
rect 15565 10965 15577 10999
rect 15611 10996 15623 10999
rect 15654 10996 15660 11008
rect 15611 10968 15660 10996
rect 15611 10965 15623 10968
rect 15565 10959 15623 10965
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2869 10795 2927 10801
rect 2869 10792 2881 10795
rect 2464 10764 2881 10792
rect 2464 10752 2470 10764
rect 2869 10761 2881 10764
rect 2915 10761 2927 10795
rect 2869 10755 2927 10761
rect 3234 10752 3240 10804
rect 3292 10792 3298 10804
rect 3292 10764 4752 10792
rect 3292 10752 3298 10764
rect 2958 10684 2964 10736
rect 3016 10724 3022 10736
rect 3145 10727 3203 10733
rect 3145 10724 3157 10727
rect 3016 10696 3157 10724
rect 3016 10684 3022 10696
rect 3145 10693 3157 10696
rect 3191 10724 3203 10727
rect 3191 10696 4660 10724
rect 3191 10693 3203 10696
rect 3145 10687 3203 10693
rect 1486 10656 1492 10668
rect 1447 10628 1492 10656
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 2648 10628 3709 10656
rect 2648 10616 2654 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 1756 10591 1814 10597
rect 1756 10557 1768 10591
rect 1802 10588 1814 10591
rect 2608 10588 2636 10616
rect 1802 10560 2636 10588
rect 1802 10557 1814 10560
rect 1756 10551 1814 10557
rect 2866 10548 2872 10600
rect 2924 10588 2930 10600
rect 3970 10588 3976 10600
rect 2924 10560 3976 10588
rect 2924 10548 2930 10560
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4632 10588 4660 10696
rect 4724 10665 4752 10764
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6236 10764 6377 10792
rect 6236 10752 6242 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 7742 10792 7748 10804
rect 7607 10764 7748 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 8389 10795 8447 10801
rect 8389 10761 8401 10795
rect 8435 10792 8447 10795
rect 10226 10792 10232 10804
rect 8435 10764 9628 10792
rect 10187 10764 10232 10792
rect 8435 10761 8447 10764
rect 8389 10755 8447 10761
rect 8294 10724 8300 10736
rect 7116 10696 8300 10724
rect 7116 10665 7144 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 8202 10656 8208 10668
rect 8163 10628 8208 10656
rect 7101 10619 7159 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 4632 10560 8401 10588
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8527 10560 8585 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8840 10591 8898 10597
rect 8840 10557 8852 10591
rect 8886 10588 8898 10591
rect 9122 10588 9128 10600
rect 8886 10560 9128 10588
rect 8886 10557 8898 10560
rect 8840 10551 8898 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9600 10588 9628 10764
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 13354 10752 13360 10804
rect 13412 10792 13418 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13412 10764 13921 10792
rect 13412 10752 13418 10764
rect 13909 10761 13921 10764
rect 13955 10761 13967 10795
rect 13909 10755 13967 10761
rect 16206 10752 16212 10804
rect 16264 10792 16270 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 16264 10764 17233 10792
rect 16264 10752 16270 10764
rect 17221 10761 17233 10764
rect 17267 10761 17279 10795
rect 17221 10755 17279 10761
rect 9950 10724 9956 10736
rect 9863 10696 9956 10724
rect 9950 10684 9956 10696
rect 10008 10724 10014 10736
rect 13078 10724 13084 10736
rect 10008 10696 13084 10724
rect 10008 10684 10014 10696
rect 10888 10665 10916 10696
rect 13078 10684 13084 10696
rect 13136 10724 13142 10736
rect 14277 10727 14335 10733
rect 14277 10724 14289 10727
rect 13136 10696 14289 10724
rect 13136 10684 13142 10696
rect 14277 10693 14289 10696
rect 14323 10693 14335 10727
rect 14277 10687 14335 10693
rect 14458 10684 14464 10736
rect 14516 10724 14522 10736
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 14516 10696 15025 10724
rect 14516 10684 14522 10696
rect 15013 10693 15025 10696
rect 15059 10693 15071 10727
rect 17236 10724 17264 10755
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 17460 10764 19809 10792
rect 17460 10752 17466 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 17954 10724 17960 10736
rect 17236 10696 17960 10724
rect 15013 10687 15071 10693
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18506 10684 18512 10736
rect 18564 10724 18570 10736
rect 19061 10727 19119 10733
rect 19061 10724 19073 10727
rect 18564 10696 19073 10724
rect 18564 10684 18570 10696
rect 19061 10693 19073 10696
rect 19107 10693 19119 10727
rect 19426 10724 19432 10736
rect 19387 10696 19432 10724
rect 19061 10687 19119 10693
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 14182 10616 14188 10668
rect 14240 10656 14246 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 14240 10628 15761 10656
rect 14240 10616 14246 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 17586 10656 17592 10668
rect 17547 10628 17592 10656
rect 15749 10619 15807 10625
rect 17586 10616 17592 10628
rect 17644 10616 17650 10668
rect 10502 10588 10508 10600
rect 9600 10560 10508 10588
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10594 10548 10600 10600
rect 10652 10548 10658 10600
rect 11425 10591 11483 10597
rect 11425 10557 11437 10591
rect 11471 10588 11483 10591
rect 11606 10588 11612 10600
rect 11471 10560 11612 10588
rect 11471 10557 11483 10560
rect 11425 10551 11483 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 13998 10588 14004 10600
rect 11900 10560 14004 10588
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 3786 10520 3792 10532
rect 3651 10492 3792 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 3786 10480 3792 10492
rect 3844 10480 3850 10532
rect 4982 10529 4988 10532
rect 4976 10520 4988 10529
rect 4943 10492 4988 10520
rect 4976 10483 4988 10492
rect 4982 10480 4988 10483
rect 5040 10480 5046 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 5408 10492 6132 10520
rect 5408 10480 5414 10492
rect 3510 10452 3516 10464
rect 3471 10424 3516 10452
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 4249 10455 4307 10461
rect 4249 10421 4261 10455
rect 4295 10452 4307 10455
rect 5994 10452 6000 10464
rect 4295 10424 6000 10452
rect 4295 10421 4307 10424
rect 4249 10415 4307 10421
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6104 10461 6132 10492
rect 7466 10480 7472 10532
rect 7524 10520 7530 10532
rect 10042 10520 10048 10532
rect 7524 10492 10048 10520
rect 7524 10480 7530 10492
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 6089 10455 6147 10461
rect 6089 10421 6101 10455
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7800 10424 7941 10452
rect 7800 10412 7806 10424
rect 7929 10421 7941 10424
rect 7975 10421 7987 10455
rect 7929 10415 7987 10421
rect 8021 10455 8079 10461
rect 8021 10421 8033 10455
rect 8067 10452 8079 10455
rect 8202 10452 8208 10464
rect 8067 10424 8208 10452
rect 8067 10421 8079 10424
rect 8021 10415 8079 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 9122 10452 9128 10464
rect 8527 10424 9128 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 9674 10452 9680 10464
rect 9548 10424 9680 10452
rect 9548 10412 9554 10424
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 10612 10461 10640 10548
rect 10689 10523 10747 10529
rect 10689 10489 10701 10523
rect 10735 10520 10747 10523
rect 10778 10520 10784 10532
rect 10735 10492 10784 10520
rect 10735 10489 10747 10492
rect 10689 10483 10747 10489
rect 10778 10480 10784 10492
rect 10836 10520 10842 10532
rect 11701 10523 11759 10529
rect 11701 10520 11713 10523
rect 10836 10492 11713 10520
rect 10836 10480 10842 10492
rect 11701 10489 11713 10492
rect 11747 10489 11759 10523
rect 11701 10483 11759 10489
rect 10597 10455 10655 10461
rect 10597 10421 10609 10455
rect 10643 10421 10655 10455
rect 11238 10452 11244 10464
rect 11199 10424 11244 10452
rect 10597 10415 10655 10421
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11330 10412 11336 10464
rect 11388 10452 11394 10464
rect 11900 10452 11928 10560
rect 13998 10548 14004 10560
rect 14056 10588 14062 10600
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14056 10560 14657 10588
rect 14056 10548 14062 10560
rect 14645 10557 14657 10560
rect 14691 10588 14703 10591
rect 15010 10588 15016 10600
rect 14691 10560 15016 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 18138 10588 18144 10600
rect 18099 10560 18144 10588
rect 18138 10548 18144 10560
rect 18196 10588 18202 10600
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18196 10560 18705 10588
rect 18196 10548 18202 10560
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 16117 10523 16175 10529
rect 16117 10520 16129 10523
rect 12676 10492 16129 10520
rect 12676 10480 12682 10492
rect 16117 10489 16129 10492
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 12066 10452 12072 10464
rect 11388 10424 11928 10452
rect 12027 10424 12072 10452
rect 11388 10412 11394 10424
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 12986 10452 12992 10464
rect 12943 10424 12992 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13262 10452 13268 10464
rect 13223 10424 13268 10452
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 13538 10452 13544 10464
rect 13499 10424 13544 10452
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 15381 10455 15439 10461
rect 15381 10452 15393 10455
rect 13780 10424 15393 10452
rect 13780 10412 13786 10424
rect 15381 10421 15393 10424
rect 15427 10421 15439 10455
rect 15381 10415 15439 10421
rect 16577 10455 16635 10461
rect 16577 10421 16589 10455
rect 16623 10452 16635 10455
rect 16666 10452 16672 10464
rect 16623 10424 16672 10452
rect 16623 10421 16635 10424
rect 16577 10415 16635 10421
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16942 10452 16948 10464
rect 16903 10424 16948 10452
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 18325 10455 18383 10461
rect 18325 10421 18337 10455
rect 18371 10452 18383 10455
rect 18966 10452 18972 10464
rect 18371 10424 18972 10452
rect 18371 10421 18383 10424
rect 18325 10415 18383 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 2130 10248 2136 10260
rect 2091 10220 2136 10248
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3510 10248 3516 10260
rect 3191 10220 3516 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3510 10208 3516 10220
rect 3568 10248 3574 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 3568 10220 3617 10248
rect 3568 10208 3574 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 3605 10211 3663 10217
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 5721 10251 5779 10257
rect 5721 10248 5733 10251
rect 4028 10220 5733 10248
rect 4028 10208 4034 10220
rect 5721 10217 5733 10220
rect 5767 10217 5779 10251
rect 5721 10211 5779 10217
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 6052 10220 6101 10248
rect 6052 10208 6058 10220
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 6089 10211 6147 10217
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 7340 10220 8493 10248
rect 7340 10208 7346 10220
rect 8481 10217 8493 10220
rect 8527 10248 8539 10251
rect 8570 10248 8576 10260
rect 8527 10220 8576 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 11790 10248 11796 10260
rect 8680 10220 11796 10248
rect 3050 10140 3056 10192
rect 3108 10180 3114 10192
rect 7009 10183 7067 10189
rect 7009 10180 7021 10183
rect 3108 10152 7021 10180
rect 3108 10140 3114 10152
rect 7009 10149 7021 10152
rect 7055 10149 7067 10183
rect 7009 10143 7067 10149
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2041 10115 2099 10121
rect 2041 10112 2053 10115
rect 1719 10084 2053 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2041 10081 2053 10084
rect 2087 10112 2099 10115
rect 4332 10115 4390 10121
rect 4332 10112 4344 10115
rect 2087 10084 4344 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 4332 10081 4344 10084
rect 4378 10112 4390 10115
rect 4706 10112 4712 10124
rect 4378 10084 4712 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 5592 10084 6193 10112
rect 5592 10072 5598 10084
rect 6181 10081 6193 10084
rect 6227 10112 6239 10115
rect 6733 10115 6791 10121
rect 6227 10084 6408 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 2682 10004 2688 10056
rect 2740 10044 2746 10056
rect 3510 10044 3516 10056
rect 2740 10016 3516 10044
rect 2740 10004 2746 10016
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3752 10016 4077 10044
rect 3752 10004 3758 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6288 9976 6316 10007
rect 5460 9948 6316 9976
rect 6380 9976 6408 10084
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 7190 10112 7196 10124
rect 6779 10084 7196 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 8680 10121 8708 10220
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13044 10220 13553 10248
rect 13044 10208 13050 10220
rect 13541 10217 13553 10220
rect 13587 10248 13599 10251
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 13587 10220 13829 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 13817 10211 13875 10217
rect 14001 10251 14059 10257
rect 14001 10217 14013 10251
rect 14047 10248 14059 10251
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14047 10220 14749 10248
rect 14047 10217 14059 10220
rect 14001 10211 14059 10217
rect 14737 10217 14749 10220
rect 14783 10217 14795 10251
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 14737 10211 14795 10217
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 17310 10248 17316 10260
rect 17271 10220 17316 10248
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17773 10251 17831 10257
rect 17773 10217 17785 10251
rect 17819 10248 17831 10251
rect 17954 10248 17960 10260
rect 17819 10220 17960 10248
rect 17819 10217 17831 10220
rect 17773 10211 17831 10217
rect 17954 10208 17960 10220
rect 18012 10248 18018 10260
rect 18049 10251 18107 10257
rect 18049 10248 18061 10251
rect 18012 10220 18061 10248
rect 18012 10208 18018 10220
rect 18049 10217 18061 10220
rect 18095 10217 18107 10251
rect 18049 10211 18107 10217
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 18656 10220 19165 10248
rect 18656 10208 18662 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 19153 10211 19211 10217
rect 19426 10208 19432 10260
rect 19484 10248 19490 10260
rect 19521 10251 19579 10257
rect 19521 10248 19533 10251
rect 19484 10220 19533 10248
rect 19484 10208 19490 10220
rect 19521 10217 19533 10220
rect 19567 10248 19579 10251
rect 19889 10251 19947 10257
rect 19889 10248 19901 10251
rect 19567 10220 19901 10248
rect 19567 10217 19579 10220
rect 19521 10211 19579 10217
rect 19889 10217 19901 10220
rect 19935 10248 19947 10251
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 19935 10220 20269 10248
rect 19935 10217 19947 10220
rect 19889 10211 19947 10217
rect 20257 10217 20269 10220
rect 20303 10248 20315 10251
rect 20438 10248 20444 10260
rect 20303 10220 20444 10248
rect 20303 10217 20315 10220
rect 20257 10211 20315 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 16945 10183 17003 10189
rect 16945 10180 16957 10183
rect 8956 10152 16957 10180
rect 8665 10115 8723 10121
rect 8665 10081 8677 10115
rect 8711 10081 8723 10115
rect 8665 10075 8723 10081
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8846 10044 8852 10056
rect 8067 10016 8852 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 8956 9976 8984 10152
rect 16945 10149 16957 10152
rect 16991 10149 17003 10183
rect 16945 10143 17003 10149
rect 17586 10140 17592 10192
rect 17644 10180 17650 10192
rect 17862 10180 17868 10192
rect 17644 10152 17868 10180
rect 17644 10140 17650 10152
rect 17862 10140 17868 10152
rect 17920 10180 17926 10192
rect 18417 10183 18475 10189
rect 18417 10180 18429 10183
rect 17920 10152 18429 10180
rect 17920 10140 17926 10152
rect 18417 10149 18429 10152
rect 18463 10180 18475 10183
rect 18785 10183 18843 10189
rect 18785 10180 18797 10183
rect 18463 10152 18797 10180
rect 18463 10149 18475 10152
rect 18417 10143 18475 10149
rect 18785 10149 18797 10152
rect 18831 10149 18843 10183
rect 18785 10143 18843 10149
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 10962 10112 10968 10124
rect 10367 10084 10968 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 9324 10044 9352 10075
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 11882 10072 11888 10124
rect 11940 10112 11946 10124
rect 12434 10121 12440 10124
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 11940 10084 12173 10112
rect 11940 10072 11946 10084
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 12428 10075 12440 10121
rect 12492 10112 12498 10124
rect 13262 10112 13268 10124
rect 12492 10084 13268 10112
rect 12434 10072 12440 10075
rect 12492 10072 12498 10084
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 11238 10044 11244 10056
rect 9324 10016 11244 10044
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 13722 10044 13728 10056
rect 13188 10016 13728 10044
rect 6380 9948 8984 9976
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 4982 9908 4988 9920
rect 1820 9880 4988 9908
rect 1820 9868 1826 9880
rect 4982 9868 4988 9880
rect 5040 9908 5046 9920
rect 5460 9917 5488 9948
rect 9030 9936 9036 9988
rect 9088 9976 9094 9988
rect 12066 9976 12072 9988
rect 9088 9948 12072 9976
rect 9088 9936 9094 9948
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 5040 9880 5457 9908
rect 5040 9868 5046 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 5445 9871 5503 9877
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 7469 9911 7527 9917
rect 7469 9908 7481 9911
rect 6144 9880 7481 9908
rect 6144 9868 6150 9880
rect 7469 9877 7481 9880
rect 7515 9877 7527 9911
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7469 9871 7527 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8720 9880 8953 9908
rect 8720 9868 8726 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 9122 9908 9128 9920
rect 9035 9880 9128 9908
rect 8941 9871 8999 9877
rect 9122 9868 9128 9880
rect 9180 9908 9186 9920
rect 9766 9908 9772 9920
rect 9180 9880 9772 9908
rect 9180 9868 9186 9880
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 9950 9908 9956 9920
rect 9911 9880 9956 9908
rect 9950 9868 9956 9880
rect 10008 9908 10014 9920
rect 10318 9908 10324 9920
rect 10008 9880 10324 9908
rect 10008 9868 10014 9880
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 11790 9908 11796 9920
rect 11751 9880 11796 9908
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13188 9908 13216 10016
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 14056 10016 15485 10044
rect 14056 10004 14062 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 14645 9979 14703 9985
rect 14645 9945 14657 9979
rect 14691 9976 14703 9979
rect 15930 9976 15936 9988
rect 14691 9948 15936 9976
rect 14691 9945 14703 9948
rect 14645 9939 14703 9945
rect 13136 9880 13216 9908
rect 13136 9868 13142 9880
rect 13354 9868 13360 9920
rect 13412 9908 13418 9920
rect 14001 9911 14059 9917
rect 14001 9908 14013 9911
rect 13412 9880 14013 9908
rect 13412 9868 13418 9880
rect 14001 9877 14013 9880
rect 14047 9877 14059 9911
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 14001 9871 14059 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 14274 9868 14280 9920
rect 14332 9908 14338 9920
rect 14660 9908 14688 9939
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 14332 9880 14688 9908
rect 14737 9911 14795 9917
rect 14332 9868 14338 9880
rect 14737 9877 14749 9911
rect 14783 9908 14795 9911
rect 15841 9911 15899 9917
rect 15841 9908 15853 9911
rect 14783 9880 15853 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 15841 9877 15853 9880
rect 15887 9877 15899 9911
rect 16298 9908 16304 9920
rect 16259 9880 16304 9908
rect 15841 9871 15899 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16574 9908 16580 9920
rect 16535 9880 16580 9908
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 2317 9707 2375 9713
rect 2317 9673 2329 9707
rect 2363 9704 2375 9707
rect 2498 9704 2504 9716
rect 2363 9676 2504 9704
rect 2363 9673 2375 9676
rect 2317 9667 2375 9673
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 7466 9704 7472 9716
rect 2648 9676 7472 9704
rect 2648 9664 2654 9676
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 16574 9704 16580 9716
rect 9508 9676 16580 9704
rect 1762 9636 1768 9648
rect 1723 9608 1768 9636
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 2038 9596 2044 9648
rect 2096 9636 2102 9648
rect 3786 9636 3792 9648
rect 2096 9608 3792 9636
rect 2096 9596 2102 9608
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 4617 9639 4675 9645
rect 4617 9605 4629 9639
rect 4663 9636 4675 9639
rect 5534 9636 5540 9648
rect 4663 9608 5540 9636
rect 4663 9605 4675 9608
rect 4617 9599 4675 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 5684 9608 5729 9636
rect 5684 9596 5690 9608
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 6052 9608 7021 9636
rect 6052 9596 6058 9608
rect 7009 9605 7021 9608
rect 7055 9605 7067 9639
rect 7190 9636 7196 9648
rect 7151 9608 7196 9636
rect 7009 9599 7067 9605
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 9508 9645 9536 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18601 9707 18659 9713
rect 18601 9704 18613 9707
rect 18012 9676 18613 9704
rect 18012 9664 18018 9676
rect 18601 9673 18613 9676
rect 18647 9704 18659 9707
rect 18969 9707 19027 9713
rect 18969 9704 18981 9707
rect 18647 9676 18981 9704
rect 18647 9673 18659 9676
rect 18601 9667 18659 9673
rect 18969 9673 18981 9676
rect 19015 9704 19027 9707
rect 19150 9704 19156 9716
rect 19015 9676 19156 9704
rect 19015 9673 19027 9676
rect 18969 9667 19027 9673
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 20438 9704 20444 9716
rect 20399 9676 20444 9704
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 9493 9639 9551 9645
rect 9493 9605 9505 9639
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9600 9608 13952 9636
rect 2958 9568 2964 9580
rect 2871 9540 2964 9568
rect 2958 9528 2964 9540
rect 3016 9568 3022 9580
rect 4062 9568 4068 9580
rect 3016 9540 4068 9568
rect 3016 9528 3022 9540
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4764 9540 5181 9568
rect 4764 9528 4770 9540
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5408 9540 6193 9568
rect 5408 9528 5414 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 1360 9472 2789 9500
rect 1360 9460 1366 9472
rect 2777 9469 2789 9472
rect 2823 9500 2835 9503
rect 3418 9500 3424 9512
rect 2823 9472 3424 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 7760 9500 7788 9531
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8205 9571 8263 9577
rect 8205 9568 8217 9571
rect 7892 9540 8217 9568
rect 7892 9528 7898 9540
rect 8205 9537 8217 9540
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8628 9540 9045 9568
rect 8628 9528 8634 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 8294 9500 8300 9512
rect 3835 9472 8300 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 7116 9444 7144 9472
rect 8294 9460 8300 9472
rect 8352 9500 8358 9512
rect 8754 9500 8760 9512
rect 8352 9472 8760 9500
rect 8352 9460 8358 9472
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 9508 9500 9536 9599
rect 8895 9472 9536 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9432 4583 9435
rect 4571 9404 5120 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 1210 9324 1216 9376
rect 1268 9364 1274 9376
rect 2133 9367 2191 9373
rect 2133 9364 2145 9367
rect 1268 9336 2145 9364
rect 1268 9324 1274 9336
rect 2133 9333 2145 9336
rect 2179 9364 2191 9367
rect 2682 9364 2688 9376
rect 2179 9336 2688 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 4065 9367 4123 9373
rect 4065 9364 4077 9367
rect 3292 9336 4077 9364
rect 3292 9324 3298 9336
rect 4065 9333 4077 9336
rect 4111 9364 4123 9367
rect 4982 9364 4988 9376
rect 4111 9336 4988 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5092 9373 5120 9404
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 6089 9435 6147 9441
rect 6089 9432 6101 9435
rect 5960 9404 6101 9432
rect 5960 9392 5966 9404
rect 6089 9401 6101 9404
rect 6135 9401 6147 9435
rect 6089 9395 6147 9401
rect 7098 9392 7104 9444
rect 7156 9392 7162 9444
rect 7653 9435 7711 9441
rect 7653 9401 7665 9435
rect 7699 9432 7711 9435
rect 9600 9432 9628 9608
rect 9674 9528 9680 9580
rect 9732 9528 9738 9580
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 10962 9568 10968 9580
rect 10183 9540 10968 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 12434 9568 12440 9580
rect 11931 9540 12440 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13924 9568 13952 9608
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 16942 9636 16948 9648
rect 15804 9608 16948 9636
rect 15804 9596 15810 9608
rect 16942 9596 16948 9608
rect 17000 9636 17006 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17000 9608 18245 9636
rect 17000 9596 17006 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 20806 9636 20812 9648
rect 20767 9608 20812 9636
rect 18233 9599 18291 9605
rect 20806 9596 20812 9608
rect 20864 9636 20870 9648
rect 21177 9639 21235 9645
rect 21177 9636 21189 9639
rect 20864 9608 21189 9636
rect 20864 9596 20870 9608
rect 21177 9605 21189 9608
rect 21223 9605 21235 9639
rect 21177 9599 21235 9605
rect 13924 9540 14044 9568
rect 9692 9500 9720 9528
rect 11057 9503 11115 9509
rect 11057 9500 11069 9503
rect 9692 9472 11069 9500
rect 11057 9469 11069 9472
rect 11103 9500 11115 9503
rect 11146 9500 11152 9512
rect 11103 9472 11152 9500
rect 11103 9469 11115 9472
rect 11057 9463 11115 9469
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11514 9460 11520 9512
rect 11572 9500 11578 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11572 9472 11713 9500
rect 11572 9460 11578 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 13265 9503 13323 9509
rect 13265 9500 13277 9503
rect 11701 9463 11759 9469
rect 12544 9472 13277 9500
rect 9953 9435 10011 9441
rect 9953 9432 9965 9435
rect 7699 9404 9628 9432
rect 9692 9404 9965 9432
rect 7699 9401 7711 9404
rect 7653 9395 7711 9401
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5442 9364 5448 9376
rect 5123 9336 5448 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 6178 9364 6184 9376
rect 6043 9336 6184 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 7742 9364 7748 9376
rect 7607 9336 7748 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8496 9373 8524 9404
rect 8481 9367 8539 9373
rect 8481 9333 8493 9367
rect 8527 9333 8539 9367
rect 8481 9327 8539 9333
rect 8941 9367 8999 9373
rect 8941 9333 8953 9367
rect 8987 9364 8999 9367
rect 9214 9364 9220 9376
rect 8987 9336 9220 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 9692 9364 9720 9404
rect 9953 9401 9965 9404
rect 9999 9432 10011 9435
rect 10505 9435 10563 9441
rect 10505 9432 10517 9435
rect 9999 9404 10517 9432
rect 9999 9401 10011 9404
rect 9953 9395 10011 9401
rect 10505 9401 10517 9404
rect 10551 9432 10563 9435
rect 10594 9432 10600 9444
rect 10551 9404 10600 9432
rect 10551 9401 10563 9404
rect 10505 9395 10563 9401
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 12544 9432 12572 9472
rect 13265 9469 13277 9472
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13872 9472 13921 9500
rect 13872 9460 13878 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 12802 9432 12808 9444
rect 11256 9404 12572 9432
rect 12715 9404 12808 9432
rect 9456 9336 9720 9364
rect 9456 9324 9462 9336
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 11256 9373 11284 9404
rect 12802 9392 12808 9404
rect 12860 9432 12866 9444
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 12860 9404 13461 9432
rect 12860 9392 12866 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 14016 9432 14044 9540
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 15068 9540 17049 9568
rect 15068 9528 15074 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 18656 9540 19472 9568
rect 18656 9528 18662 9540
rect 14182 9509 14188 9512
rect 14176 9500 14188 9509
rect 14143 9472 14188 9500
rect 14176 9463 14188 9472
rect 14182 9460 14188 9463
rect 14240 9460 14246 9512
rect 14642 9460 14648 9512
rect 14700 9500 14706 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 14700 9472 15945 9500
rect 14700 9460 14706 9472
rect 15933 9469 15945 9472
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 16206 9460 16212 9512
rect 16264 9500 16270 9512
rect 16669 9503 16727 9509
rect 16669 9500 16681 9503
rect 16264 9472 16681 9500
rect 16264 9460 16270 9472
rect 16669 9469 16681 9472
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 19444 9441 19472 9540
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 14016 9404 17417 9432
rect 13449 9395 13507 9401
rect 17405 9401 17417 9404
rect 17451 9401 17463 9435
rect 17405 9395 17463 9401
rect 19429 9435 19487 9441
rect 19429 9401 19441 9435
rect 19475 9432 19487 9435
rect 19797 9435 19855 9441
rect 19797 9432 19809 9435
rect 19475 9404 19809 9432
rect 19475 9401 19487 9404
rect 19429 9395 19487 9401
rect 19797 9401 19809 9404
rect 19843 9432 19855 9435
rect 19843 9404 20116 9432
rect 19843 9401 19855 9404
rect 19797 9395 19855 9401
rect 20088 9376 20116 9404
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 9824 9336 9873 9364
rect 9824 9324 9830 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 11241 9367 11299 9373
rect 11241 9333 11253 9367
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11388 9336 11621 9364
rect 11388 9324 11394 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12710 9364 12716 9376
rect 12483 9336 12716 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 12943 9336 13277 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 13265 9333 13277 9336
rect 13311 9364 13323 9367
rect 14366 9364 14372 9376
rect 13311 9336 14372 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 14608 9336 15301 9364
rect 14608 9324 14614 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 15657 9367 15715 9373
rect 15657 9333 15669 9367
rect 15703 9364 15715 9367
rect 15930 9364 15936 9376
rect 15703 9336 15936 9364
rect 15703 9333 15715 9336
rect 15657 9327 15715 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16390 9364 16396 9376
rect 16351 9336 16396 9364
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17276 9336 17785 9364
rect 17276 9324 17282 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 20070 9364 20076 9376
rect 20031 9336 20076 9364
rect 17773 9327 17831 9333
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1673 9163 1731 9169
rect 1673 9129 1685 9163
rect 1719 9160 1731 9163
rect 1719 9132 3740 9160
rect 1719 9129 1731 9132
rect 1673 9123 1731 9129
rect 2032 9095 2090 9101
rect 2032 9061 2044 9095
rect 2078 9092 2090 9095
rect 2958 9092 2964 9104
rect 2078 9064 2964 9092
rect 2078 9061 2090 9064
rect 2032 9055 2090 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 3712 9092 3740 9132
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 3844 9132 4261 9160
rect 3844 9120 3850 9132
rect 4249 9129 4261 9132
rect 4295 9160 4307 9163
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 4295 9132 4905 9160
rect 4295 9129 4307 9132
rect 4249 9123 4307 9129
rect 4893 9129 4905 9132
rect 4939 9129 4951 9163
rect 4893 9123 4951 9129
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 5626 9160 5632 9172
rect 5316 9132 5632 9160
rect 5316 9120 5322 9132
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7929 9163 7987 9169
rect 7432 9132 7696 9160
rect 7432 9120 7438 9132
rect 5350 9092 5356 9104
rect 3712 9064 5356 9092
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 6730 9052 6736 9104
rect 6788 9101 6794 9104
rect 6788 9095 6852 9101
rect 6788 9061 6806 9095
rect 6840 9092 6852 9095
rect 7668 9092 7696 9132
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8294 9160 8300 9172
rect 7975 9132 8300 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8665 9163 8723 9169
rect 8665 9129 8677 9163
rect 8711 9160 8723 9163
rect 9306 9160 9312 9172
rect 8711 9132 9312 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 12618 9160 12624 9172
rect 9539 9132 12624 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 12768 9132 14136 9160
rect 12768 9120 12774 9132
rect 8757 9095 8815 9101
rect 8757 9092 8769 9095
rect 6840 9064 7604 9092
rect 7668 9064 8769 9092
rect 6840 9061 6852 9064
rect 6788 9055 6852 9061
rect 6788 9052 6794 9055
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 1765 9027 1823 9033
rect 1765 9024 1777 9027
rect 1728 8996 1777 9024
rect 1728 8984 1734 8996
rect 1765 8993 1777 8996
rect 1811 9024 1823 9027
rect 3694 9024 3700 9036
rect 1811 8996 3700 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 4798 9024 4804 9036
rect 4759 8996 4804 9024
rect 4798 8984 4804 8996
rect 4856 9024 4862 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 4856 8996 5457 9024
rect 4856 8984 4862 8996
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 6546 9024 6552 9036
rect 6507 8996 6552 9024
rect 5445 8987 5503 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 3292 8928 3433 8956
rect 3292 8916 3298 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 5074 8956 5080 8968
rect 5035 8928 5080 8956
rect 3421 8919 3479 8925
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 7576 8956 7604 9064
rect 8757 9061 8769 9064
rect 8803 9092 8815 9095
rect 9030 9092 9036 9104
rect 8803 9064 9036 9092
rect 8803 9061 8815 9064
rect 8757 9055 8815 9061
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 9125 9095 9183 9101
rect 9125 9061 9137 9095
rect 9171 9092 9183 9095
rect 9944 9095 10002 9101
rect 9944 9092 9956 9095
rect 9171 9064 9956 9092
rect 9171 9061 9183 9064
rect 9125 9055 9183 9061
rect 9944 9061 9956 9064
rect 9990 9092 10002 9095
rect 10226 9092 10232 9104
rect 9990 9064 10232 9092
rect 9990 9061 10002 9064
rect 9944 9055 10002 9061
rect 10226 9052 10232 9064
rect 10284 9092 10290 9104
rect 10962 9092 10968 9104
rect 10284 9064 10968 9092
rect 10284 9052 10290 9064
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 12152 9095 12210 9101
rect 12152 9061 12164 9095
rect 12198 9092 12210 9095
rect 12986 9092 12992 9104
rect 12198 9064 12992 9092
rect 12198 9061 12210 9064
rect 12152 9055 12210 9061
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 14108 9092 14136 9132
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 14921 9163 14979 9169
rect 14921 9160 14933 9163
rect 14240 9132 14933 9160
rect 14240 9120 14246 9132
rect 14921 9129 14933 9132
rect 14967 9160 14979 9163
rect 15102 9160 15108 9172
rect 14967 9132 15108 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 19429 9163 19487 9169
rect 19429 9160 19441 9163
rect 19208 9132 19441 9160
rect 19208 9120 19214 9132
rect 19429 9129 19441 9132
rect 19475 9129 19487 9163
rect 19429 9123 19487 9129
rect 17126 9092 17132 9104
rect 13320 9064 13952 9092
rect 14108 9064 17132 9092
rect 13320 9052 13326 9064
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 11698 9024 11704 9036
rect 8352 8996 11704 9024
rect 8352 8984 8358 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 11882 8984 11888 8996
rect 11940 9024 11946 9036
rect 13446 9024 13452 9036
rect 11940 8996 13452 9024
rect 11940 8984 11946 8996
rect 13446 8984 13452 8996
rect 13504 9024 13510 9036
rect 13814 9033 13820 9036
rect 13541 9027 13599 9033
rect 13541 9024 13553 9027
rect 13504 8996 13553 9024
rect 13504 8984 13510 8996
rect 13541 8993 13553 8996
rect 13587 8993 13599 9027
rect 13808 9024 13820 9033
rect 13775 8996 13820 9024
rect 13541 8987 13599 8993
rect 13808 8987 13820 8996
rect 13814 8984 13820 8987
rect 13872 8984 13878 9036
rect 13924 9024 13952 9064
rect 17126 9052 17132 9064
rect 17184 9092 17190 9104
rect 17589 9095 17647 9101
rect 17589 9092 17601 9095
rect 17184 9064 17601 9092
rect 17184 9052 17190 9064
rect 17589 9061 17601 9064
rect 17635 9061 17647 9095
rect 17589 9055 17647 9061
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 19797 9095 19855 9101
rect 19797 9092 19809 9095
rect 17920 9064 19809 9092
rect 17920 9052 17926 9064
rect 19797 9061 19809 9064
rect 19843 9092 19855 9095
rect 20165 9095 20223 9101
rect 20165 9092 20177 9095
rect 19843 9064 20177 9092
rect 19843 9061 19855 9064
rect 19797 9055 19855 9061
rect 20165 9061 20177 9064
rect 20211 9092 20223 9095
rect 20714 9092 20720 9104
rect 20211 9064 20720 9092
rect 20211 9061 20223 9064
rect 20165 9055 20223 9061
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 14550 9024 14556 9036
rect 13924 8996 14556 9024
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 17221 9027 17279 9033
rect 17221 9024 17233 9027
rect 16908 8996 17233 9024
rect 16908 8984 16914 8996
rect 17221 8993 17233 8996
rect 17267 8993 17279 9027
rect 17221 8987 17279 8993
rect 8570 8956 8576 8968
rect 5592 8928 6500 8956
rect 7576 8928 8576 8956
rect 5592 8916 5598 8928
rect 3326 8848 3332 8900
rect 3384 8888 3390 8900
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 3384 8860 3801 8888
rect 3384 8848 3390 8860
rect 3789 8857 3801 8860
rect 3835 8888 3847 8891
rect 6086 8888 6092 8900
rect 3835 8860 6092 8888
rect 3835 8857 3847 8860
rect 3789 8851 3847 8857
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 6365 8891 6423 8897
rect 6365 8888 6377 8891
rect 6236 8860 6377 8888
rect 6236 8848 6242 8860
rect 6365 8857 6377 8860
rect 6411 8857 6423 8891
rect 6365 8851 6423 8857
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 3510 8820 3516 8832
rect 3191 8792 3516 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 5074 8820 5080 8832
rect 4479 8792 5080 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5960 8792 6009 8820
rect 5960 8780 5966 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 6472 8820 6500 8928
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8956 8999 8959
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8987 8928 9137 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9674 8956 9680 8968
rect 9635 8928 9680 8956
rect 9125 8919 9183 8925
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 11422 8956 11428 8968
rect 10888 8928 11428 8956
rect 8297 8891 8355 8897
rect 8297 8857 8309 8891
rect 8343 8888 8355 8891
rect 8754 8888 8760 8900
rect 8343 8860 8760 8888
rect 8343 8857 8355 8860
rect 8297 8851 8355 8857
rect 8754 8848 8760 8860
rect 8812 8888 8818 8900
rect 9493 8891 9551 8897
rect 9493 8888 9505 8891
rect 8812 8860 9505 8888
rect 8812 8848 8818 8860
rect 9493 8857 9505 8860
rect 9539 8857 9551 8891
rect 9493 8851 9551 8857
rect 10888 8832 10916 8928
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8956 15347 8959
rect 15562 8956 15568 8968
rect 15335 8928 15568 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 16114 8956 16120 8968
rect 16075 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8956 16178 8968
rect 17770 8956 17776 8968
rect 16172 8928 17776 8956
rect 16172 8916 16178 8928
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11020 8860 11183 8888
rect 11020 8848 11026 8860
rect 10778 8820 10784 8832
rect 6472 8792 10784 8820
rect 5997 8783 6055 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10928 8792 11069 8820
rect 10928 8780 10934 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11155 8820 11183 8860
rect 11514 8848 11520 8900
rect 11572 8888 11578 8900
rect 11698 8888 11704 8900
rect 11572 8860 11704 8888
rect 11572 8848 11578 8860
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 15010 8848 15016 8900
rect 15068 8888 15074 8900
rect 16853 8891 16911 8897
rect 16853 8888 16865 8891
rect 15068 8860 16865 8888
rect 15068 8848 15074 8860
rect 16853 8857 16865 8860
rect 16899 8857 16911 8891
rect 16853 8851 16911 8857
rect 18049 8891 18107 8897
rect 18049 8857 18061 8891
rect 18095 8888 18107 8891
rect 18598 8888 18604 8900
rect 18095 8860 18604 8888
rect 18095 8857 18107 8860
rect 18049 8851 18107 8857
rect 18598 8848 18604 8860
rect 18656 8848 18662 8900
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 11155 8792 13277 8820
rect 11057 8783 11115 8789
rect 13265 8789 13277 8792
rect 13311 8820 13323 8823
rect 13538 8820 13544 8832
rect 13311 8792 13544 8820
rect 13311 8789 13323 8792
rect 13265 8783 13323 8789
rect 13538 8780 13544 8792
rect 13596 8820 13602 8832
rect 15749 8823 15807 8829
rect 15749 8820 15761 8823
rect 13596 8792 15761 8820
rect 13596 8780 13602 8792
rect 15749 8789 15761 8792
rect 15795 8789 15807 8823
rect 16574 8820 16580 8832
rect 16535 8792 16580 8820
rect 15749 8783 15807 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 18417 8823 18475 8829
rect 18417 8789 18429 8823
rect 18463 8820 18475 8823
rect 18506 8820 18512 8832
rect 18463 8792 18512 8820
rect 18463 8789 18475 8792
rect 18417 8783 18475 8789
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 18690 8820 18696 8832
rect 18651 8792 18696 8820
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 19061 8823 19119 8829
rect 19061 8820 19073 8823
rect 18840 8792 19073 8820
rect 18840 8780 18846 8792
rect 19061 8789 19073 8792
rect 19107 8789 19119 8823
rect 19061 8783 19119 8789
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 20625 8823 20683 8829
rect 20625 8820 20637 8823
rect 20128 8792 20637 8820
rect 20128 8780 20134 8792
rect 20625 8789 20637 8792
rect 20671 8820 20683 8823
rect 21174 8820 21180 8832
rect 20671 8792 21180 8820
rect 20671 8789 20683 8792
rect 20625 8783 20683 8789
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 1857 8619 1915 8625
rect 1857 8585 1869 8619
rect 1903 8616 1915 8619
rect 2133 8619 2191 8625
rect 2133 8616 2145 8619
rect 1903 8588 2145 8616
rect 1903 8585 1915 8588
rect 1857 8579 1915 8585
rect 2133 8585 2145 8588
rect 2179 8616 2191 8619
rect 2406 8616 2412 8628
rect 2179 8588 2412 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 2501 8619 2559 8625
rect 2501 8585 2513 8619
rect 2547 8616 2559 8619
rect 3326 8616 3332 8628
rect 2547 8588 3332 8616
rect 2547 8585 2559 8588
rect 2501 8579 2559 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 5258 8616 5264 8628
rect 3476 8588 5120 8616
rect 5171 8588 5264 8616
rect 3476 8576 3482 8588
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 2685 8551 2743 8557
rect 2685 8548 2697 8551
rect 2648 8520 2697 8548
rect 2648 8508 2654 8520
rect 2685 8517 2697 8520
rect 2731 8517 2743 8551
rect 3786 8548 3792 8560
rect 2685 8511 2743 8517
rect 3160 8520 3792 8548
rect 3160 8489 3188 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 5092 8480 5120 8588
rect 5258 8576 5264 8588
rect 5316 8616 5322 8628
rect 5534 8616 5540 8628
rect 5316 8588 5540 8616
rect 5316 8576 5322 8588
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6730 8616 6736 8628
rect 6052 8588 6736 8616
rect 6052 8576 6058 8588
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 6847 8588 7788 8616
rect 6454 8548 6460 8560
rect 6012 8520 6460 8548
rect 6012 8489 6040 8520
rect 6454 8508 6460 8520
rect 6512 8548 6518 8560
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 6512 8520 6561 8548
rect 6512 8508 6518 8520
rect 6549 8517 6561 8520
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5092 8452 6009 8480
rect 3237 8443 3295 8449
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 6178 8480 6184 8492
rect 6091 8452 6184 8480
rect 5997 8443 6055 8449
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3252 8412 3280 8443
rect 6178 8440 6184 8452
rect 6236 8480 6242 8492
rect 6847 8480 6875 8588
rect 7760 8548 7788 8588
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 7984 8588 8493 8616
rect 7984 8576 7990 8588
rect 8481 8585 8493 8588
rect 8527 8616 8539 8619
rect 11146 8616 11152 8628
rect 8527 8588 11152 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11606 8616 11612 8628
rect 11519 8588 11612 8616
rect 11606 8576 11612 8588
rect 11664 8616 11670 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11664 8588 11897 8616
rect 11664 8576 11670 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 12124 8588 13369 8616
rect 12124 8576 12130 8588
rect 13357 8585 13369 8588
rect 13403 8616 13415 8619
rect 13446 8616 13452 8628
rect 13403 8588 13452 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 13541 8619 13599 8625
rect 13541 8585 13553 8619
rect 13587 8616 13599 8619
rect 15010 8616 15016 8628
rect 13587 8588 15016 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15381 8619 15439 8625
rect 15120 8588 15332 8616
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 7760 8520 8217 8548
rect 8205 8517 8217 8520
rect 8251 8548 8263 8551
rect 8294 8548 8300 8560
rect 8251 8520 8300 8548
rect 8251 8517 8263 8520
rect 8205 8511 8263 8517
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 8628 8520 9168 8548
rect 8628 8508 8634 8520
rect 9140 8489 9168 8520
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9677 8551 9735 8557
rect 9677 8548 9689 8551
rect 9364 8520 9689 8548
rect 9364 8508 9370 8520
rect 9677 8517 9689 8520
rect 9723 8548 9735 8551
rect 13081 8551 13139 8557
rect 9723 8520 12296 8548
rect 9723 8517 9735 8520
rect 9677 8511 9735 8517
rect 9125 8483 9183 8489
rect 6236 8452 6875 8480
rect 8404 8452 9045 8480
rect 6236 8440 6242 8452
rect 3016 8384 3280 8412
rect 3016 8372 3022 8384
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 3881 8415 3939 8421
rect 3881 8412 3893 8415
rect 3752 8384 3893 8412
rect 3752 8372 3758 8384
rect 3881 8381 3893 8384
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4148 8415 4206 8421
rect 4148 8381 4160 8415
rect 4194 8412 4206 8415
rect 5166 8412 5172 8424
rect 4194 8384 5172 8412
rect 4194 8381 4206 8384
rect 4148 8375 4206 8381
rect 4264 8356 4292 8384
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 6454 8412 6460 8424
rect 5491 8384 6460 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 7098 8421 7104 8424
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8381 6883 8415
rect 7092 8412 7104 8421
rect 7059 8384 7104 8412
rect 6825 8375 6883 8381
rect 7092 8375 7104 8384
rect 3786 8344 3792 8356
rect 3747 8316 3792 8344
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 4246 8304 4252 8356
rect 4304 8304 4310 8356
rect 6840 8344 6868 8375
rect 7098 8372 7104 8375
rect 7156 8372 7162 8424
rect 8404 8344 8432 8452
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8628 8384 8861 8412
rect 8628 8372 8634 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 6840 8316 8432 8344
rect 9017 8344 9045 8452
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9140 8412 9168 8443
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9272 8452 9505 8480
rect 9272 8440 9278 8452
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 10226 8480 10232 8492
rect 10187 8452 10232 8480
rect 9493 8443 9551 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11563 8452 12112 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 12084 8424 12112 8452
rect 9950 8412 9956 8424
rect 9140 8384 9956 8412
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10137 8415 10195 8421
rect 10137 8381 10149 8415
rect 10183 8412 10195 8415
rect 10594 8412 10600 8424
rect 10183 8384 10600 8412
rect 10183 8381 10195 8384
rect 10137 8375 10195 8381
rect 10594 8372 10600 8384
rect 10652 8412 10658 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10652 8384 10701 8412
rect 10652 8372 10658 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 11790 8412 11796 8424
rect 11751 8384 11796 8412
rect 10689 8375 10747 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12066 8412 12072 8424
rect 12027 8384 12072 8412
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12268 8412 12296 8520
rect 13081 8517 13093 8551
rect 13127 8548 13139 8551
rect 13814 8548 13820 8560
rect 13127 8520 13820 8548
rect 13127 8517 13139 8520
rect 13081 8511 13139 8517
rect 13814 8508 13820 8520
rect 13872 8548 13878 8560
rect 13872 8520 14228 8548
rect 13872 8508 13878 8520
rect 14200 8492 14228 8520
rect 14274 8508 14280 8560
rect 14332 8548 14338 8560
rect 15120 8548 15148 8588
rect 14332 8520 15148 8548
rect 14332 8508 14338 8520
rect 15194 8508 15200 8560
rect 15252 8508 15258 8560
rect 15304 8548 15332 8588
rect 15381 8585 15393 8619
rect 15427 8616 15439 8619
rect 15562 8616 15568 8628
rect 15427 8588 15568 8616
rect 15427 8585 15439 8588
rect 15381 8579 15439 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 19705 8619 19763 8625
rect 19705 8616 19717 8619
rect 15712 8588 19717 8616
rect 15712 8576 15718 8588
rect 19705 8585 19717 8588
rect 19751 8585 19763 8619
rect 19705 8579 19763 8585
rect 20533 8619 20591 8625
rect 20533 8585 20545 8619
rect 20579 8616 20591 8619
rect 20714 8616 20720 8628
rect 20579 8588 20720 8616
rect 20579 8585 20591 8588
rect 20533 8579 20591 8585
rect 20714 8576 20720 8588
rect 20772 8616 20778 8628
rect 20809 8619 20867 8625
rect 20809 8616 20821 8619
rect 20772 8588 20821 8616
rect 20772 8576 20778 8588
rect 20809 8585 20821 8588
rect 20855 8585 20867 8619
rect 21174 8616 21180 8628
rect 21135 8588 21180 8616
rect 20809 8579 20867 8585
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 18969 8551 19027 8557
rect 18969 8548 18981 8551
rect 15304 8520 18981 8548
rect 18969 8517 18981 8520
rect 19015 8517 19027 8551
rect 18969 8511 19027 8517
rect 19150 8508 19156 8560
rect 19208 8548 19214 8560
rect 20073 8551 20131 8557
rect 20073 8548 20085 8551
rect 19208 8520 20085 8548
rect 19208 8508 19214 8520
rect 20073 8517 20085 8520
rect 20119 8517 20131 8551
rect 20073 8511 20131 8517
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12802 8480 12808 8492
rect 12483 8452 12808 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 14090 8480 14096 8492
rect 13280 8452 14096 8480
rect 13280 8412 13308 8452
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 15105 8483 15163 8489
rect 14240 8452 14285 8480
rect 14240 8440 14246 8452
rect 15105 8449 15117 8483
rect 15151 8480 15163 8483
rect 15212 8480 15240 8508
rect 15151 8452 15240 8480
rect 17405 8483 17463 8489
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17451 8452 17632 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 12268 8384 13308 8412
rect 13446 8372 13452 8424
rect 13504 8412 13510 8424
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 13504 8384 13921 8412
rect 13504 8372 13510 8384
rect 13909 8381 13921 8384
rect 13955 8381 13967 8415
rect 13909 8375 13967 8381
rect 14366 8372 14372 8424
rect 14424 8412 14430 8424
rect 14826 8412 14832 8424
rect 14424 8384 14832 8412
rect 14424 8372 14430 8384
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8412 14979 8415
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 14967 8384 15393 8412
rect 14967 8381 14979 8384
rect 14921 8375 14979 8381
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 16393 8415 16451 8421
rect 16393 8381 16405 8415
rect 16439 8412 16451 8415
rect 16850 8412 16856 8424
rect 16439 8384 16856 8412
rect 16439 8381 16451 8384
rect 16393 8375 16451 8381
rect 9674 8344 9680 8356
rect 9017 8316 9680 8344
rect 9674 8304 9680 8316
rect 9732 8304 9738 8356
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 9916 8316 10057 8344
rect 9916 8304 9922 8316
rect 10045 8313 10057 8316
rect 10091 8313 10103 8347
rect 11054 8344 11060 8356
rect 11015 8316 11060 8344
rect 10045 8307 10103 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 11885 8347 11943 8353
rect 11885 8313 11897 8347
rect 11931 8344 11943 8347
rect 12526 8344 12532 8356
rect 11931 8316 12532 8344
rect 11931 8313 11943 8316
rect 11885 8307 11943 8313
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 16408 8344 16436 8375
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17604 8412 17632 8452
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 17920 8452 18613 8480
rect 17920 8440 17926 8452
rect 18601 8449 18613 8452
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 18874 8412 18880 8424
rect 17604 8384 18880 8412
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 14568 8316 16436 8344
rect 16669 8347 16727 8353
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 3053 8279 3111 8285
rect 3053 8276 3065 8279
rect 1636 8248 3065 8276
rect 1636 8236 1642 8248
rect 3053 8245 3065 8248
rect 3099 8276 3111 8279
rect 3234 8276 3240 8288
rect 3099 8248 3240 8276
rect 3099 8245 3111 8248
rect 3053 8239 3111 8245
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 4948 8248 5457 8276
rect 4948 8236 4954 8248
rect 5445 8245 5457 8248
rect 5491 8276 5503 8279
rect 5537 8279 5595 8285
rect 5537 8276 5549 8279
rect 5491 8248 5549 8276
rect 5491 8245 5503 8248
rect 5445 8239 5503 8245
rect 5537 8245 5549 8248
rect 5583 8245 5595 8279
rect 5537 8239 5595 8245
rect 5626 8236 5632 8288
rect 5684 8276 5690 8288
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 5684 8248 5917 8276
rect 5684 8236 5690 8248
rect 5905 8245 5917 8248
rect 5951 8276 5963 8279
rect 5994 8276 6000 8288
rect 5951 8248 6000 8276
rect 5951 8245 5963 8248
rect 5905 8239 5963 8245
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 6454 8236 6460 8288
rect 6512 8276 6518 8288
rect 7190 8276 7196 8288
rect 6512 8248 7196 8276
rect 6512 8236 6518 8248
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 8202 8276 8208 8288
rect 7432 8248 8208 8276
rect 7432 8236 7438 8248
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 8812 8248 8953 8276
rect 8812 8236 8818 8248
rect 8941 8245 8953 8248
rect 8987 8245 8999 8279
rect 8941 8239 8999 8245
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 13262 8276 13268 8288
rect 9088 8248 13268 8276
rect 9088 8236 9094 8248
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 14001 8279 14059 8285
rect 14001 8245 14013 8279
rect 14047 8276 14059 8279
rect 14090 8276 14096 8288
rect 14047 8248 14096 8276
rect 14047 8245 14059 8248
rect 14001 8239 14059 8245
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 14568 8285 14596 8316
rect 16669 8313 16681 8347
rect 16715 8344 16727 8347
rect 16942 8344 16948 8356
rect 16715 8316 16948 8344
rect 16715 8313 16727 8316
rect 16669 8307 16727 8313
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 18046 8304 18052 8356
rect 18104 8344 18110 8356
rect 18690 8344 18696 8356
rect 18104 8316 18696 8344
rect 18104 8304 18110 8316
rect 18690 8304 18696 8316
rect 18748 8304 18754 8356
rect 19334 8344 19340 8356
rect 19295 8316 19340 8344
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 14553 8279 14611 8285
rect 14553 8245 14565 8279
rect 14599 8245 14611 8279
rect 15010 8276 15016 8288
rect 14971 8248 15016 8276
rect 14553 8239 14611 8245
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 15470 8236 15476 8288
rect 15528 8276 15534 8288
rect 16025 8279 16083 8285
rect 16025 8276 16037 8279
rect 15528 8248 16037 8276
rect 15528 8236 15534 8248
rect 16025 8245 16037 8248
rect 16071 8276 16083 8279
rect 17310 8276 17316 8288
rect 16071 8248 17316 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 18322 8236 18328 8288
rect 18380 8276 18386 8288
rect 18380 8248 18425 8276
rect 18380 8236 18386 8248
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2958 8032 2964 8084
rect 3016 8072 3022 8084
rect 3053 8075 3111 8081
rect 3053 8072 3065 8075
rect 3016 8044 3065 8072
rect 3016 8032 3022 8044
rect 3053 8041 3065 8044
rect 3099 8041 3111 8075
rect 3053 8035 3111 8041
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 4246 8072 4252 8084
rect 3844 8044 4252 8072
rect 3844 8032 3850 8044
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 4706 8072 4712 8084
rect 4387 8044 4712 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 4890 8072 4896 8084
rect 4847 8044 4896 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 5000 8044 6776 8072
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 5000 8004 5028 8044
rect 4028 7976 5028 8004
rect 5712 8007 5770 8013
rect 4028 7964 4034 7976
rect 5712 7973 5724 8007
rect 5758 8004 5770 8007
rect 6178 8004 6184 8016
rect 5758 7976 6184 8004
rect 5758 7973 5770 7976
rect 5712 7967 5770 7973
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 1946 7945 1952 7948
rect 1940 7936 1952 7945
rect 1907 7908 1952 7936
rect 1940 7899 1952 7908
rect 1946 7896 1952 7899
rect 2004 7896 2010 7948
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 3752 7908 5365 7936
rect 3752 7896 3758 7908
rect 5353 7905 5365 7908
rect 5399 7936 5411 7939
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5399 7908 5457 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5552 7908 6684 7936
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 4890 7828 4896 7880
rect 4948 7868 4954 7880
rect 5077 7871 5135 7877
rect 4948 7840 4993 7868
rect 4948 7828 4954 7840
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5166 7868 5172 7880
rect 5123 7840 5172 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5166 7828 5172 7840
rect 5224 7868 5230 7880
rect 5552 7868 5580 7908
rect 5224 7840 5580 7868
rect 5224 7828 5230 7840
rect 3050 7760 3056 7812
rect 3108 7800 3114 7812
rect 4798 7800 4804 7812
rect 3108 7772 4804 7800
rect 3108 7760 3114 7772
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 3513 7735 3571 7741
rect 3513 7701 3525 7735
rect 3559 7732 3571 7735
rect 3602 7732 3608 7744
rect 3559 7704 3608 7732
rect 3559 7701 3571 7704
rect 3513 7695 3571 7701
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 3786 7732 3792 7744
rect 3747 7704 3792 7732
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 4706 7732 4712 7744
rect 4479 7704 4712 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 5166 7692 5172 7744
rect 5224 7732 5230 7744
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 5224 7704 5365 7732
rect 5224 7692 5230 7704
rect 5353 7701 5365 7704
rect 5399 7732 5411 7735
rect 6454 7732 6460 7744
rect 5399 7704 6460 7732
rect 5399 7701 5411 7704
rect 5353 7695 5411 7701
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 6656 7732 6684 7908
rect 6748 7868 6776 8044
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 6972 8044 7113 8072
rect 6972 8032 6978 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 8846 8072 8852 8084
rect 8807 8044 8852 8072
rect 7101 8035 7159 8041
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 14274 8072 14280 8084
rect 8956 8044 14280 8072
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 8956 8004 8984 8044
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 15013 8075 15071 8081
rect 15013 8041 15025 8075
rect 15059 8072 15071 8075
rect 15102 8072 15108 8084
rect 15059 8044 15108 8072
rect 15059 8041 15071 8044
rect 15013 8035 15071 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 16666 8072 16672 8084
rect 15804 8044 16672 8072
rect 15804 8032 15810 8044
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17310 8072 17316 8084
rect 17271 8044 17316 8072
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 18690 8072 18696 8084
rect 17552 8044 18696 8072
rect 17552 8032 17558 8044
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 21085 8075 21143 8081
rect 21085 8072 21097 8075
rect 20772 8044 21097 8072
rect 20772 8032 20778 8044
rect 21085 8041 21097 8044
rect 21131 8041 21143 8075
rect 21085 8035 21143 8041
rect 15470 8004 15476 8016
rect 7248 7976 8984 8004
rect 9140 7976 15476 8004
rect 7248 7964 7254 7976
rect 7282 7936 7288 7948
rect 7243 7908 7288 7936
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 9030 7936 9036 7948
rect 7392 7908 9036 7936
rect 7392 7868 7420 7908
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 6748 7840 7420 7868
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 9140 7868 9168 7976
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 16574 8004 16580 8016
rect 15764 7976 16580 8004
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 10502 7936 10508 7948
rect 9272 7908 10508 7936
rect 9272 7896 9278 7908
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 11140 7939 11198 7945
rect 11140 7905 11152 7939
rect 11186 7936 11198 7939
rect 12066 7936 12072 7948
rect 11186 7908 12072 7936
rect 11186 7905 11198 7908
rect 11140 7899 11198 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 15764 7936 15792 7976
rect 16574 7964 16580 7976
rect 16632 8004 16638 8016
rect 17957 8007 18015 8013
rect 17957 8004 17969 8007
rect 16632 7976 17969 8004
rect 16632 7964 16638 7976
rect 17957 7973 17969 7976
rect 18003 7973 18015 8007
rect 17957 7967 18015 7973
rect 14240 7908 15792 7936
rect 14240 7896 14246 7908
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 16189 7939 16247 7945
rect 16189 7936 16201 7939
rect 15896 7908 16201 7936
rect 15896 7896 15902 7908
rect 16189 7905 16201 7908
rect 16235 7905 16247 7939
rect 16189 7899 16247 7905
rect 16666 7896 16672 7948
rect 16724 7936 16730 7948
rect 20533 7939 20591 7945
rect 20533 7936 20545 7939
rect 16724 7908 20545 7936
rect 16724 7896 16730 7908
rect 20533 7905 20545 7908
rect 20579 7905 20591 7939
rect 20533 7899 20591 7905
rect 7524 7840 9168 7868
rect 7524 7828 7530 7840
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 9732 7840 10885 7868
rect 9732 7828 9738 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7868 12587 7871
rect 12802 7868 12808 7880
rect 12575 7840 12808 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 15746 7868 15752 7880
rect 12943 7840 15752 7868
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 8573 7803 8631 7809
rect 8573 7769 8585 7803
rect 8619 7800 8631 7803
rect 9030 7800 9036 7812
rect 8619 7772 9036 7800
rect 8619 7769 8631 7772
rect 8573 7763 8631 7769
rect 9030 7760 9036 7772
rect 9088 7800 9094 7812
rect 9217 7803 9275 7809
rect 9217 7800 9229 7803
rect 9088 7772 9229 7800
rect 9088 7760 9094 7772
rect 9217 7769 9229 7772
rect 9263 7800 9275 7803
rect 9582 7800 9588 7812
rect 9263 7772 9588 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 9858 7760 9864 7812
rect 9916 7800 9922 7812
rect 10045 7803 10103 7809
rect 10045 7800 10057 7803
rect 9916 7772 10057 7800
rect 9916 7760 9922 7772
rect 10045 7769 10057 7772
rect 10091 7769 10103 7803
rect 13357 7803 13415 7809
rect 13357 7800 13369 7803
rect 10045 7763 10103 7769
rect 12268 7772 13369 7800
rect 6825 7735 6883 7741
rect 6825 7732 6837 7735
rect 6656 7704 6837 7732
rect 6825 7701 6837 7704
rect 6871 7732 6883 7735
rect 7190 7732 7196 7744
rect 6871 7704 7196 7732
rect 6871 7701 6883 7704
rect 6825 7695 6883 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7340 7704 7573 7732
rect 7340 7692 7346 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 7742 7692 7748 7744
rect 7800 7732 7806 7744
rect 7929 7735 7987 7741
rect 7929 7732 7941 7735
rect 7800 7704 7941 7732
rect 7800 7692 7806 7704
rect 7929 7701 7941 7704
rect 7975 7701 7987 7735
rect 7929 7695 7987 7701
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 9122 7732 9128 7744
rect 8076 7704 9128 7732
rect 8076 7692 8082 7704
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 11790 7732 11796 7744
rect 10827 7704 11796 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 11790 7692 11796 7704
rect 11848 7732 11854 7744
rect 12268 7741 12296 7772
rect 13096 7744 13124 7772
rect 13357 7769 13369 7772
rect 13403 7769 13415 7803
rect 13357 7763 13415 7769
rect 14001 7803 14059 7809
rect 14001 7769 14013 7803
rect 14047 7800 14059 7803
rect 14090 7800 14096 7812
rect 14047 7772 14096 7800
rect 14047 7769 14059 7772
rect 14001 7763 14059 7769
rect 14090 7760 14096 7772
rect 14148 7800 14154 7812
rect 15102 7800 15108 7812
rect 14148 7772 15108 7800
rect 14148 7760 14154 7772
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 15286 7760 15292 7812
rect 15344 7800 15350 7812
rect 15562 7800 15568 7812
rect 15344 7772 15568 7800
rect 15344 7760 15350 7772
rect 15562 7760 15568 7772
rect 15620 7800 15626 7812
rect 15948 7800 15976 7831
rect 16942 7828 16948 7880
rect 17000 7868 17006 7880
rect 19061 7871 19119 7877
rect 19061 7868 19073 7871
rect 17000 7840 19073 7868
rect 17000 7828 17006 7840
rect 19061 7837 19073 7840
rect 19107 7837 19119 7871
rect 19061 7831 19119 7837
rect 15620 7772 15976 7800
rect 15620 7760 15626 7772
rect 17034 7760 17040 7812
rect 17092 7800 17098 7812
rect 18325 7803 18383 7809
rect 18325 7800 18337 7803
rect 17092 7772 18337 7800
rect 17092 7760 17098 7772
rect 18325 7769 18337 7772
rect 18371 7769 18383 7803
rect 18325 7763 18383 7769
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 11848 7704 12265 7732
rect 11848 7692 11854 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 12805 7735 12863 7741
rect 12805 7732 12817 7735
rect 12768 7704 12817 7732
rect 12768 7692 12774 7704
rect 12805 7701 12817 7704
rect 12851 7701 12863 7735
rect 12986 7732 12992 7744
rect 12947 7704 12992 7732
rect 12805 7695 12863 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13078 7692 13084 7744
rect 13136 7692 13142 7744
rect 14550 7732 14556 7744
rect 14511 7704 14556 7732
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 15838 7732 15844 7744
rect 15799 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 15930 7692 15936 7744
rect 15988 7732 15994 7744
rect 17589 7735 17647 7741
rect 17589 7732 17601 7735
rect 15988 7704 17601 7732
rect 15988 7692 15994 7704
rect 17589 7701 17601 7704
rect 17635 7701 17647 7735
rect 17589 7695 17647 7701
rect 17770 7692 17776 7744
rect 17828 7732 17834 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 17828 7704 18705 7732
rect 17828 7692 17834 7704
rect 18693 7701 18705 7704
rect 18739 7701 18751 7735
rect 19518 7732 19524 7744
rect 19479 7704 19524 7732
rect 18693 7695 18751 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 19794 7732 19800 7744
rect 19755 7704 19800 7732
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 20162 7732 20168 7744
rect 20123 7704 20168 7732
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 3050 7528 3056 7540
rect 3011 7500 3056 7528
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3200 7500 4077 7528
rect 3200 7488 3206 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 4065 7491 4123 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4948 7500 5089 7528
rect 4948 7488 4954 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5258 7528 5264 7540
rect 5077 7491 5135 7497
rect 5184 7500 5264 7528
rect 2041 7463 2099 7469
rect 2041 7429 2053 7463
rect 2087 7460 2099 7463
rect 4430 7460 4436 7472
rect 2087 7432 4436 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 4614 7420 4620 7472
rect 4672 7420 4678 7472
rect 5184 7460 5212 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 6730 7528 6736 7540
rect 5868 7500 6736 7528
rect 5868 7488 5874 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 9030 7528 9036 7540
rect 7668 7500 8616 7528
rect 8991 7500 9036 7528
rect 4724 7432 5212 7460
rect 5276 7432 5755 7460
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3510 7392 3516 7404
rect 2731 7364 3516 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 3510 7352 3516 7364
rect 3568 7392 3574 7404
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 3568 7364 3617 7392
rect 3568 7352 3574 7364
rect 3605 7361 3617 7364
rect 3651 7392 3663 7395
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3651 7364 3893 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 3881 7361 3893 7364
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4632 7392 4660 7420
rect 4724 7401 4752 7432
rect 4571 7364 4660 7392
rect 4709 7395 4767 7401
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 5276 7392 5304 7432
rect 5626 7392 5632 7404
rect 5132 7364 5304 7392
rect 5587 7364 5632 7392
rect 5132 7352 5138 7364
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5727 7392 5755 7432
rect 5994 7420 6000 7472
rect 6052 7460 6058 7472
rect 6457 7463 6515 7469
rect 6457 7460 6469 7463
rect 6052 7432 6469 7460
rect 6052 7420 6058 7432
rect 6457 7429 6469 7432
rect 6503 7429 6515 7463
rect 7466 7460 7472 7472
rect 6457 7423 6515 7429
rect 6564 7432 7472 7460
rect 6564 7392 6592 7432
rect 7466 7420 7472 7432
rect 7524 7420 7530 7472
rect 5727 7364 6592 7392
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7668 7401 7696 7500
rect 8588 7460 8616 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 12710 7528 12716 7540
rect 9180 7500 12716 7528
rect 9180 7488 9186 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 12820 7500 15577 7528
rect 8588 7432 9260 7460
rect 9232 7404 9260 7432
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 11882 7460 11888 7472
rect 10560 7432 11888 7460
rect 10560 7420 10566 7432
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 12342 7460 12348 7472
rect 12216 7432 12348 7460
rect 12216 7420 12222 7432
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 12437 7463 12495 7469
rect 12437 7429 12449 7463
rect 12483 7460 12495 7463
rect 12618 7460 12624 7472
rect 12483 7432 12624 7460
rect 12483 7429 12495 7432
rect 12437 7423 12495 7429
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 7653 7395 7711 7401
rect 6880 7364 7604 7392
rect 6880 7352 6886 7364
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 3752 7296 5549 7324
rect 3752 7284 3758 7296
rect 5537 7293 5549 7296
rect 5583 7324 5595 7327
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5583 7296 6101 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 7576 7324 7604 7364
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9309 7395 9367 7401
rect 9309 7392 9321 7395
rect 9272 7364 9321 7392
rect 9272 7352 9278 7364
rect 9309 7361 9321 7364
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 11609 7395 11667 7401
rect 11609 7361 11621 7395
rect 11655 7392 11667 7395
rect 12066 7392 12072 7404
rect 11655 7364 12072 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 12066 7352 12072 7364
rect 12124 7392 12130 7404
rect 12820 7392 12848 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 15565 7491 15623 7497
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 16390 7528 16396 7540
rect 16347 7500 16396 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16482 7488 16488 7540
rect 16540 7528 16546 7540
rect 18509 7531 18567 7537
rect 18509 7528 18521 7531
rect 16540 7500 18521 7528
rect 16540 7488 16546 7500
rect 18509 7497 18521 7500
rect 18555 7528 18567 7531
rect 18601 7531 18659 7537
rect 18601 7528 18613 7531
rect 18555 7500 18613 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 18601 7497 18613 7500
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 19337 7531 19395 7537
rect 19337 7528 19349 7531
rect 18840 7500 19349 7528
rect 18840 7488 18846 7500
rect 19337 7497 19349 7500
rect 19383 7497 19395 7531
rect 19337 7491 19395 7497
rect 15470 7420 15476 7472
rect 15528 7460 15534 7472
rect 20809 7463 20867 7469
rect 20809 7460 20821 7463
rect 15528 7432 20821 7460
rect 15528 7420 15534 7432
rect 20809 7429 20821 7432
rect 20855 7429 20867 7463
rect 20809 7423 20867 7429
rect 13078 7392 13084 7404
rect 12124 7364 12848 7392
rect 13039 7364 13084 7392
rect 12124 7352 12130 7364
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 13320 7364 14320 7392
rect 13320 7352 13326 7364
rect 12802 7324 12808 7336
rect 7576 7296 9444 7324
rect 6089 7287 6147 7293
rect 9416 7268 9444 7296
rect 9692 7296 12204 7324
rect 12763 7296 12808 7324
rect 2409 7259 2467 7265
rect 2409 7256 2421 7259
rect 1872 7228 2421 7256
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 1872 7197 1900 7228
rect 2409 7225 2421 7228
rect 2455 7225 2467 7259
rect 2409 7219 2467 7225
rect 3326 7216 3332 7268
rect 3384 7256 3390 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 3384 7228 3525 7256
rect 3384 7216 3390 7228
rect 3513 7225 3525 7228
rect 3559 7256 3571 7259
rect 3970 7256 3976 7268
rect 3559 7228 3976 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3970 7216 3976 7228
rect 4028 7216 4034 7268
rect 4433 7259 4491 7265
rect 4433 7225 4445 7259
rect 4479 7256 4491 7259
rect 5074 7256 5080 7268
rect 4479 7228 5080 7256
rect 4479 7225 4491 7228
rect 4433 7219 4491 7225
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 7926 7265 7932 7268
rect 5184 7228 7328 7256
rect 1857 7191 1915 7197
rect 1857 7188 1869 7191
rect 1820 7160 1869 7188
rect 1820 7148 1826 7160
rect 1857 7157 1869 7160
rect 1903 7157 1915 7191
rect 1857 7151 1915 7157
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 3200 7160 3433 7188
rect 3200 7148 3206 7160
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3421 7151 3479 7157
rect 3881 7191 3939 7197
rect 3881 7157 3893 7191
rect 3927 7188 3939 7191
rect 5184 7188 5212 7228
rect 3927 7160 5212 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 5408 7160 5457 7188
rect 5408 7148 5414 7160
rect 5445 7157 5457 7160
rect 5491 7157 5503 7191
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 5445 7151 5503 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7300 7188 7328 7228
rect 7920 7219 7932 7265
rect 7984 7256 7990 7268
rect 8018 7256 8024 7268
rect 7984 7228 8024 7256
rect 7926 7216 7932 7219
rect 7984 7216 7990 7228
rect 8018 7216 8024 7228
rect 8076 7256 8082 7268
rect 9306 7256 9312 7268
rect 8076 7228 9312 7256
rect 8076 7216 8082 7228
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 9398 7216 9404 7268
rect 9456 7216 9462 7268
rect 9582 7265 9588 7268
rect 9565 7259 9588 7265
rect 9565 7225 9577 7259
rect 9565 7219 9588 7225
rect 9582 7216 9588 7219
rect 9640 7216 9646 7268
rect 9692 7188 9720 7296
rect 12176 7256 12204 7296
rect 12802 7284 12808 7296
rect 12860 7324 12866 7336
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 12860 7296 13461 7324
rect 12860 7284 12866 7296
rect 13449 7293 13461 7296
rect 13495 7293 13507 7327
rect 13449 7287 13507 7293
rect 13538 7284 13544 7336
rect 13596 7324 13602 7336
rect 14182 7324 14188 7336
rect 13596 7296 14188 7324
rect 13596 7284 13602 7296
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 14292 7324 14320 7364
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 16022 7392 16028 7404
rect 15252 7364 16028 7392
rect 15252 7352 15258 7364
rect 16022 7352 16028 7364
rect 16080 7392 16086 7404
rect 16945 7395 17003 7401
rect 16080 7364 16896 7392
rect 16080 7352 16086 7364
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 14292 7296 16129 7324
rect 16117 7293 16129 7296
rect 16163 7324 16175 7327
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 16163 7296 16773 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 16868 7324 16896 7364
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17310 7392 17316 7404
rect 16991 7364 17316 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 20441 7395 20499 7401
rect 20441 7392 20453 7395
rect 18012 7364 20453 7392
rect 18012 7352 18018 7364
rect 20441 7361 20453 7364
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 18509 7327 18567 7333
rect 16868 7296 17172 7324
rect 16761 7287 16819 7293
rect 14452 7259 14510 7265
rect 10980 7228 12112 7256
rect 12176 7228 14136 7256
rect 7300 7160 9720 7188
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 10980 7197 11008 7228
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10560 7160 10701 7188
rect 10560 7148 10566 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11296 7160 11345 7188
rect 11296 7148 11302 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 11425 7191 11483 7197
rect 11425 7157 11437 7191
rect 11471 7188 11483 7191
rect 11698 7188 11704 7200
rect 11471 7160 11704 7188
rect 11471 7157 11483 7160
rect 11425 7151 11483 7157
rect 11698 7148 11704 7160
rect 11756 7188 11762 7200
rect 11977 7191 12035 7197
rect 11977 7188 11989 7191
rect 11756 7160 11989 7188
rect 11756 7148 11762 7160
rect 11977 7157 11989 7160
rect 12023 7157 12035 7191
rect 12084 7188 12112 7228
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12084 7160 12909 7188
rect 11977 7151 12035 7157
rect 12897 7157 12909 7160
rect 12943 7188 12955 7191
rect 13814 7188 13820 7200
rect 12943 7160 13820 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 13998 7188 14004 7200
rect 13959 7160 14004 7188
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14108 7188 14136 7228
rect 14452 7225 14464 7259
rect 14498 7256 14510 7259
rect 14550 7256 14556 7268
rect 14498 7228 14556 7256
rect 14498 7225 14510 7228
rect 14452 7219 14510 7225
rect 14550 7216 14556 7228
rect 14608 7216 14614 7268
rect 16669 7259 16727 7265
rect 16669 7225 16681 7259
rect 16715 7256 16727 7259
rect 17144 7256 17172 7296
rect 18509 7293 18521 7327
rect 18555 7324 18567 7327
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18555 7296 18981 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 18969 7293 18981 7296
rect 19015 7324 19027 7327
rect 19150 7324 19156 7336
rect 19015 7296 19156 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 21177 7259 21235 7265
rect 21177 7256 21189 7259
rect 16715 7228 17080 7256
rect 17144 7228 21189 7256
rect 16715 7225 16727 7228
rect 16669 7219 16727 7225
rect 16482 7188 16488 7200
rect 14108 7160 16488 7188
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 17052 7188 17080 7228
rect 21177 7225 21189 7228
rect 21223 7225 21235 7259
rect 21177 7219 21235 7225
rect 17313 7191 17371 7197
rect 17313 7188 17325 7191
rect 17052 7160 17325 7188
rect 17313 7157 17325 7160
rect 17359 7188 17371 7191
rect 17773 7191 17831 7197
rect 17773 7188 17785 7191
rect 17359 7160 17785 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 17773 7157 17785 7160
rect 17819 7157 17831 7191
rect 18230 7188 18236 7200
rect 18191 7160 18236 7188
rect 17773 7151 17831 7157
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 19702 7188 19708 7200
rect 19663 7160 19708 7188
rect 19702 7148 19708 7160
rect 19760 7148 19766 7200
rect 20070 7188 20076 7200
rect 20031 7160 20076 7188
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2777 6987 2835 6993
rect 2777 6984 2789 6987
rect 2004 6956 2789 6984
rect 2004 6944 2010 6956
rect 2777 6953 2789 6956
rect 2823 6984 2835 6987
rect 2869 6987 2927 6993
rect 2869 6984 2881 6987
rect 2823 6956 2881 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 2869 6953 2881 6956
rect 2915 6953 2927 6987
rect 2869 6947 2927 6953
rect 2961 6987 3019 6993
rect 2961 6953 2973 6987
rect 3007 6984 3019 6987
rect 3145 6987 3203 6993
rect 3145 6984 3157 6987
rect 3007 6956 3157 6984
rect 3007 6953 3019 6956
rect 2961 6947 3019 6953
rect 3145 6953 3157 6956
rect 3191 6984 3203 6987
rect 3786 6984 3792 6996
rect 3191 6956 3792 6984
rect 3191 6953 3203 6956
rect 3145 6947 3203 6953
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 6641 6987 6699 6993
rect 6641 6984 6653 6987
rect 4120 6956 6653 6984
rect 4120 6944 4126 6956
rect 6641 6953 6653 6956
rect 6687 6984 6699 6987
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 6687 6956 7573 6984
rect 6687 6953 6699 6956
rect 6641 6947 6699 6953
rect 7561 6953 7573 6956
rect 7607 6953 7619 6987
rect 7561 6947 7619 6953
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6984 8539 6987
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8527 6956 9045 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 9033 6953 9045 6956
rect 9079 6984 9091 6987
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9079 6956 9413 6984
rect 9079 6953 9091 6956
rect 9033 6947 9091 6953
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9401 6947 9459 6953
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10505 6987 10563 6993
rect 10505 6984 10517 6987
rect 10008 6956 10517 6984
rect 10008 6944 10014 6956
rect 10505 6953 10517 6956
rect 10551 6984 10563 6987
rect 10962 6984 10968 6996
rect 10551 6956 10968 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11606 6944 11612 6996
rect 11664 6984 11670 6996
rect 11790 6984 11796 6996
rect 11664 6956 11796 6984
rect 11664 6944 11670 6956
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 11882 6944 11888 6996
rect 11940 6984 11946 6996
rect 17218 6984 17224 6996
rect 11940 6956 17224 6984
rect 11940 6944 11946 6956
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17310 6944 17316 6996
rect 17368 6984 17374 6996
rect 17773 6987 17831 6993
rect 17773 6984 17785 6987
rect 17368 6956 17785 6984
rect 17368 6944 17374 6956
rect 17773 6953 17785 6956
rect 17819 6984 17831 6987
rect 17862 6984 17868 6996
rect 17819 6956 17868 6984
rect 17819 6953 17831 6956
rect 17773 6947 17831 6953
rect 17862 6944 17868 6956
rect 17920 6984 17926 6996
rect 18141 6987 18199 6993
rect 18141 6984 18153 6987
rect 17920 6956 18153 6984
rect 17920 6944 17926 6956
rect 18141 6953 18153 6956
rect 18187 6984 18199 6987
rect 18230 6984 18236 6996
rect 18187 6956 18236 6984
rect 18187 6953 18199 6956
rect 18141 6947 18199 6953
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 1664 6919 1722 6925
rect 1664 6885 1676 6919
rect 1710 6916 1722 6919
rect 3510 6916 3516 6928
rect 1710 6888 3516 6916
rect 1710 6885 1722 6888
rect 1664 6879 1722 6885
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 11149 6919 11207 6925
rect 11149 6916 11161 6919
rect 4028 6888 11161 6916
rect 4028 6876 4034 6888
rect 11149 6885 11161 6888
rect 11195 6916 11207 6919
rect 11238 6916 11244 6928
rect 11195 6888 11244 6916
rect 11195 6885 11207 6888
rect 11149 6879 11207 6885
rect 11238 6876 11244 6888
rect 11296 6876 11302 6928
rect 11440 6888 12388 6916
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 3421 6851 3479 6857
rect 3421 6848 3433 6851
rect 2004 6820 3433 6848
rect 2004 6808 2010 6820
rect 3421 6817 3433 6820
rect 3467 6848 3479 6851
rect 3881 6851 3939 6857
rect 3881 6848 3893 6851
rect 3467 6820 3893 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 3881 6817 3893 6820
rect 3927 6848 3939 6851
rect 4062 6848 4068 6860
rect 3927 6820 4068 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4430 6848 4436 6860
rect 4391 6820 4436 6848
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 4798 6848 4804 6860
rect 4571 6820 4804 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 5307 6820 6193 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 6181 6817 6193 6820
rect 6227 6848 6239 6851
rect 6822 6848 6828 6860
rect 6227 6820 6828 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7524 6820 7665 6848
rect 7524 6808 7530 6820
rect 7653 6817 7665 6820
rect 7699 6848 7711 6851
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7699 6820 8217 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 8938 6848 8944 6860
rect 8899 6820 8944 6848
rect 8205 6811 8263 6817
rect 8938 6808 8944 6820
rect 8996 6848 9002 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 8996 6820 9689 6848
rect 8996 6808 9002 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10134 6848 10140 6860
rect 9916 6820 10140 6848
rect 9916 6808 9922 6820
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 11440 6848 11468 6888
rect 11606 6857 11612 6860
rect 11600 6848 11612 6857
rect 10735 6820 11468 6848
rect 11567 6820 11612 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 11600 6811 11612 6820
rect 11606 6808 11612 6811
rect 11664 6808 11670 6860
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 4706 6780 4712 6792
rect 2915 6752 4712 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5537 6783 5595 6789
rect 5537 6780 5549 6783
rect 5408 6752 5549 6780
rect 5408 6740 5414 6752
rect 5537 6749 5549 6752
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7742 6780 7748 6792
rect 6972 6752 7748 6780
rect 6972 6740 6978 6752
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 9088 6752 9137 6780
rect 9088 6740 9094 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9364 6752 10548 6780
rect 9364 6740 9370 6752
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2464 6684 2973 6712
rect 2464 6672 2470 6684
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 3936 6684 4077 6712
rect 3936 6672 3942 6684
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 5077 6715 5135 6721
rect 5077 6681 5089 6715
rect 5123 6712 5135 6715
rect 5166 6712 5172 6724
rect 5123 6684 5172 6712
rect 5123 6681 5135 6684
rect 5077 6675 5135 6681
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 6638 6712 6644 6724
rect 5776 6684 6644 6712
rect 5776 6672 5782 6684
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 7193 6715 7251 6721
rect 7193 6681 7205 6715
rect 7239 6712 7251 6715
rect 8481 6715 8539 6721
rect 8481 6712 8493 6715
rect 7239 6684 8493 6712
rect 7239 6681 7251 6684
rect 7193 6675 7251 6681
rect 8481 6681 8493 6684
rect 8527 6681 8539 6715
rect 8481 6675 8539 6681
rect 9401 6715 9459 6721
rect 9401 6681 9413 6715
rect 9447 6712 9459 6715
rect 10410 6712 10416 6724
rect 9447 6684 10416 6712
rect 9447 6681 9459 6684
rect 9401 6675 9459 6681
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 2866 6644 2872 6656
rect 2740 6616 2872 6644
rect 2740 6604 2746 6616
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 5997 6647 6055 6653
rect 5997 6644 6009 6647
rect 5868 6616 6009 6644
rect 5868 6604 5874 6616
rect 5997 6613 6009 6616
rect 6043 6613 6055 6647
rect 7006 6644 7012 6656
rect 6967 6616 7012 6644
rect 5997 6607 6055 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 8202 6644 8208 6656
rect 7432 6616 8208 6644
rect 7432 6604 7438 6616
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8570 6644 8576 6656
rect 8531 6616 8576 6644
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 10134 6644 10140 6656
rect 10095 6616 10140 6644
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10520 6644 10548 6752
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 11020 6752 11345 6780
rect 11020 6740 11026 6752
rect 11333 6749 11345 6752
rect 11379 6749 11391 6783
rect 12360 6780 12388 6888
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 15194 6916 15200 6928
rect 12584 6888 15200 6916
rect 12584 6876 12590 6888
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13188 6857 13216 6888
rect 15194 6876 15200 6888
rect 15252 6876 15258 6928
rect 15562 6876 15568 6928
rect 15620 6916 15626 6928
rect 16022 6916 16028 6928
rect 15620 6888 16028 6916
rect 15620 6876 15626 6888
rect 16022 6876 16028 6888
rect 16080 6876 16086 6928
rect 16224 6888 16988 6916
rect 13173 6851 13231 6857
rect 12492 6820 13124 6848
rect 12492 6808 12498 6820
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 12360 6752 12817 6780
rect 11333 6743 11391 6749
rect 12805 6749 12817 6752
rect 12851 6749 12863 6783
rect 13096 6780 13124 6820
rect 13173 6817 13185 6851
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13538 6848 13544 6860
rect 13495 6820 13544 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13464 6780 13492 6811
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 13716 6851 13774 6857
rect 13716 6817 13728 6851
rect 13762 6848 13774 6851
rect 13998 6848 14004 6860
rect 13762 6820 14004 6848
rect 13762 6817 13774 6820
rect 13716 6811 13774 6817
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 14148 6820 15301 6848
rect 14148 6808 14154 6820
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 15841 6851 15899 6857
rect 15841 6848 15853 6851
rect 15335 6820 15853 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15841 6817 15853 6820
rect 15887 6817 15899 6851
rect 16224 6848 16252 6888
rect 15841 6811 15899 6817
rect 15948 6820 16252 6848
rect 16292 6851 16350 6857
rect 15470 6780 15476 6792
rect 13096 6752 13492 6780
rect 15431 6752 15476 6780
rect 12805 6743 12863 6749
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 12526 6672 12532 6724
rect 12584 6712 12590 6724
rect 15948 6712 15976 6820
rect 16292 6817 16304 6851
rect 16338 6848 16350 6851
rect 16850 6848 16856 6860
rect 16338 6820 16856 6848
rect 16338 6817 16350 6820
rect 16292 6811 16350 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 16960 6848 16988 6888
rect 18690 6848 18696 6860
rect 16960 6820 18696 6848
rect 18690 6808 18696 6820
rect 18748 6848 18754 6860
rect 18785 6851 18843 6857
rect 18785 6848 18797 6851
rect 18748 6820 18797 6848
rect 18748 6808 18754 6820
rect 18785 6817 18797 6820
rect 18831 6817 18843 6851
rect 18785 6811 18843 6817
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 18932 6820 20269 6848
rect 18932 6808 18938 6820
rect 20257 6817 20269 6820
rect 20303 6817 20315 6851
rect 20257 6811 20315 6817
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 18414 6780 18420 6792
rect 16080 6752 16125 6780
rect 18375 6752 18420 6780
rect 16080 6740 16086 6752
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 19334 6780 19340 6792
rect 19208 6752 19340 6780
rect 19208 6740 19214 6752
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 20717 6783 20775 6789
rect 20717 6749 20729 6783
rect 20763 6780 20775 6783
rect 20806 6780 20812 6792
rect 20763 6752 20812 6780
rect 20763 6749 20775 6752
rect 20717 6743 20775 6749
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 12584 6684 13492 6712
rect 12584 6672 12590 6684
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 10520 6616 12725 6644
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 12805 6647 12863 6653
rect 12805 6613 12817 6647
rect 12851 6644 12863 6647
rect 12989 6647 13047 6653
rect 12989 6644 13001 6647
rect 12851 6616 13001 6644
rect 12851 6613 12863 6616
rect 12805 6607 12863 6613
rect 12989 6613 13001 6616
rect 13035 6644 13047 6647
rect 13078 6644 13084 6656
rect 13035 6616 13084 6644
rect 13035 6613 13047 6616
rect 12989 6607 13047 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13464 6644 13492 6684
rect 14476 6684 15976 6712
rect 16951 6684 17632 6712
rect 14476 6644 14504 6684
rect 13464 6616 14504 6644
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14829 6647 14887 6653
rect 14829 6644 14841 6647
rect 14608 6616 14841 6644
rect 14608 6604 14614 6616
rect 14829 6613 14841 6616
rect 14875 6613 14887 6647
rect 14829 6607 14887 6613
rect 15841 6647 15899 6653
rect 15841 6613 15853 6647
rect 15887 6644 15899 6647
rect 16951 6644 16979 6684
rect 15887 6616 16979 6644
rect 17405 6647 17463 6653
rect 15887 6613 15899 6616
rect 15841 6607 15899 6613
rect 17405 6613 17417 6647
rect 17451 6644 17463 6647
rect 17494 6644 17500 6656
rect 17451 6616 17500 6644
rect 17451 6613 17463 6616
rect 17405 6607 17463 6613
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 17604 6644 17632 6684
rect 18506 6672 18512 6724
rect 18564 6712 18570 6724
rect 19889 6715 19947 6721
rect 19889 6712 19901 6715
rect 18564 6684 19901 6712
rect 18564 6672 18570 6684
rect 19889 6681 19901 6684
rect 19935 6681 19947 6715
rect 19889 6675 19947 6681
rect 18598 6644 18604 6656
rect 17604 6616 18604 6644
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 19150 6644 19156 6656
rect 19111 6616 19156 6644
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19518 6644 19524 6656
rect 19479 6616 19524 6644
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 20162 6604 20168 6656
rect 20220 6644 20226 6656
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 20220 6616 21097 6644
rect 20220 6604 20226 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 2406 6440 2412 6452
rect 1719 6412 2412 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 3510 6400 3516 6452
rect 3568 6440 3574 6452
rect 3605 6443 3663 6449
rect 3605 6440 3617 6443
rect 3568 6412 3617 6440
rect 3568 6400 3574 6412
rect 3605 6409 3617 6412
rect 3651 6409 3663 6443
rect 3605 6403 3663 6409
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 13446 6440 13452 6452
rect 4120 6412 13452 6440
rect 4120 6400 4126 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 19150 6440 19156 6452
rect 13556 6412 19156 6440
rect 5166 6332 5172 6384
rect 5224 6372 5230 6384
rect 5537 6375 5595 6381
rect 5537 6372 5549 6375
rect 5224 6344 5549 6372
rect 5224 6332 5230 6344
rect 5537 6341 5549 6344
rect 5583 6372 5595 6375
rect 5583 6344 7512 6372
rect 5583 6341 5595 6344
rect 5537 6335 5595 6341
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6914 6304 6920 6316
rect 6227 6276 6920 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7156 6276 7389 6304
rect 7156 6264 7162 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7484 6304 7512 6344
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 10042 6372 10048 6384
rect 9456 6344 10048 6372
rect 9456 6332 9462 6344
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 11701 6375 11759 6381
rect 11701 6341 11713 6375
rect 11747 6341 11759 6375
rect 11701 6335 11759 6341
rect 7484 6276 8432 6304
rect 7377 6267 7435 6273
rect 1394 6196 1400 6248
rect 1452 6236 1458 6248
rect 1854 6236 1860 6248
rect 1452 6208 1860 6236
rect 1452 6196 1458 6208
rect 1854 6196 1860 6208
rect 1912 6236 1918 6248
rect 2225 6239 2283 6245
rect 2225 6236 2237 6239
rect 1912 6208 2237 6236
rect 1912 6196 1918 6208
rect 2225 6205 2237 6208
rect 2271 6236 2283 6239
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 2271 6208 4169 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 4157 6205 4169 6208
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4424 6239 4482 6245
rect 4424 6205 4436 6239
rect 4470 6236 4482 6239
rect 5258 6236 5264 6248
rect 4470 6208 5264 6236
rect 4470 6205 4482 6208
rect 4424 6199 4482 6205
rect 2492 6171 2550 6177
rect 2492 6137 2504 6171
rect 2538 6168 2550 6171
rect 3142 6168 3148 6180
rect 2538 6140 3148 6168
rect 2538 6137 2550 6140
rect 2492 6131 2550 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 4172 6168 4200 6199
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 5626 6236 5632 6248
rect 5539 6208 5632 6236
rect 5552 6168 5580 6208
rect 5626 6196 5632 6208
rect 5684 6236 5690 6248
rect 5810 6236 5816 6248
rect 5684 6208 5816 6236
rect 5684 6196 5690 6208
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 6273 6239 6331 6245
rect 6273 6205 6285 6239
rect 6319 6236 6331 6239
rect 7190 6236 7196 6248
rect 6319 6208 7196 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6205 8355 6239
rect 8404 6236 8432 6276
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 9950 6304 9956 6316
rect 9640 6276 9956 6304
rect 9640 6264 9646 6276
rect 9950 6264 9956 6276
rect 10008 6304 10014 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 10008 6276 10333 6304
rect 10008 6264 10014 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 8404 6208 10241 6236
rect 8297 6199 8355 6205
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 7006 6168 7012 6180
rect 4172 6140 5580 6168
rect 5644 6140 7012 6168
rect 3970 6100 3976 6112
rect 3931 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 5644 6100 5672 6140
rect 7006 6128 7012 6140
rect 7064 6168 7070 6180
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 7064 6140 7297 6168
rect 7064 6128 7070 6140
rect 7285 6137 7297 6140
rect 7331 6137 7343 6171
rect 7285 6131 7343 6137
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 7742 6168 7748 6180
rect 7432 6140 7748 6168
rect 7432 6128 7438 6140
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 4120 6072 5672 6100
rect 4120 6060 4126 6072
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6822 6100 6828 6112
rect 6420 6072 6828 6100
rect 6420 6060 6426 6072
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7466 6100 7472 6112
rect 6972 6072 7472 6100
rect 6972 6060 6978 6072
rect 7466 6060 7472 6072
rect 7524 6100 7530 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7524 6072 7849 6100
rect 7524 6060 7530 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 8312 6100 8340 6199
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 11716 6236 11744 6335
rect 12434 6304 12440 6316
rect 12395 6276 12440 6304
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 12526 6236 12532 6248
rect 10468 6208 11376 6236
rect 11716 6208 12532 6236
rect 10468 6196 10474 6208
rect 8564 6171 8622 6177
rect 8564 6137 8576 6171
rect 8610 6168 8622 6171
rect 8662 6168 8668 6180
rect 8610 6140 8668 6168
rect 8610 6137 8622 6140
rect 8564 6131 8622 6137
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 10566 6171 10624 6177
rect 10566 6168 10578 6171
rect 9692 6140 10578 6168
rect 9214 6100 9220 6112
rect 8312 6072 9220 6100
rect 7837 6063 7895 6069
rect 9214 6060 9220 6072
rect 9272 6100 9278 6112
rect 9582 6100 9588 6112
rect 9272 6072 9588 6100
rect 9272 6060 9278 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9692 6109 9720 6140
rect 10566 6137 10578 6140
rect 10612 6168 10624 6171
rect 11238 6168 11244 6180
rect 10612 6140 11244 6168
rect 10612 6137 10624 6140
rect 10566 6131 10624 6137
rect 11238 6128 11244 6140
rect 11296 6128 11302 6180
rect 11348 6168 11376 6208
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 13556 6236 13584 6412
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19334 6440 19340 6452
rect 19295 6412 19340 6440
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 13817 6375 13875 6381
rect 13817 6341 13829 6375
rect 13863 6341 13875 6375
rect 16209 6375 16267 6381
rect 16209 6372 16221 6375
rect 13817 6335 13875 6341
rect 15672 6344 16221 6372
rect 13832 6304 13860 6335
rect 13998 6304 14004 6316
rect 13832 6276 14004 6304
rect 13998 6264 14004 6276
rect 14056 6304 14062 6316
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 14056 6276 14749 6304
rect 14056 6264 14062 6276
rect 14737 6273 14749 6276
rect 14783 6304 14795 6307
rect 15010 6304 15016 6316
rect 14783 6276 15016 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15672 6313 15700 6344
rect 16209 6341 16221 6344
rect 16255 6372 16267 6375
rect 20809 6375 20867 6381
rect 20809 6372 20821 6375
rect 16255 6344 20821 6372
rect 16255 6341 16267 6344
rect 16209 6335 16267 6341
rect 20809 6341 20821 6344
rect 20855 6341 20867 6375
rect 20809 6335 20867 6341
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6273 15715 6307
rect 15838 6304 15844 6316
rect 15751 6276 15844 6304
rect 15657 6267 15715 6273
rect 15838 6264 15844 6276
rect 15896 6304 15902 6316
rect 16850 6304 16856 6316
rect 15896 6276 16712 6304
rect 16763 6276 16856 6304
rect 15896 6264 15902 6276
rect 12636 6208 13584 6236
rect 12636 6168 12664 6208
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 15378 6236 15384 6248
rect 13780 6208 15384 6236
rect 13780 6196 13786 6208
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6236 15623 6239
rect 16390 6236 16396 6248
rect 15611 6208 16396 6236
rect 15611 6205 15623 6208
rect 15565 6199 15623 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 16577 6239 16635 6245
rect 16577 6236 16589 6239
rect 16540 6208 16589 6236
rect 16540 6196 16546 6208
rect 16577 6205 16589 6208
rect 16623 6205 16635 6239
rect 16684 6236 16712 6276
rect 16850 6264 16856 6276
rect 16908 6304 16914 6316
rect 17310 6304 17316 6316
rect 16908 6276 17316 6304
rect 16908 6264 16914 6276
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17552 6276 18245 6304
rect 17552 6264 17558 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 18656 6276 19717 6304
rect 18656 6264 18662 6276
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 17512 6236 17540 6264
rect 16684 6208 17540 6236
rect 16577 6199 16635 6205
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 17736 6208 18797 6236
rect 17736 6196 17742 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 18932 6208 20085 6236
rect 18932 6196 18938 6208
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 20073 6199 20131 6205
rect 12710 6177 12716 6180
rect 11348 6140 12664 6168
rect 12704 6131 12716 6177
rect 12768 6168 12774 6180
rect 12986 6168 12992 6180
rect 12768 6140 12992 6168
rect 12710 6128 12716 6131
rect 12768 6128 12774 6140
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 14274 6128 14280 6180
rect 14332 6168 14338 6180
rect 14461 6171 14519 6177
rect 14461 6168 14473 6171
rect 14332 6140 14473 6168
rect 14332 6128 14338 6140
rect 14461 6137 14473 6140
rect 14507 6168 14519 6171
rect 15930 6168 15936 6180
rect 14507 6140 15936 6168
rect 14507 6137 14519 6140
rect 14461 6131 14519 6137
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 16850 6168 16856 6180
rect 16592 6140 16856 6168
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6069 9735 6103
rect 9677 6063 9735 6069
rect 10229 6103 10287 6109
rect 10229 6069 10241 6103
rect 10275 6100 10287 6103
rect 11882 6100 11888 6112
rect 10275 6072 11888 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12158 6100 12164 6112
rect 12115 6072 12164 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 14090 6100 14096 6112
rect 14051 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 15102 6100 15108 6112
rect 14599 6072 15108 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 16592 6100 16620 6140
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 16951 6140 17724 6168
rect 15243 6072 16620 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 16951 6100 16979 6140
rect 17696 6112 17724 6140
rect 18046 6128 18052 6180
rect 18104 6168 18110 6180
rect 20441 6171 20499 6177
rect 20441 6168 20453 6171
rect 18104 6140 20453 6168
rect 18104 6128 18110 6140
rect 20441 6137 20453 6140
rect 20487 6137 20499 6171
rect 20441 6131 20499 6137
rect 16724 6072 16979 6100
rect 17313 6103 17371 6109
rect 16724 6060 16730 6072
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 17494 6100 17500 6112
rect 17359 6072 17500 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 17678 6100 17684 6112
rect 17639 6072 17684 6100
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18601 6103 18659 6109
rect 18601 6100 18613 6103
rect 17828 6072 18613 6100
rect 17828 6060 17834 6072
rect 18601 6069 18613 6072
rect 18647 6069 18659 6103
rect 18601 6063 18659 6069
rect 18785 6103 18843 6109
rect 18785 6069 18797 6103
rect 18831 6100 18843 6103
rect 18969 6103 19027 6109
rect 18969 6100 18981 6103
rect 18831 6072 18981 6100
rect 18831 6069 18843 6072
rect 18785 6063 18843 6069
rect 18969 6069 18981 6072
rect 19015 6069 19027 6103
rect 21174 6100 21180 6112
rect 21135 6072 21180 6100
rect 18969 6063 19027 6069
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2498 5896 2504 5908
rect 2455 5868 2504 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3970 5896 3976 5908
rect 3559 5868 3976 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3970 5856 3976 5868
rect 4028 5896 4034 5908
rect 6546 5896 6552 5908
rect 4028 5868 6552 5896
rect 4028 5856 4034 5868
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7098 5896 7104 5908
rect 6963 5868 7104 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 8938 5896 8944 5908
rect 8899 5868 8944 5896
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9766 5896 9772 5908
rect 9539 5868 9772 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 11057 5899 11115 5905
rect 9876 5868 10171 5896
rect 3878 5788 3884 5840
rect 3936 5828 3942 5840
rect 5445 5831 5503 5837
rect 3936 5800 5396 5828
rect 3936 5788 3942 5800
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 3050 5760 3056 5772
rect 2832 5732 3056 5760
rect 2832 5720 2838 5732
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4304 5732 4445 5760
rect 4304 5720 4310 5732
rect 4433 5729 4445 5732
rect 4479 5760 4491 5763
rect 4890 5760 4896 5772
rect 4479 5732 4896 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 2866 5692 2872 5704
rect 2372 5664 2872 5692
rect 2372 5652 2378 5664
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 2406 5584 2412 5636
rect 2464 5624 2470 5636
rect 2976 5624 3004 5655
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 4062 5692 4068 5704
rect 3384 5664 4068 5692
rect 3384 5652 3390 5664
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4212 5664 4537 5692
rect 4212 5652 4218 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4706 5692 4712 5704
rect 4619 5664 4712 5692
rect 4525 5655 4583 5661
rect 4706 5652 4712 5664
rect 4764 5692 4770 5704
rect 5166 5692 5172 5704
rect 4764 5664 5172 5692
rect 4764 5652 4770 5664
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 3142 5624 3148 5636
rect 2464 5596 2636 5624
rect 2976 5596 3148 5624
rect 2464 5584 2470 5596
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 2498 5556 2504 5568
rect 2363 5528 2504 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 2608 5556 2636 5596
rect 3142 5584 3148 5596
rect 3200 5624 3206 5636
rect 4724 5624 4752 5652
rect 3200 5596 4752 5624
rect 3200 5584 3206 5596
rect 3602 5556 3608 5568
rect 2608 5528 3608 5556
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 5368 5556 5396 5800
rect 5445 5797 5457 5831
rect 5491 5828 5503 5831
rect 7282 5828 7288 5840
rect 5491 5800 7288 5828
rect 5491 5797 5503 5800
rect 5445 5791 5503 5797
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 8386 5828 8392 5840
rect 7576 5800 8392 5828
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 5626 5760 5632 5772
rect 5583 5732 5632 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 5804 5763 5862 5769
rect 5804 5729 5816 5763
rect 5850 5760 5862 5763
rect 6086 5760 6092 5772
rect 5850 5732 6092 5760
rect 5850 5729 5862 5732
rect 5804 5723 5862 5729
rect 6086 5720 6092 5732
rect 6144 5760 6150 5772
rect 6914 5760 6920 5772
rect 6144 5732 6920 5760
rect 6144 5720 6150 5732
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7098 5720 7104 5772
rect 7156 5760 7162 5772
rect 7449 5763 7507 5769
rect 7449 5760 7461 5763
rect 7156 5732 7461 5760
rect 7156 5720 7162 5732
rect 7449 5729 7461 5732
rect 7495 5760 7507 5763
rect 7576 5760 7604 5800
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 8570 5788 8576 5840
rect 8628 5828 8634 5840
rect 9876 5828 9904 5868
rect 10045 5831 10103 5837
rect 10045 5828 10057 5831
rect 8628 5800 9904 5828
rect 9968 5800 10057 5828
rect 8628 5788 8634 5800
rect 9968 5772 9996 5800
rect 10045 5797 10057 5800
rect 10091 5797 10103 5831
rect 10143 5828 10171 5868
rect 11057 5865 11069 5899
rect 11103 5896 11115 5899
rect 11146 5896 11152 5908
rect 11103 5868 11152 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 12802 5896 12808 5908
rect 11296 5868 12808 5896
rect 11296 5856 11302 5868
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 12986 5896 12992 5908
rect 12947 5868 12992 5896
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13630 5896 13636 5908
rect 13320 5868 13636 5896
rect 13320 5856 13326 5868
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 14056 5868 14105 5896
rect 14056 5856 14062 5868
rect 14093 5865 14105 5868
rect 14139 5896 14151 5899
rect 19429 5899 19487 5905
rect 19429 5896 19441 5899
rect 14139 5868 19441 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 19429 5865 19441 5868
rect 19475 5865 19487 5899
rect 19429 5859 19487 5865
rect 11609 5831 11667 5837
rect 11609 5828 11621 5831
rect 10143 5800 11621 5828
rect 10045 5791 10103 5797
rect 11609 5797 11621 5800
rect 11655 5797 11667 5831
rect 11790 5828 11796 5840
rect 11751 5800 11796 5828
rect 11609 5791 11667 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 12345 5831 12403 5837
rect 12345 5797 12357 5831
rect 12391 5828 12403 5831
rect 12710 5828 12716 5840
rect 12391 5800 12716 5828
rect 12391 5797 12403 5800
rect 12345 5791 12403 5797
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 13078 5788 13084 5840
rect 13136 5828 13142 5840
rect 13136 5800 14596 5828
rect 13136 5788 13142 5800
rect 7495 5732 7604 5760
rect 7495 5729 7507 5732
rect 7449 5723 7507 5729
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 9766 5760 9772 5772
rect 7800 5732 9772 5760
rect 7800 5720 7806 5732
rect 9766 5720 9772 5732
rect 9824 5760 9830 5772
rect 9824 5732 9904 5760
rect 9824 5720 9830 5732
rect 7190 5692 7196 5704
rect 7151 5664 7196 5692
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 9674 5692 9680 5704
rect 8352 5664 9680 5692
rect 8352 5652 8358 5664
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 9876 5692 9904 5732
rect 9950 5720 9956 5772
rect 10008 5720 10014 5772
rect 10060 5732 10364 5760
rect 10060 5692 10088 5732
rect 10336 5701 10364 5732
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 11149 5763 11207 5769
rect 11149 5760 11161 5763
rect 10468 5732 11161 5760
rect 10468 5720 10474 5732
rect 11149 5729 11161 5732
rect 11195 5760 11207 5763
rect 11808 5760 11836 5788
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 11195 5732 11836 5760
rect 11900 5732 13369 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 9876 5664 10088 5692
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10502 5692 10508 5704
rect 10367 5664 10508 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 9493 5627 9551 5633
rect 9493 5624 9505 5627
rect 8496 5596 9505 5624
rect 8496 5556 8524 5596
rect 9493 5593 9505 5596
rect 9539 5593 9551 5627
rect 9493 5587 9551 5593
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10152 5624 10180 5655
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 11238 5692 11244 5704
rect 11199 5664 11244 5692
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5692 11667 5695
rect 11900 5692 11928 5732
rect 13357 5729 13369 5732
rect 13403 5760 13415 5763
rect 13538 5760 13544 5772
rect 13403 5732 13544 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 14458 5760 14464 5772
rect 14419 5732 14464 5760
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 14568 5760 14596 5800
rect 15010 5788 15016 5840
rect 15068 5828 15074 5840
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 15068 5800 16313 5828
rect 15068 5788 15074 5800
rect 16301 5797 16313 5800
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 16574 5788 16580 5840
rect 16632 5828 16638 5840
rect 17494 5828 17500 5840
rect 16632 5800 17500 5828
rect 16632 5788 16638 5800
rect 17494 5788 17500 5800
rect 17552 5788 17558 5840
rect 17770 5788 17776 5840
rect 17828 5828 17834 5840
rect 18325 5831 18383 5837
rect 18325 5828 18337 5831
rect 17828 5800 18337 5828
rect 17828 5788 17834 5800
rect 18325 5797 18337 5800
rect 18371 5797 18383 5831
rect 18690 5828 18696 5840
rect 18651 5800 18696 5828
rect 18325 5791 18383 5797
rect 18690 5788 18696 5800
rect 18748 5828 18754 5840
rect 19061 5831 19119 5837
rect 19061 5828 19073 5831
rect 18748 5800 19073 5828
rect 18748 5788 18754 5800
rect 19061 5797 19073 5800
rect 19107 5797 19119 5831
rect 19061 5791 19119 5797
rect 15654 5760 15660 5772
rect 14568 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 16540 5732 16681 5760
rect 16540 5720 16546 5732
rect 16669 5729 16681 5732
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 16936 5763 16994 5769
rect 16936 5729 16948 5763
rect 16982 5760 16994 5763
rect 17402 5760 17408 5772
rect 16982 5732 17408 5760
rect 16982 5729 16994 5732
rect 16936 5723 16994 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 17678 5720 17684 5772
rect 17736 5760 17742 5772
rect 19518 5760 19524 5772
rect 17736 5732 19524 5760
rect 17736 5720 17742 5732
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 11655 5664 11928 5692
rect 12437 5695 12495 5701
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5692 12679 5695
rect 12986 5692 12992 5704
rect 12667 5664 12992 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 10100 5596 10180 5624
rect 10689 5627 10747 5633
rect 10100 5584 10106 5596
rect 10689 5593 10701 5627
rect 10735 5624 10747 5627
rect 12452 5624 12480 5655
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5692 13691 5695
rect 13722 5692 13728 5704
rect 13679 5664 13728 5692
rect 13679 5661 13691 5664
rect 13633 5655 13691 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 14090 5652 14096 5704
rect 14148 5692 14154 5704
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14148 5664 14565 5692
rect 14148 5652 14154 5664
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 12894 5624 12900 5636
rect 10735 5596 12900 5624
rect 10735 5593 10747 5596
rect 10689 5587 10747 5593
rect 12894 5584 12900 5596
rect 12952 5584 12958 5636
rect 14568 5624 14596 5655
rect 14642 5652 14648 5704
rect 14700 5692 14706 5704
rect 14700 5664 14745 5692
rect 14700 5652 14706 5664
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 20533 5695 20591 5701
rect 20533 5692 20545 5695
rect 18932 5664 20545 5692
rect 18932 5652 18938 5664
rect 20533 5661 20545 5664
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 14568 5596 15608 5624
rect 5368 5528 8524 5556
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9306 5556 9312 5568
rect 8628 5528 8673 5556
rect 9267 5528 9312 5556
rect 8628 5516 8634 5528
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 11606 5556 11612 5568
rect 9723 5528 11612 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 11606 5516 11612 5528
rect 11664 5516 11670 5568
rect 11977 5559 12035 5565
rect 11977 5525 11989 5559
rect 12023 5556 12035 5559
rect 13262 5556 13268 5568
rect 12023 5528 13268 5556
rect 12023 5525 12035 5528
rect 11977 5519 12035 5525
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 15378 5516 15384 5568
rect 15436 5556 15442 5568
rect 15473 5559 15531 5565
rect 15473 5556 15485 5559
rect 15436 5528 15485 5556
rect 15436 5516 15442 5528
rect 15473 5525 15485 5528
rect 15519 5525 15531 5559
rect 15580 5556 15608 5596
rect 17862 5584 17868 5636
rect 17920 5624 17926 5636
rect 18049 5627 18107 5633
rect 18049 5624 18061 5627
rect 17920 5596 18061 5624
rect 17920 5584 17926 5596
rect 18049 5593 18061 5596
rect 18095 5593 18107 5627
rect 19334 5624 19340 5636
rect 18049 5587 18107 5593
rect 18156 5596 19340 5624
rect 18156 5556 18184 5596
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 20165 5627 20223 5633
rect 20165 5624 20177 5627
rect 19444 5596 20177 5624
rect 15580 5528 18184 5556
rect 15473 5519 15531 5525
rect 18598 5516 18604 5568
rect 18656 5556 18662 5568
rect 19444 5556 19472 5596
rect 20165 5593 20177 5596
rect 20211 5593 20223 5627
rect 20165 5587 20223 5593
rect 18656 5528 19472 5556
rect 18656 5516 18662 5528
rect 19518 5516 19524 5568
rect 19576 5556 19582 5568
rect 19797 5559 19855 5565
rect 19797 5556 19809 5559
rect 19576 5528 19809 5556
rect 19576 5516 19582 5528
rect 19797 5525 19809 5528
rect 19843 5525 19855 5559
rect 19797 5519 19855 5525
rect 19886 5516 19892 5568
rect 19944 5556 19950 5568
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 19944 5528 21097 5556
rect 19944 5516 19950 5528
rect 21085 5525 21097 5528
rect 21131 5525 21143 5559
rect 21085 5519 21143 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3789 5355 3847 5361
rect 3789 5352 3801 5355
rect 3476 5324 3801 5352
rect 3476 5312 3482 5324
rect 3789 5321 3801 5324
rect 3835 5321 3847 5355
rect 3789 5315 3847 5321
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5169 5355 5227 5361
rect 5169 5352 5181 5355
rect 4948 5324 5181 5352
rect 4948 5312 4954 5324
rect 5169 5321 5181 5324
rect 5215 5321 5227 5355
rect 7929 5355 7987 5361
rect 7929 5352 7941 5355
rect 5169 5315 5227 5321
rect 6288 5324 7941 5352
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4801 5287 4859 5293
rect 4801 5284 4813 5287
rect 4212 5256 4813 5284
rect 4212 5244 4218 5256
rect 4801 5253 4813 5256
rect 4847 5253 4859 5287
rect 6288 5284 6316 5324
rect 7929 5321 7941 5324
rect 7975 5321 7987 5355
rect 13814 5352 13820 5364
rect 7929 5315 7987 5321
rect 8496 5324 13820 5352
rect 4801 5247 4859 5253
rect 6196 5256 6316 5284
rect 7009 5287 7067 5293
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4706 5216 4712 5228
rect 4479 5188 4712 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 6196 5225 6224 5256
rect 7009 5253 7021 5287
rect 7055 5284 7067 5287
rect 8496 5284 8524 5324
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 14642 5352 14648 5364
rect 13955 5324 14648 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 15010 5312 15016 5364
rect 15068 5352 15074 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 15068 5324 15209 5352
rect 15068 5312 15074 5324
rect 15197 5321 15209 5324
rect 15243 5321 15255 5355
rect 17402 5352 17408 5364
rect 15197 5315 15255 5321
rect 15672 5324 17080 5352
rect 17363 5324 17408 5352
rect 7055 5256 8524 5284
rect 7055 5253 7067 5256
rect 7009 5247 7067 5253
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5185 6239 5219
rect 6181 5179 6239 5185
rect 6273 5219 6331 5225
rect 6273 5185 6285 5219
rect 6319 5216 6331 5219
rect 6638 5216 6644 5228
rect 6319 5188 6644 5216
rect 6319 5185 6331 5188
rect 6273 5179 6331 5185
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 6972 5188 7573 5216
rect 6972 5176 6978 5188
rect 7561 5185 7573 5188
rect 7607 5216 7619 5219
rect 7742 5216 7748 5228
rect 7607 5188 7748 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 8496 5225 8524 5256
rect 10873 5287 10931 5293
rect 10873 5253 10885 5287
rect 10919 5284 10931 5287
rect 10962 5284 10968 5296
rect 10919 5256 10968 5284
rect 10919 5253 10931 5256
rect 10873 5247 10931 5253
rect 10962 5244 10968 5256
rect 11020 5284 11026 5296
rect 11020 5256 15608 5284
rect 11020 5244 11026 5256
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 11606 5216 11612 5228
rect 11567 5188 11612 5216
rect 8573 5179 8631 5185
rect 5718 5148 5724 5160
rect 4172 5120 5724 5148
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5080 1915 5083
rect 2498 5080 2504 5092
rect 1903 5052 2504 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 2498 5040 2504 5052
rect 2556 5040 2562 5092
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 4172 5089 4200 5120
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6362 5148 6368 5160
rect 6135 5120 6368 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 8386 5108 8392 5160
rect 8444 5148 8450 5160
rect 8588 5148 8616 5179
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11808 5225 11836 5256
rect 15580 5228 15608 5256
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5185 11851 5219
rect 12710 5216 12716 5228
rect 11793 5179 11851 5185
rect 12544 5188 12716 5216
rect 8444 5120 8616 5148
rect 8849 5151 8907 5157
rect 8444 5108 8450 5120
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9493 5151 9551 5157
rect 8895 5120 9444 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 3605 5083 3663 5089
rect 3605 5080 3617 5083
rect 2648 5052 3617 5080
rect 2648 5040 2654 5052
rect 3605 5049 3617 5052
rect 3651 5080 3663 5083
rect 4157 5083 4215 5089
rect 4157 5080 4169 5083
rect 3651 5052 4169 5080
rect 3651 5049 3663 5052
rect 3605 5043 3663 5049
rect 4157 5049 4169 5052
rect 4203 5049 4215 5083
rect 4157 5043 4215 5049
rect 4890 5040 4896 5092
rect 4948 5080 4954 5092
rect 7006 5080 7012 5092
rect 4948 5052 7012 5080
rect 4948 5040 4954 5052
rect 7006 5040 7012 5052
rect 7064 5080 7070 5092
rect 7377 5083 7435 5089
rect 7377 5080 7389 5083
rect 7064 5052 7389 5080
rect 7064 5040 7070 5052
rect 7377 5049 7389 5052
rect 7423 5049 7435 5083
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 7377 5043 7435 5049
rect 7484 5052 9045 5080
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 2464 4984 2789 5012
rect 2464 4972 2470 4984
rect 2777 4981 2789 4984
rect 2823 5012 2835 5015
rect 2866 5012 2872 5024
rect 2823 4984 2872 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 3145 5015 3203 5021
rect 3145 5012 3157 5015
rect 3108 4984 3157 5012
rect 3108 4972 3114 4984
rect 3145 4981 3157 4984
rect 3191 4981 3203 5015
rect 3145 4975 3203 4981
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 4249 5015 4307 5021
rect 4249 5012 4261 5015
rect 4028 4984 4261 5012
rect 4028 4972 4034 4984
rect 4249 4981 4261 4984
rect 4295 4981 4307 5015
rect 4249 4975 4307 4981
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5408 4984 5549 5012
rect 5408 4972 5414 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 5537 4975 5595 4981
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 7098 5012 7104 5024
rect 5767 4984 7104 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 7484 5021 7512 5052
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9416 5080 9444 5120
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 9582 5148 9588 5160
rect 9539 5120 9588 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9766 5157 9772 5160
rect 9760 5148 9772 5157
rect 9727 5120 9772 5148
rect 9760 5111 9772 5120
rect 9766 5108 9772 5111
rect 9824 5108 9830 5160
rect 11624 5148 11652 5176
rect 12250 5148 12256 5160
rect 11624 5120 12256 5148
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12544 5148 12572 5188
rect 12710 5176 12716 5188
rect 12768 5216 12774 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12768 5188 12909 5216
rect 12768 5176 12774 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13004 5188 14136 5216
rect 12483 5120 12572 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 13004 5148 13032 5188
rect 13998 5148 14004 5160
rect 12676 5120 13032 5148
rect 13959 5120 14004 5148
rect 12676 5108 12682 5120
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 14108 5148 14136 5188
rect 14458 5176 14464 5228
rect 14516 5216 14522 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14516 5188 14749 5216
rect 14516 5176 14522 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 15562 5216 15568 5228
rect 15523 5188 15568 5216
rect 14737 5179 14795 5185
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 15672 5148 15700 5324
rect 17052 5216 17080 5324
rect 17402 5312 17408 5324
rect 17460 5352 17466 5364
rect 18233 5355 18291 5361
rect 18233 5352 18245 5355
rect 17460 5324 18245 5352
rect 17460 5312 17466 5324
rect 18233 5321 18245 5324
rect 18279 5321 18291 5355
rect 18233 5315 18291 5321
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 18969 5355 19027 5361
rect 18969 5352 18981 5355
rect 18748 5324 18981 5352
rect 18748 5312 18754 5324
rect 18969 5321 18981 5324
rect 19015 5321 19027 5355
rect 19334 5352 19340 5364
rect 19295 5324 19340 5352
rect 18969 5315 19027 5321
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 17126 5244 17132 5296
rect 17184 5284 17190 5296
rect 19705 5287 19763 5293
rect 19705 5284 19717 5287
rect 17184 5256 19717 5284
rect 17184 5244 17190 5256
rect 19705 5253 19717 5256
rect 19751 5253 19763 5287
rect 19705 5247 19763 5253
rect 20530 5216 20536 5228
rect 17052 5188 20536 5216
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 16022 5148 16028 5160
rect 14108 5120 15700 5148
rect 15983 5120 16028 5148
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 20441 5151 20499 5157
rect 20441 5148 20453 5151
rect 16132 5120 20453 5148
rect 9950 5080 9956 5092
rect 9416 5052 9956 5080
rect 9033 5043 9091 5049
rect 7469 5015 7527 5021
rect 7469 5012 7481 5015
rect 7340 4984 7481 5012
rect 7340 4972 7346 4984
rect 7469 4981 7481 4984
rect 7515 4981 7527 5015
rect 7469 4975 7527 4981
rect 7929 5015 7987 5021
rect 7929 4981 7941 5015
rect 7975 5012 7987 5015
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7975 4984 8033 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8021 4981 8033 4984
rect 8067 5012 8079 5015
rect 8202 5012 8208 5024
rect 8067 4984 8208 5012
rect 8067 4981 8079 4984
rect 8021 4975 8079 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8386 5012 8392 5024
rect 8299 4984 8392 5012
rect 8386 4972 8392 4984
rect 8444 5012 8450 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 8444 4984 8861 5012
rect 8444 4972 8450 4984
rect 8849 4981 8861 4984
rect 8895 4981 8907 5015
rect 9048 5012 9076 5043
rect 9950 5040 9956 5052
rect 10008 5040 10014 5092
rect 10502 5040 10508 5092
rect 10560 5080 10566 5092
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 10560 5052 11529 5080
rect 10560 5040 10566 5052
rect 11517 5049 11529 5052
rect 11563 5080 11575 5083
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 11563 5052 13277 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 13265 5049 13277 5052
rect 13311 5049 13323 5083
rect 14277 5083 14335 5089
rect 13265 5043 13323 5049
rect 13740 5052 13952 5080
rect 10778 5012 10784 5024
rect 9048 4984 10784 5012
rect 8849 4975 8907 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11146 5012 11152 5024
rect 11107 4984 11152 5012
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 11296 4984 12173 5012
rect 11296 4972 11302 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12161 4975 12219 4981
rect 12250 4972 12256 5024
rect 12308 5012 12314 5024
rect 13740 5012 13768 5052
rect 12308 4984 13768 5012
rect 13924 5012 13952 5052
rect 14277 5049 14289 5083
rect 14323 5080 14335 5083
rect 14366 5080 14372 5092
rect 14323 5052 14372 5080
rect 14323 5049 14335 5052
rect 14277 5043 14335 5049
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 16132 5080 16160 5120
rect 20441 5117 20453 5120
rect 20487 5117 20499 5151
rect 20441 5111 20499 5117
rect 15120 5052 16160 5080
rect 16292 5083 16350 5089
rect 15120 5012 15148 5052
rect 16292 5049 16304 5083
rect 16338 5080 16350 5083
rect 16850 5080 16856 5092
rect 16338 5052 16856 5080
rect 16338 5049 16350 5052
rect 16292 5043 16350 5049
rect 16850 5040 16856 5052
rect 16908 5040 16914 5092
rect 20809 5083 20867 5089
rect 20809 5080 20821 5083
rect 16960 5052 20821 5080
rect 13924 4984 15148 5012
rect 12308 4972 12314 4984
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 16574 5012 16580 5024
rect 16264 4984 16580 5012
rect 16264 4972 16270 4984
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 16960 5012 16988 5052
rect 20809 5049 20821 5052
rect 20855 5049 20867 5083
rect 20809 5043 20867 5049
rect 17770 5012 17776 5024
rect 16724 4984 16988 5012
rect 17731 4984 17776 5012
rect 16724 4972 16730 4984
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18414 4972 18420 5024
rect 18472 5012 18478 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 18472 4984 18613 5012
rect 18472 4972 18478 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 18601 4975 18659 4981
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 20073 5015 20131 5021
rect 20073 5012 20085 5015
rect 19392 4984 20085 5012
rect 19392 4972 19398 4984
rect 20073 4981 20085 4984
rect 20119 4981 20131 5015
rect 20073 4975 20131 4981
rect 21269 5015 21327 5021
rect 21269 4981 21281 5015
rect 21315 5012 21327 5015
rect 21729 5015 21787 5021
rect 21729 5012 21741 5015
rect 21315 4984 21741 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 21729 4981 21741 4984
rect 21775 4981 21787 5015
rect 21729 4975 21787 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4777 1823 4811
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 1765 4771 1823 4777
rect 1780 4740 1808 4771
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 3142 4808 3148 4820
rect 3103 4780 3148 4808
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4120 4780 5181 4808
rect 4120 4768 4126 4780
rect 5169 4777 5181 4780
rect 5215 4808 5227 4811
rect 5626 4808 5632 4820
rect 5215 4780 5632 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4808 6791 4811
rect 6822 4808 6828 4820
rect 6779 4780 6828 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 8386 4808 8392 4820
rect 7423 4780 8392 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9582 4768 9588 4820
rect 9640 4768 9646 4820
rect 10042 4808 10048 4820
rect 10003 4780 10048 4808
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10229 4811 10287 4817
rect 10229 4777 10241 4811
rect 10275 4808 10287 4811
rect 10502 4808 10508 4820
rect 10275 4780 10508 4808
rect 10275 4777 10287 4780
rect 10229 4771 10287 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10796 4780 11100 4808
rect 3160 4740 3188 4768
rect 1780 4712 3188 4740
rect 3602 4700 3608 4752
rect 3660 4740 3666 4752
rect 3660 4712 5948 4740
rect 3660 4700 3666 4712
rect 1486 4632 1492 4684
rect 1544 4672 1550 4684
rect 1673 4675 1731 4681
rect 1673 4672 1685 4675
rect 1544 4644 1685 4672
rect 1544 4632 1550 4644
rect 1673 4641 1685 4644
rect 1719 4672 1731 4675
rect 2133 4675 2191 4681
rect 2133 4672 2145 4675
rect 1719 4644 2145 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 2133 4641 2145 4644
rect 2179 4641 2191 4675
rect 2133 4635 2191 4641
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3510 4672 3516 4684
rect 3283 4644 3516 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3510 4632 3516 4644
rect 3568 4632 3574 4684
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5718 4672 5724 4684
rect 4939 4644 5724 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2498 4604 2504 4616
rect 2455 4576 2504 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3384 4576 3433 4604
rect 3384 4564 3390 4576
rect 3421 4573 3433 4576
rect 3467 4604 3479 4607
rect 3786 4604 3792 4616
rect 3467 4576 3792 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 5350 4604 5356 4616
rect 3988 4576 5356 4604
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 2832 4508 2877 4536
rect 2832 4496 2838 4508
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3988 4536 4016 4576
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5810 4604 5816 4616
rect 5771 4576 5816 4604
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 5920 4613 5948 4712
rect 7098 4700 7104 4752
rect 7156 4740 7162 4752
rect 7156 4712 9536 4740
rect 7156 4700 7162 4712
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 6604 4644 6960 4672
rect 6604 4632 6610 4644
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 5994 4604 6000 4616
rect 5951 4576 6000 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6454 4604 6460 4616
rect 6144 4576 6460 4604
rect 6144 4564 6150 4576
rect 6454 4564 6460 4576
rect 6512 4604 6518 4616
rect 6932 4613 6960 4644
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 7064 4644 7757 4672
rect 7064 4632 7070 4644
rect 7745 4641 7757 4644
rect 7791 4672 7803 4675
rect 8570 4672 8576 4684
rect 7791 4644 8576 4672
rect 7791 4641 7803 4644
rect 7745 4635 7803 4641
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6512 4576 6837 4604
rect 6512 4564 6518 4576
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 7834 4604 7840 4616
rect 7795 4576 7840 4604
rect 6917 4567 6975 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 7926 4564 7932 4616
rect 7984 4604 7990 4616
rect 7984 4576 8029 4604
rect 7984 4564 7990 4576
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 9508 4604 9536 4712
rect 9600 4672 9628 4768
rect 10796 4740 10824 4780
rect 10962 4749 10968 4752
rect 10956 4740 10968 4749
rect 10704 4712 10824 4740
rect 10923 4712 10968 4740
rect 10704 4681 10732 4712
rect 10956 4703 10968 4712
rect 10962 4700 10968 4703
rect 11020 4700 11026 4752
rect 11072 4740 11100 4780
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 14182 4808 14188 4820
rect 11204 4780 14188 4808
rect 11204 4768 11210 4780
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 14458 4808 14464 4820
rect 14419 4780 14464 4808
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 14921 4811 14979 4817
rect 14921 4777 14933 4811
rect 14967 4808 14979 4811
rect 15562 4808 15568 4820
rect 14967 4780 15568 4808
rect 14967 4777 14979 4780
rect 14921 4771 14979 4777
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 16390 4768 16396 4820
rect 16448 4808 16454 4820
rect 17405 4811 17463 4817
rect 17405 4808 17417 4811
rect 16448 4780 17417 4808
rect 16448 4768 16454 4780
rect 17405 4777 17417 4780
rect 17451 4808 17463 4811
rect 18046 4808 18052 4820
rect 17451 4780 18052 4808
rect 17451 4777 17463 4780
rect 17405 4771 17463 4777
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18138 4768 18144 4820
rect 18196 4808 18202 4820
rect 18506 4808 18512 4820
rect 18196 4780 18512 4808
rect 18196 4768 18202 4780
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 18690 4768 18696 4820
rect 18748 4808 18754 4820
rect 18969 4811 19027 4817
rect 18969 4808 18981 4811
rect 18748 4780 18981 4808
rect 18748 4768 18754 4780
rect 18969 4777 18981 4780
rect 19015 4777 19027 4811
rect 20530 4808 20536 4820
rect 20491 4780 20536 4808
rect 18969 4771 19027 4777
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 12612 4743 12670 4749
rect 12612 4740 12624 4743
rect 11072 4712 12112 4740
rect 10689 4675 10747 4681
rect 10689 4672 10701 4675
rect 9600 4644 10701 4672
rect 10689 4641 10701 4644
rect 10735 4641 10747 4675
rect 11974 4672 11980 4684
rect 10689 4635 10747 4641
rect 10796 4644 11980 4672
rect 10796 4604 10824 4644
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12084 4672 12112 4712
rect 12544 4712 12624 4740
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12084 4644 12357 4672
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12544 4672 12572 4712
rect 12612 4709 12624 4712
rect 12658 4740 12670 4743
rect 16574 4740 16580 4752
rect 12658 4712 16580 4740
rect 12658 4709 12670 4712
rect 12612 4703 12670 4709
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 17126 4700 17132 4752
rect 17184 4740 17190 4752
rect 19426 4749 19432 4752
rect 18325 4743 18383 4749
rect 18325 4740 18337 4743
rect 17184 4712 18337 4740
rect 17184 4700 17190 4712
rect 18325 4709 18337 4712
rect 18371 4709 18383 4743
rect 19420 4740 19432 4749
rect 19387 4712 19432 4740
rect 18325 4703 18383 4709
rect 19420 4703 19432 4712
rect 19426 4700 19432 4703
rect 19484 4700 19490 4752
rect 12345 4635 12403 4641
rect 12452 4644 12572 4672
rect 15289 4675 15347 4681
rect 12452 4604 12480 4644
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15378 4672 15384 4684
rect 15335 4644 15384 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 13998 4604 14004 4616
rect 8260 4576 9260 4604
rect 9508 4576 10824 4604
rect 12084 4576 12480 4604
rect 13959 4576 14004 4604
rect 8260 4564 8266 4576
rect 3016 4508 4016 4536
rect 3016 4496 3022 4508
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 8754 4536 8760 4548
rect 4120 4508 8760 4536
rect 4120 4496 4126 4508
rect 8754 4496 8760 4508
rect 8812 4496 8818 4548
rect 2222 4428 2228 4480
rect 2280 4468 2286 4480
rect 3970 4468 3976 4480
rect 2280 4440 3976 4468
rect 2280 4428 2286 4440
rect 3970 4428 3976 4440
rect 4028 4468 4034 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 4028 4440 4261 4468
rect 4028 4428 4034 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 5353 4471 5411 4477
rect 5353 4437 5365 4471
rect 5399 4468 5411 4471
rect 6822 4468 6828 4480
rect 5399 4440 6828 4468
rect 5399 4437 5411 4440
rect 5353 4431 5411 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4468 8539 4471
rect 8570 4468 8576 4480
rect 8527 4440 8576 4468
rect 8527 4437 8539 4440
rect 8481 4431 8539 4437
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 9088 4440 9137 4468
rect 9088 4428 9094 4440
rect 9125 4437 9137 4440
rect 9171 4437 9183 4471
rect 9232 4468 9260 4576
rect 12084 4548 12112 4576
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14642 4564 14648 4616
rect 14700 4604 14706 4616
rect 15304 4604 15332 4635
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 15556 4675 15614 4681
rect 15556 4641 15568 4675
rect 15602 4672 15614 4675
rect 15930 4672 15936 4684
rect 15602 4644 15936 4672
rect 15602 4641 15614 4644
rect 15556 4635 15614 4641
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 17310 4672 17316 4684
rect 17271 4644 17316 4672
rect 17310 4632 17316 4644
rect 17368 4672 17374 4684
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17368 4644 17969 4672
rect 17368 4632 17374 4644
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4672 18291 4675
rect 18509 4675 18567 4681
rect 18509 4672 18521 4675
rect 18279 4644 18521 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 18509 4641 18521 4644
rect 18555 4672 18567 4675
rect 18690 4672 18696 4684
rect 18555 4644 18696 4672
rect 18555 4641 18567 4644
rect 18509 4635 18567 4641
rect 18690 4632 18696 4644
rect 18748 4632 18754 4684
rect 14700 4576 15332 4604
rect 14700 4564 14706 4576
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 17460 4576 17509 4604
rect 17460 4564 17466 4576
rect 17497 4573 17509 4576
rect 17543 4604 17555 4607
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 17543 4576 18797 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 18785 4573 18797 4576
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4604 19027 4607
rect 19153 4607 19211 4613
rect 19153 4604 19165 4607
rect 19015 4576 19165 4604
rect 19015 4573 19027 4576
rect 18969 4567 19027 4573
rect 19153 4573 19165 4576
rect 19199 4573 19211 4607
rect 19153 4567 19211 4573
rect 12066 4536 12072 4548
rect 11979 4508 12072 4536
rect 12066 4496 12072 4508
rect 12124 4496 12130 4548
rect 14090 4536 14096 4548
rect 13556 4508 14096 4536
rect 13556 4468 13584 4508
rect 14090 4496 14096 4508
rect 14148 4496 14154 4548
rect 16669 4539 16727 4545
rect 16669 4505 16681 4539
rect 16715 4536 16727 4539
rect 16850 4536 16856 4548
rect 16715 4508 16856 4536
rect 16715 4505 16727 4508
rect 16669 4499 16727 4505
rect 16850 4496 16856 4508
rect 16908 4536 16914 4548
rect 18414 4536 18420 4548
rect 16908 4508 18420 4536
rect 16908 4496 16914 4508
rect 18414 4496 18420 4508
rect 18472 4496 18478 4548
rect 9232 4440 13584 4468
rect 9125 4431 9183 4437
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 13725 4471 13783 4477
rect 13725 4468 13737 4471
rect 13688 4440 13737 4468
rect 13688 4428 13694 4440
rect 13725 4437 13737 4440
rect 13771 4437 13783 4471
rect 13725 4431 13783 4437
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 15102 4468 15108 4480
rect 13872 4440 15108 4468
rect 13872 4428 13878 4440
rect 15102 4428 15108 4440
rect 15160 4428 15166 4480
rect 16942 4468 16948 4480
rect 16903 4440 16948 4468
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17218 4428 17224 4480
rect 17276 4468 17282 4480
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 17276 4440 18245 4468
rect 17276 4428 17282 4440
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 18325 4471 18383 4477
rect 18325 4437 18337 4471
rect 18371 4468 18383 4471
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 18371 4440 21097 4468
rect 18371 4437 18383 4440
rect 18325 4431 18383 4437
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3326 4264 3332 4276
rect 3287 4236 3332 4264
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 4890 4264 4896 4276
rect 3476 4236 4896 4264
rect 3476 4224 3482 4236
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 4985 4267 5043 4273
rect 4985 4233 4997 4267
rect 5031 4264 5043 4267
rect 5074 4264 5080 4276
rect 5031 4236 5080 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 5074 4224 5080 4236
rect 5132 4264 5138 4276
rect 6178 4264 6184 4276
rect 5132 4236 6184 4264
rect 5132 4224 5138 4236
rect 1486 4128 1492 4140
rect 1447 4100 1492 4128
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 5828 4137 5856 4236
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 7190 4264 7196 4276
rect 6840 4236 7196 4264
rect 6840 4140 6868 4236
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 7926 4224 7932 4276
rect 7984 4264 7990 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 7984 4236 8217 4264
rect 7984 4224 7990 4236
rect 8205 4233 8217 4236
rect 8251 4233 8263 4267
rect 8205 4227 8263 4233
rect 9030 4224 9036 4276
rect 9088 4264 9094 4276
rect 16206 4264 16212 4276
rect 9088 4236 16212 4264
rect 9088 4224 9094 4236
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 16301 4267 16359 4273
rect 16301 4233 16313 4267
rect 16347 4264 16359 4267
rect 16390 4264 16396 4276
rect 16347 4236 16396 4264
rect 16347 4233 16359 4236
rect 16301 4227 16359 4233
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 18693 4267 18751 4273
rect 18693 4264 18705 4267
rect 16632 4236 18705 4264
rect 16632 4224 16638 4236
rect 18693 4233 18705 4236
rect 18739 4264 18751 4267
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 18739 4236 18981 4264
rect 18739 4233 18751 4236
rect 18693 4227 18751 4233
rect 18969 4233 18981 4236
rect 19015 4233 19027 4267
rect 19426 4264 19432 4276
rect 19387 4236 19432 4264
rect 18969 4227 19027 4233
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 11241 4199 11299 4205
rect 11241 4165 11253 4199
rect 11287 4196 11299 4199
rect 11422 4196 11428 4208
rect 11287 4168 11428 4196
rect 11287 4165 11299 4168
rect 11241 4159 11299 4165
rect 11422 4156 11428 4168
rect 11480 4156 11486 4208
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 11790 4196 11796 4208
rect 11664 4168 11796 4196
rect 11664 4156 11670 4168
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 12584 4168 13032 4196
rect 12584 4156 12590 4168
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1912 4100 1961 4128
rect 1912 4088 1918 4100
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 5813 4131 5871 4137
rect 1949 4091 2007 4097
rect 5460 4100 5764 4128
rect 1964 4060 1992 4091
rect 3602 4060 3608 4072
rect 1964 4032 3608 4060
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 5460 4060 5488 4100
rect 5626 4060 5632 4072
rect 3988 4032 5488 4060
rect 5587 4032 5632 4060
rect 3988 4004 4016 4032
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5736 4060 5764 4100
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 6822 4128 6828 4140
rect 6735 4100 6828 4128
rect 5813 4091 5871 4097
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 9030 4128 9036 4140
rect 8711 4100 9036 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 9030 4088 9036 4100
rect 9088 4128 9094 4140
rect 9217 4131 9275 4137
rect 9217 4128 9229 4131
rect 9088 4100 9229 4128
rect 9088 4088 9094 4100
rect 9217 4097 9229 4100
rect 9263 4097 9275 4131
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9217 4091 9275 4097
rect 9324 4100 9413 4128
rect 9324 4072 9352 4100
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 7834 4060 7840 4072
rect 5736 4032 7840 4060
rect 7834 4020 7840 4032
rect 7892 4060 7898 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 7892 4032 8493 4060
rect 7892 4020 7898 4032
rect 8481 4029 8493 4032
rect 8527 4060 8539 4063
rect 8570 4060 8576 4072
rect 8527 4032 8576 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8812 4032 9137 4060
rect 8812 4020 8818 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10428 4060 10456 4091
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10928 4100 11069 4128
rect 10928 4088 10934 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12066 4128 12072 4140
rect 11931 4100 12072 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 13004 4137 13032 4168
rect 15930 4156 15936 4208
rect 15988 4196 15994 4208
rect 16025 4199 16083 4205
rect 16025 4196 16037 4199
rect 15988 4168 16037 4196
rect 15988 4156 15994 4168
rect 16025 4165 16037 4168
rect 16071 4196 16083 4199
rect 17770 4196 17776 4208
rect 16071 4168 17776 4196
rect 16071 4165 16083 4168
rect 16025 4159 16083 4165
rect 16684 4140 16712 4168
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 21729 4199 21787 4205
rect 21729 4196 21741 4199
rect 17880 4168 21741 4196
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 14642 4128 14648 4140
rect 14603 4100 14648 4128
rect 12989 4091 13047 4097
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 16850 4128 16856 4140
rect 16811 4100 16856 4128
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 17880 4128 17908 4168
rect 21729 4165 21741 4168
rect 21775 4165 21787 4199
rect 21729 4159 21787 4165
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 17644 4100 17908 4128
rect 17972 4100 20177 4128
rect 17644 4088 17650 4100
rect 12621 4063 12679 4069
rect 12621 4060 12633 4063
rect 10008 4032 12633 4060
rect 10008 4020 10014 4032
rect 12621 4029 12633 4032
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 13256 4063 13314 4069
rect 13256 4029 13268 4063
rect 13302 4060 13314 4063
rect 13630 4060 13636 4072
rect 13302 4032 13636 4060
rect 13302 4029 13314 4032
rect 13256 4023 13314 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 13731 4032 16773 4060
rect 2216 3995 2274 4001
rect 2216 3961 2228 3995
rect 2262 3992 2274 3995
rect 2498 3992 2504 4004
rect 2262 3964 2504 3992
rect 2262 3961 2274 3964
rect 2216 3955 2274 3961
rect 2498 3952 2504 3964
rect 2556 3952 2562 4004
rect 3786 3952 3792 4004
rect 3844 4001 3850 4004
rect 3844 3995 3908 4001
rect 3844 3961 3862 3995
rect 3896 3961 3908 3995
rect 3844 3955 3908 3961
rect 3844 3952 3850 3955
rect 3970 3952 3976 4004
rect 4028 3952 4034 4004
rect 5810 3992 5816 4004
rect 5276 3964 5816 3992
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 4890 3924 4896 3936
rect 2372 3896 4896 3924
rect 2372 3884 2378 3896
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5276 3933 5304 3964
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 6604 3964 7082 3992
rect 6604 3952 6610 3964
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7070 3955 7128 3961
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 8938 3992 8944 4004
rect 8352 3964 8944 3992
rect 8352 3952 8358 3964
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 10137 3995 10195 4001
rect 10137 3961 10149 3995
rect 10183 3992 10195 3995
rect 10778 3992 10784 4004
rect 10183 3964 10784 3992
rect 10183 3961 10195 3964
rect 10137 3955 10195 3961
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 13731 3992 13759 4032
rect 16761 4029 16773 4032
rect 16807 4060 16819 4063
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16807 4032 17325 4060
rect 16807 4029 16819 4032
rect 16761 4023 16819 4029
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 11020 3964 13759 3992
rect 14912 3995 14970 4001
rect 11020 3952 11026 3964
rect 14912 3961 14924 3995
rect 14958 3961 14970 3995
rect 16666 3992 16672 4004
rect 16627 3964 16672 3992
rect 14912 3955 14970 3961
rect 5261 3927 5319 3933
rect 5261 3893 5273 3927
rect 5307 3893 5319 3927
rect 5261 3887 5319 3893
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5408 3896 5733 3924
rect 5408 3884 5414 3896
rect 5721 3893 5733 3896
rect 5767 3924 5779 3927
rect 6273 3927 6331 3933
rect 6273 3924 6285 3927
rect 5767 3896 6285 3924
rect 5767 3893 5779 3896
rect 5721 3887 5779 3893
rect 6273 3893 6285 3896
rect 6319 3924 6331 3927
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 6319 3896 8677 3924
rect 6319 3893 6331 3896
rect 6273 3887 6331 3893
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 8665 3887 8723 3893
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 9122 3924 9128 3936
rect 8803 3896 9128 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9766 3924 9772 3936
rect 9727 3896 9772 3924
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 10502 3924 10508 3936
rect 10275 3896 10508 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 10928 3896 11621 3924
rect 10928 3884 10934 3896
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 11609 3887 11667 3893
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 11790 3924 11796 3936
rect 11747 3896 11796 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 14369 3927 14427 3933
rect 14369 3893 14381 3927
rect 14415 3924 14427 3927
rect 14550 3924 14556 3936
rect 14415 3896 14556 3924
rect 14415 3893 14427 3896
rect 14369 3887 14427 3893
rect 14550 3884 14556 3896
rect 14608 3924 14614 3936
rect 14927 3924 14955 3955
rect 16666 3952 16672 3964
rect 16724 3992 16730 4004
rect 17681 3995 17739 4001
rect 17681 3992 17693 3995
rect 16724 3964 17693 3992
rect 16724 3952 16730 3964
rect 17681 3961 17693 3964
rect 17727 3961 17739 3995
rect 17681 3955 17739 3961
rect 17218 3924 17224 3936
rect 14608 3896 17224 3924
rect 14608 3884 14614 3896
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 17972 3924 18000 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 19886 4060 19892 4072
rect 19300 4032 19892 4060
rect 19300 4020 19306 4032
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 18414 3952 18420 4004
rect 18472 3992 18478 4004
rect 19797 3995 19855 4001
rect 19797 3992 19809 3995
rect 18472 3964 19809 3992
rect 18472 3952 18478 3964
rect 19797 3961 19809 3964
rect 19843 3961 19855 3995
rect 19797 3955 19855 3961
rect 18230 3924 18236 3936
rect 17920 3896 18000 3924
rect 18191 3896 18236 3924
rect 17920 3884 17926 3896
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 18380 3896 20545 3924
rect 18380 3884 18386 3896
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 20898 3924 20904 3936
rect 20859 3896 20904 3924
rect 20533 3887 20591 3893
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 4062 3720 4068 3732
rect 4023 3692 4068 3720
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 4522 3720 4528 3732
rect 4479 3692 4528 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 6546 3680 6552 3732
rect 6604 3720 6610 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 6604 3692 6837 3720
rect 6604 3680 6610 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9674 3720 9680 3732
rect 9355 3692 9680 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9674 3680 9680 3692
rect 9732 3720 9738 3732
rect 9950 3720 9956 3732
rect 9732 3692 9956 3720
rect 9732 3680 9738 3692
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 10100 3692 10425 3720
rect 10100 3680 10106 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 11422 3680 11428 3732
rect 11480 3720 11486 3732
rect 12989 3723 13047 3729
rect 11480 3692 12296 3720
rect 11480 3680 11486 3692
rect 1670 3652 1676 3664
rect 1504 3624 1676 3652
rect 1504 3593 1532 3624
rect 1670 3612 1676 3624
rect 1728 3652 1734 3664
rect 3786 3652 3792 3664
rect 1728 3624 3792 3652
rect 1728 3612 1734 3624
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 5712 3655 5770 3661
rect 5712 3621 5724 3655
rect 5758 3652 5770 3655
rect 5994 3652 6000 3664
rect 5758 3624 6000 3652
rect 5758 3621 5770 3624
rect 5712 3615 5770 3621
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 7742 3612 7748 3664
rect 7800 3652 7806 3664
rect 8202 3661 8208 3664
rect 8174 3655 8208 3661
rect 8174 3652 8186 3655
rect 7800 3624 8186 3652
rect 7800 3612 7806 3624
rect 8174 3621 8186 3624
rect 8260 3652 8266 3664
rect 8260 3624 8322 3652
rect 8174 3615 8208 3621
rect 8202 3612 8208 3615
rect 8260 3612 8266 3624
rect 8570 3612 8576 3664
rect 8628 3652 8634 3664
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 8628 3624 11621 3652
rect 8628 3612 8634 3624
rect 11609 3621 11621 3624
rect 11655 3652 11667 3655
rect 11790 3652 11796 3664
rect 11655 3624 11796 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 1762 3593 1768 3596
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3553 1547 3587
rect 1756 3584 1768 3593
rect 1723 3556 1768 3584
rect 1489 3547 1547 3553
rect 1756 3547 1768 3556
rect 1762 3544 1768 3547
rect 1820 3544 1826 3596
rect 3234 3584 3240 3596
rect 3195 3556 3240 3584
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4706 3584 4712 3596
rect 4571 3556 4712 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 6822 3584 6828 3596
rect 5491 3556 6828 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 6822 3544 6828 3556
rect 6880 3584 6886 3596
rect 7929 3587 7987 3593
rect 7929 3584 7941 3587
rect 6880 3556 7941 3584
rect 6880 3544 6886 3556
rect 7929 3553 7941 3556
rect 7975 3584 7987 3587
rect 8754 3584 8760 3596
rect 7975 3556 8760 3584
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 11885 3587 11943 3593
rect 11885 3584 11897 3587
rect 10367 3556 11897 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 11885 3553 11897 3556
rect 11931 3553 11943 3587
rect 11885 3547 11943 3553
rect 11974 3544 11980 3596
rect 12032 3584 12038 3596
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 12032 3556 12173 3584
rect 12032 3544 12038 3556
rect 12161 3553 12173 3556
rect 12207 3553 12219 3587
rect 12268 3584 12296 3692
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 15286 3720 15292 3732
rect 13035 3692 15292 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 15286 3680 15292 3692
rect 15344 3680 15350 3732
rect 15841 3723 15899 3729
rect 15841 3689 15853 3723
rect 15887 3720 15899 3723
rect 17126 3720 17132 3732
rect 15887 3692 17132 3720
rect 15887 3689 15899 3692
rect 15841 3683 15899 3689
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 17405 3723 17463 3729
rect 17405 3720 17417 3723
rect 17368 3692 17417 3720
rect 17368 3680 17374 3692
rect 17405 3689 17417 3692
rect 17451 3689 17463 3723
rect 17405 3683 17463 3689
rect 17770 3680 17776 3732
rect 17828 3720 17834 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 17828 3692 18153 3720
rect 17828 3680 17834 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 18598 3680 18604 3732
rect 18656 3720 18662 3732
rect 18877 3723 18935 3729
rect 18877 3720 18889 3723
rect 18656 3692 18889 3720
rect 18656 3680 18662 3692
rect 18877 3689 18889 3692
rect 18923 3689 18935 3723
rect 18877 3683 18935 3689
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 19426 3720 19432 3732
rect 19116 3692 19432 3720
rect 19116 3680 19122 3692
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 12437 3655 12495 3661
rect 12437 3621 12449 3655
rect 12483 3652 12495 3655
rect 12618 3652 12624 3664
rect 12483 3624 12624 3652
rect 12483 3621 12495 3624
rect 12437 3615 12495 3621
rect 12618 3612 12624 3624
rect 12676 3652 12682 3664
rect 13170 3652 13176 3664
rect 12676 3624 13176 3652
rect 12676 3612 12682 3624
rect 13170 3612 13176 3624
rect 13228 3612 13234 3664
rect 13357 3655 13415 3661
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 13998 3652 14004 3664
rect 13403 3624 14004 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 13998 3612 14004 3624
rect 14056 3612 14062 3664
rect 17865 3655 17923 3661
rect 17865 3652 17877 3655
rect 14108 3624 17877 3652
rect 13449 3587 13507 3593
rect 13449 3584 13461 3587
rect 12268 3556 13461 3584
rect 12161 3547 12219 3553
rect 13449 3553 13461 3556
rect 13495 3584 13507 3587
rect 13814 3584 13820 3596
rect 13495 3556 13820 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 4062 3516 4068 3528
rect 3559 3488 4068 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 2869 3451 2927 3457
rect 2869 3417 2881 3451
rect 2915 3448 2927 3451
rect 4632 3448 4660 3479
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 10505 3519 10563 3525
rect 10505 3516 10517 3519
rect 9364 3488 10517 3516
rect 9364 3476 9370 3488
rect 10505 3485 10517 3488
rect 10551 3516 10563 3519
rect 10962 3516 10968 3528
rect 10551 3488 10968 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10962 3476 10968 3488
rect 11020 3516 11026 3528
rect 12066 3516 12072 3528
rect 11020 3488 12072 3516
rect 11020 3476 11026 3488
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 13630 3516 13636 3528
rect 13543 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3516 13694 3528
rect 14108 3516 14136 3624
rect 17865 3621 17877 3624
rect 17911 3652 17923 3655
rect 18230 3652 18236 3664
rect 17911 3624 18236 3652
rect 17911 3621 17923 3624
rect 17865 3615 17923 3621
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 18509 3655 18567 3661
rect 18509 3621 18521 3655
rect 18555 3652 18567 3655
rect 18690 3652 18696 3664
rect 18555 3624 18696 3652
rect 18555 3621 18567 3624
rect 18509 3615 18567 3621
rect 18690 3612 18696 3624
rect 18748 3612 18754 3664
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 14332 3556 14381 3584
rect 14332 3544 14338 3556
rect 14369 3553 14381 3556
rect 14415 3584 14427 3587
rect 15013 3587 15071 3593
rect 15013 3584 15025 3587
rect 14415 3556 15025 3584
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 15013 3553 15025 3556
rect 15059 3553 15071 3587
rect 15286 3584 15292 3596
rect 15199 3556 15292 3584
rect 15013 3547 15071 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3584 15623 3587
rect 15841 3587 15899 3593
rect 15841 3584 15853 3587
rect 15611 3556 15853 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 15841 3553 15853 3556
rect 15887 3553 15899 3587
rect 16390 3584 16396 3596
rect 15841 3547 15899 3553
rect 15948 3556 16396 3584
rect 13688 3488 14136 3516
rect 14461 3519 14519 3525
rect 13688 3476 13694 3488
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14642 3516 14648 3528
rect 14603 3488 14648 3516
rect 14461 3479 14519 3485
rect 5350 3448 5356 3460
rect 2915 3420 4660 3448
rect 5184 3420 5356 3448
rect 2915 3417 2927 3420
rect 2869 3411 2927 3417
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2884 3380 2912 3411
rect 2556 3352 2912 3380
rect 2556 3340 2562 3352
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 5184 3380 5212 3420
rect 5350 3408 5356 3420
rect 5408 3408 5414 3460
rect 7742 3448 7748 3460
rect 7300 3420 7748 3448
rect 3292 3352 5212 3380
rect 3292 3340 3298 3352
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 5316 3352 5361 3380
rect 5316 3340 5322 3352
rect 6178 3340 6184 3392
rect 6236 3380 6242 3392
rect 7300 3380 7328 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 14366 3448 14372 3460
rect 13924 3420 14372 3448
rect 7466 3380 7472 3392
rect 6236 3352 7328 3380
rect 7427 3352 7472 3380
rect 6236 3340 6242 3352
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7837 3383 7895 3389
rect 7837 3349 7849 3383
rect 7883 3380 7895 3383
rect 8294 3380 8300 3392
rect 7883 3352 8300 3380
rect 7883 3349 7895 3352
rect 7837 3343 7895 3349
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 9950 3380 9956 3392
rect 9911 3352 9956 3380
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10870 3340 10876 3392
rect 10928 3380 10934 3392
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10928 3352 10977 3380
rect 10928 3340 10934 3352
rect 10965 3349 10977 3352
rect 11011 3380 11023 3383
rect 11698 3380 11704 3392
rect 11011 3352 11704 3380
rect 11011 3349 11023 3352
rect 10965 3343 11023 3349
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 11885 3383 11943 3389
rect 11885 3349 11897 3383
rect 11931 3380 11943 3383
rect 12158 3380 12164 3392
rect 11931 3352 12164 3380
rect 11931 3349 11943 3352
rect 11885 3343 11943 3349
rect 12158 3340 12164 3352
rect 12216 3380 12222 3392
rect 13924 3380 13952 3420
rect 14366 3408 14372 3420
rect 14424 3448 14430 3460
rect 14476 3448 14504 3479
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 15304 3516 15332 3544
rect 15948 3516 15976 3556
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 16669 3587 16727 3593
rect 16669 3553 16681 3587
rect 16715 3584 16727 3587
rect 17034 3584 17040 3596
rect 16715 3556 17040 3584
rect 16715 3553 16727 3556
rect 16669 3547 16727 3553
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 21085 3587 21143 3593
rect 21085 3584 21097 3587
rect 17276 3556 21097 3584
rect 17276 3544 17282 3556
rect 21085 3553 21097 3556
rect 21131 3553 21143 3587
rect 21085 3547 21143 3553
rect 15304 3488 15976 3516
rect 16025 3519 16083 3525
rect 16025 3485 16037 3519
rect 16071 3516 16083 3519
rect 16114 3516 16120 3528
rect 16071 3488 16120 3516
rect 16071 3485 16083 3488
rect 16025 3479 16083 3485
rect 16114 3476 16120 3488
rect 16172 3516 16178 3528
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 16172 3488 16497 3516
rect 16172 3476 16178 3488
rect 16485 3485 16497 3488
rect 16531 3485 16543 3519
rect 16850 3516 16856 3528
rect 16811 3488 16856 3516
rect 16485 3479 16543 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 20349 3519 20407 3525
rect 20349 3516 20361 3519
rect 16960 3488 20361 3516
rect 14424 3420 14504 3448
rect 14424 3408 14430 3420
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 16960 3448 16988 3488
rect 20349 3485 20361 3488
rect 20395 3485 20407 3519
rect 20349 3479 20407 3485
rect 15988 3420 16988 3448
rect 15988 3408 15994 3420
rect 18414 3408 18420 3460
rect 18472 3408 18478 3460
rect 19978 3448 19984 3460
rect 19939 3420 19984 3448
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 12216 3352 13952 3380
rect 14001 3383 14059 3389
rect 12216 3340 12222 3352
rect 14001 3349 14013 3383
rect 14047 3380 14059 3383
rect 14090 3380 14096 3392
rect 14047 3352 14096 3380
rect 14047 3349 14059 3352
rect 14001 3343 14059 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 17954 3340 17960 3392
rect 18012 3380 18018 3392
rect 18432 3380 18460 3408
rect 19242 3380 19248 3392
rect 18012 3352 18460 3380
rect 19203 3352 19248 3380
rect 18012 3340 18018 3352
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 19610 3380 19616 3392
rect 19571 3352 19616 3380
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 10134 3176 10140 3188
rect 4120 3148 9996 3176
rect 10095 3148 10140 3176
rect 4120 3136 4126 3148
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 1762 3108 1768 3120
rect 1719 3080 1768 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect 1762 3068 1768 3080
rect 1820 3108 1826 3120
rect 2041 3111 2099 3117
rect 2041 3108 2053 3111
rect 1820 3080 2053 3108
rect 1820 3068 1826 3080
rect 2041 3077 2053 3080
rect 2087 3108 2099 3111
rect 2409 3111 2467 3117
rect 2409 3108 2421 3111
rect 2087 3080 2421 3108
rect 2087 3077 2099 3080
rect 2041 3071 2099 3077
rect 2409 3077 2421 3080
rect 2455 3108 2467 3111
rect 2869 3111 2927 3117
rect 2455 3080 2820 3108
rect 2455 3077 2467 3080
rect 2409 3071 2467 3077
rect 2792 3040 2820 3080
rect 2869 3077 2881 3111
rect 2915 3108 2927 3111
rect 4430 3108 4436 3120
rect 2915 3080 4436 3108
rect 2915 3077 2927 3080
rect 2869 3071 2927 3077
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 7190 3108 7196 3120
rect 5592 3080 7196 3108
rect 5592 3068 5598 3080
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 7466 3068 7472 3120
rect 7524 3108 7530 3120
rect 8662 3108 8668 3120
rect 7524 3080 8668 3108
rect 7524 3068 7530 3080
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 9968 3108 9996 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 13446 3176 13452 3188
rect 10704 3148 13452 3176
rect 10704 3108 10732 3148
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 14550 3136 14556 3188
rect 14608 3176 14614 3188
rect 15102 3176 15108 3188
rect 14608 3148 15108 3176
rect 14608 3136 14614 3148
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 16301 3179 16359 3185
rect 16301 3176 16313 3179
rect 15427 3148 16313 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 16301 3145 16313 3148
rect 16347 3176 16359 3179
rect 17678 3176 17684 3188
rect 16347 3148 17684 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 9968 3080 10732 3108
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 11790 3108 11796 3120
rect 11204 3080 11796 3108
rect 11204 3068 11210 3080
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 11882 3068 11888 3120
rect 11940 3108 11946 3120
rect 19153 3111 19211 3117
rect 19153 3108 19165 3111
rect 11940 3080 19165 3108
rect 11940 3068 11946 3080
rect 19153 3077 19165 3080
rect 19199 3077 19211 3111
rect 19153 3071 19211 3077
rect 20165 3111 20223 3117
rect 20165 3077 20177 3111
rect 20211 3108 20223 3111
rect 20806 3108 20812 3120
rect 20211 3080 20812 3108
rect 20211 3077 20223 3080
rect 20165 3071 20223 3077
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 3510 3040 3516 3052
rect 2792 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 3660 3012 4537 3040
rect 3660 3000 3666 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 5776 3012 6193 3040
rect 5776 3000 5782 3012
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7742 3040 7748 3052
rect 7699 3012 7748 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 8294 3040 8300 3052
rect 8255 3012 8300 3040
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11057 3043 11115 3049
rect 11057 3040 11069 3043
rect 11020 3012 11069 3040
rect 11020 3000 11026 3012
rect 11057 3009 11069 3012
rect 11103 3009 11115 3043
rect 15930 3040 15936 3052
rect 11057 3003 11115 3009
rect 12636 3012 15936 3040
rect 1026 2932 1032 2984
rect 1084 2972 1090 2984
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 1084 2944 2697 2972
rect 1084 2932 1090 2944
rect 2685 2941 2697 2944
rect 2731 2972 2743 2975
rect 3237 2975 3295 2981
rect 3237 2972 3249 2975
rect 2731 2944 3249 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 3237 2941 3249 2944
rect 3283 2972 3295 2975
rect 3418 2972 3424 2984
rect 3283 2944 3424 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2972 3847 2975
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3835 2944 3893 2972
rect 3835 2941 3847 2944
rect 3789 2935 3847 2941
rect 3881 2941 3893 2944
rect 3927 2972 3939 2975
rect 4614 2972 4620 2984
rect 3927 2944 4620 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 4792 2975 4850 2981
rect 4792 2941 4804 2975
rect 4838 2972 4850 2975
rect 5074 2972 5080 2984
rect 4838 2944 5080 2972
rect 4838 2941 4850 2944
rect 4792 2935 4850 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 5368 2944 7389 2972
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 5368 2904 5396 2944
rect 7377 2941 7389 2944
rect 7423 2972 7435 2975
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7423 2944 8033 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 8021 2941 8033 2944
rect 8067 2972 8079 2975
rect 8570 2972 8576 2984
rect 8067 2944 8576 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 8754 2972 8760 2984
rect 8715 2944 8760 2972
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 9824 2944 11529 2972
rect 9824 2932 9830 2944
rect 11517 2941 11529 2944
rect 11563 2972 11575 2975
rect 11563 2944 12020 2972
rect 11563 2941 11575 2944
rect 11517 2935 11575 2941
rect 624 2876 5396 2904
rect 5460 2876 8156 2904
rect 624 2864 630 2876
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 3329 2839 3387 2845
rect 3329 2836 3341 2839
rect 256 2808 3341 2836
rect 256 2796 262 2808
rect 3329 2805 3341 2808
rect 3375 2836 3387 2839
rect 3789 2839 3847 2845
rect 3789 2836 3801 2839
rect 3375 2808 3801 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 3789 2805 3801 2808
rect 3835 2805 3847 2839
rect 4430 2836 4436 2848
rect 4343 2808 4436 2836
rect 3789 2799 3847 2805
rect 4430 2796 4436 2808
rect 4488 2836 4494 2848
rect 5460 2836 5488 2876
rect 4488 2808 5488 2836
rect 4488 2796 4494 2808
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5592 2808 5917 2836
rect 5592 2796 5598 2808
rect 5905 2805 5917 2808
rect 5951 2836 5963 2839
rect 5994 2836 6000 2848
rect 5951 2808 6000 2836
rect 5951 2805 5963 2808
rect 5905 2799 5963 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 7282 2836 7288 2848
rect 7055 2808 7288 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 7466 2836 7472 2848
rect 7427 2808 7472 2836
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 8128 2836 8156 2876
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 9002 2907 9060 2913
rect 9002 2904 9014 2907
rect 8444 2876 9014 2904
rect 8444 2864 8450 2876
rect 9002 2873 9014 2876
rect 9048 2904 9060 2907
rect 9306 2904 9312 2916
rect 9048 2876 9312 2904
rect 9048 2873 9060 2876
rect 9002 2867 9060 2873
rect 9306 2864 9312 2876
rect 9364 2864 9370 2916
rect 11793 2907 11851 2913
rect 11793 2873 11805 2907
rect 11839 2904 11851 2907
rect 11882 2904 11888 2916
rect 11839 2876 11888 2904
rect 11839 2873 11851 2876
rect 11793 2867 11851 2873
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 11992 2904 12020 2944
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 12636 2904 12664 3012
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3040 16083 3043
rect 16574 3040 16580 3052
rect 16071 3012 16580 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 16850 3000 16856 3052
rect 16908 3040 16914 3052
rect 16908 3012 18736 3040
rect 16908 3000 16914 3012
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2972 13231 2975
rect 13262 2972 13268 2984
rect 13219 2944 13268 2972
rect 13219 2941 13231 2944
rect 13173 2935 13231 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14550 2972 14556 2984
rect 14240 2944 14556 2972
rect 14240 2932 14246 2944
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 14826 2972 14832 2984
rect 14787 2944 14832 2972
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 15746 2972 15752 2984
rect 15707 2944 15752 2972
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 16301 2975 16359 2981
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 16393 2975 16451 2981
rect 16393 2972 16405 2975
rect 16347 2944 16405 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 16393 2941 16405 2944
rect 16439 2941 16451 2975
rect 16393 2935 16451 2941
rect 16942 2932 16948 2984
rect 17000 2972 17006 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 17000 2944 17141 2972
rect 17000 2932 17006 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 17770 2972 17776 2984
rect 17451 2944 17776 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 18055 2975 18113 2981
rect 18055 2941 18067 2975
rect 18101 2972 18113 2975
rect 18340 2972 18368 3012
rect 18598 2972 18604 2984
rect 18101 2944 18368 2972
rect 18559 2944 18604 2972
rect 18101 2941 18113 2944
rect 18055 2935 18113 2941
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 18708 2972 18736 3012
rect 20070 3000 20076 3052
rect 20128 3040 20134 3052
rect 22554 3040 22560 3052
rect 20128 3012 22560 3040
rect 20128 3000 20134 3012
rect 22554 3000 22560 3012
rect 22612 3000 22618 3052
rect 19794 2972 19800 2984
rect 18708 2944 19800 2972
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 20579 2944 20913 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 20901 2941 20913 2944
rect 20947 2941 20959 2975
rect 20901 2935 20959 2941
rect 11992 2876 12664 2904
rect 12710 2864 12716 2916
rect 12768 2904 12774 2916
rect 13354 2904 13360 2916
rect 12768 2876 13360 2904
rect 12768 2864 12774 2876
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 13449 2907 13507 2913
rect 13449 2873 13461 2907
rect 13495 2904 13507 2907
rect 13906 2904 13912 2916
rect 13495 2876 13912 2904
rect 13495 2873 13507 2876
rect 13449 2867 13507 2873
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 14090 2864 14096 2916
rect 14148 2904 14154 2916
rect 15841 2907 15899 2913
rect 15841 2904 15853 2907
rect 14148 2876 15853 2904
rect 14148 2864 14154 2876
rect 15841 2873 15853 2876
rect 15887 2904 15899 2907
rect 15930 2904 15936 2916
rect 15887 2876 15936 2904
rect 15887 2873 15899 2876
rect 15841 2867 15899 2873
rect 15930 2864 15936 2876
rect 15988 2864 15994 2916
rect 16669 2907 16727 2913
rect 16669 2873 16681 2907
rect 16715 2904 16727 2907
rect 17310 2904 17316 2916
rect 16715 2876 17316 2904
rect 16715 2873 16727 2876
rect 16669 2867 16727 2873
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 19521 2907 19579 2913
rect 19521 2904 19533 2907
rect 18196 2876 19533 2904
rect 18196 2864 18202 2876
rect 19521 2873 19533 2876
rect 19567 2873 19579 2907
rect 22094 2904 22100 2916
rect 19521 2867 19579 2873
rect 20732 2876 22100 2904
rect 9674 2836 9680 2848
rect 8128 2808 9680 2836
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 10505 2839 10563 2845
rect 10505 2805 10517 2839
rect 10551 2836 10563 2839
rect 10594 2836 10600 2848
rect 10551 2808 10600 2836
rect 10551 2805 10563 2808
rect 10505 2799 10563 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 10965 2839 11023 2845
rect 10965 2805 10977 2839
rect 11011 2836 11023 2839
rect 11054 2836 11060 2848
rect 11011 2808 11060 2836
rect 11011 2805 11023 2808
rect 10965 2799 11023 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11146 2796 11152 2848
rect 11204 2836 11210 2848
rect 12342 2836 12348 2848
rect 11204 2808 12348 2836
rect 11204 2796 11210 2808
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 17678 2796 17684 2848
rect 17736 2836 17742 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17736 2808 18245 2836
rect 17736 2796 17742 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 20732 2845 20760 2876
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 18785 2839 18843 2845
rect 18785 2836 18797 2839
rect 18656 2808 18797 2836
rect 18656 2796 18662 2808
rect 18785 2805 18797 2808
rect 18831 2805 18843 2839
rect 18785 2799 18843 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2805 20775 2839
rect 20717 2799 20775 2805
rect 20901 2839 20959 2845
rect 20901 2805 20913 2839
rect 20947 2836 20959 2839
rect 21177 2839 21235 2845
rect 21177 2836 21189 2839
rect 20947 2808 21189 2836
rect 20947 2805 20959 2808
rect 20901 2799 20959 2805
rect 21177 2805 21189 2808
rect 21223 2836 21235 2839
rect 21634 2836 21640 2848
rect 21223 2808 21640 2836
rect 21223 2805 21235 2808
rect 21177 2799 21235 2805
rect 21634 2796 21640 2808
rect 21692 2796 21698 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 2498 2632 2504 2644
rect 1719 2604 2504 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 2682 2592 2688 2644
rect 2740 2632 2746 2644
rect 2777 2635 2835 2641
rect 2777 2632 2789 2635
rect 2740 2604 2789 2632
rect 2740 2592 2746 2604
rect 2777 2601 2789 2604
rect 2823 2632 2835 2635
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 2823 2604 3341 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3329 2601 3341 2604
rect 3375 2632 3387 2635
rect 3970 2632 3976 2644
rect 3375 2604 3976 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 6086 2632 6092 2644
rect 5859 2604 6092 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 6273 2635 6331 2641
rect 6273 2601 6285 2635
rect 6319 2632 6331 2635
rect 7374 2632 7380 2644
rect 6319 2604 7380 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 8352 2604 9045 2632
rect 8352 2592 8358 2604
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 9033 2595 9091 2601
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10594 2632 10600 2644
rect 10275 2604 10600 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 11112 2604 11529 2632
rect 11112 2592 11118 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 12066 2632 12072 2644
rect 11940 2604 12072 2632
rect 11940 2592 11946 2604
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12618 2592 12624 2644
rect 12676 2632 12682 2644
rect 12676 2604 13768 2632
rect 12676 2592 12682 2604
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 2958 2564 2964 2576
rect 2087 2536 2964 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 3878 2564 3884 2576
rect 3344 2536 3884 2564
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 2832 2468 3249 2496
rect 2832 2456 2838 2468
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 3237 2459 3295 2465
rect 2869 2363 2927 2369
rect 2869 2329 2881 2363
rect 2915 2360 2927 2363
rect 3344 2360 3372 2536
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 4332 2567 4390 2573
rect 4332 2533 4344 2567
rect 4378 2564 4390 2567
rect 4430 2564 4436 2576
rect 4378 2536 4436 2564
rect 4378 2533 4390 2536
rect 4332 2527 4390 2533
rect 4430 2524 4436 2536
rect 4488 2524 4494 2576
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 5592 2536 6408 2564
rect 5592 2524 5598 2536
rect 3786 2456 3792 2508
rect 3844 2496 3850 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3844 2468 4077 2496
rect 3844 2456 3850 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 6181 2499 6239 2505
rect 6181 2465 6193 2499
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 3510 2428 3516 2440
rect 3423 2400 3516 2428
rect 3510 2388 3516 2400
rect 3568 2428 3574 2440
rect 3568 2400 3648 2428
rect 3568 2388 3574 2400
rect 2915 2332 3372 2360
rect 2915 2329 2927 2332
rect 2869 2323 2927 2329
rect 2409 2295 2467 2301
rect 2409 2261 2421 2295
rect 2455 2292 2467 2295
rect 2774 2292 2780 2304
rect 2455 2264 2780 2292
rect 2455 2261 2467 2264
rect 2409 2255 2467 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 3620 2292 3648 2400
rect 6196 2360 6224 2459
rect 6380 2437 6408 2536
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 7064 2536 7420 2564
rect 7064 2524 7070 2536
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7392 2505 7420 2536
rect 9950 2524 9956 2576
rect 10008 2564 10014 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 10008 2536 10149 2564
rect 10008 2524 10014 2536
rect 10137 2533 10149 2536
rect 10183 2564 10195 2567
rect 13446 2564 13452 2576
rect 10183 2536 12195 2564
rect 10183 2533 10195 2536
rect 10137 2527 10195 2533
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 7156 2468 7297 2496
rect 7156 2456 7162 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2496 7435 2499
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7423 2468 7941 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7300 2360 7328 2459
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 7742 2428 7748 2440
rect 7607 2400 7748 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 7944 2428 7972 2459
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8260 2468 9260 2496
rect 8260 2456 8266 2468
rect 9122 2428 9128 2440
rect 7944 2400 8340 2428
rect 9083 2400 9128 2428
rect 8312 2360 8340 2400
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9232 2437 9260 2468
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 10042 2496 10048 2508
rect 9732 2468 10048 2496
rect 9732 2456 9738 2468
rect 10042 2456 10048 2468
rect 10100 2496 10106 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10100 2468 10793 2496
rect 10100 2456 10106 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 11910 2499 11968 2505
rect 11910 2465 11922 2499
rect 11956 2496 11968 2499
rect 12066 2496 12072 2508
rect 11956 2468 12072 2496
rect 11956 2465 11968 2468
rect 11910 2459 11968 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12167 2496 12195 2536
rect 12636 2536 13452 2564
rect 12636 2505 12664 2536
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 12621 2499 12679 2505
rect 12167 2468 12480 2496
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 10134 2428 10140 2440
rect 9263 2400 10140 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 10134 2388 10140 2400
rect 10192 2428 10198 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10192 2400 10333 2428
rect 10192 2388 10198 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11112 2400 11253 2428
rect 11112 2388 11118 2400
rect 11241 2397 11253 2400
rect 11287 2428 11299 2431
rect 12158 2428 12164 2440
rect 11287 2400 12164 2428
rect 11287 2397 11299 2400
rect 11241 2391 11299 2397
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12452 2428 12480 2468
rect 12621 2465 12633 2499
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 12710 2456 12716 2508
rect 12768 2496 12774 2508
rect 13740 2505 13768 2604
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 16393 2635 16451 2641
rect 16393 2632 16405 2635
rect 13872 2604 16405 2632
rect 13872 2592 13878 2604
rect 16393 2601 16405 2604
rect 16439 2632 16451 2635
rect 20898 2632 20904 2644
rect 16439 2604 20904 2632
rect 16439 2601 16451 2604
rect 16393 2595 16451 2601
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 19242 2564 19248 2576
rect 13823 2536 19248 2564
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12768 2468 13185 2496
rect 12768 2456 12774 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2465 13783 2499
rect 13725 2459 13783 2465
rect 13823 2428 13851 2536
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 13964 2468 14289 2496
rect 13964 2456 13970 2468
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 12452 2400 13851 2428
rect 14292 2428 14320 2459
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14516 2468 14841 2496
rect 14516 2456 14522 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 15194 2496 15200 2508
rect 14829 2459 14887 2465
rect 14927 2468 15200 2496
rect 14927 2428 14955 2468
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16025 2499 16083 2505
rect 16025 2465 16037 2499
rect 16071 2496 16083 2499
rect 16393 2499 16451 2505
rect 16393 2496 16405 2499
rect 16071 2468 16405 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16393 2465 16405 2468
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2496 16635 2499
rect 16666 2496 16672 2508
rect 16623 2468 16672 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 17586 2456 17592 2508
rect 17644 2496 17650 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17644 2468 17693 2496
rect 17644 2456 17650 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 17770 2456 17776 2508
rect 17828 2496 17834 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17828 2468 18337 2496
rect 17828 2456 17834 2468
rect 18325 2465 18337 2468
rect 18371 2496 18383 2499
rect 18782 2496 18788 2508
rect 18371 2468 18788 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18782 2456 18788 2468
rect 18840 2456 18846 2508
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 19150 2496 19156 2508
rect 18923 2468 19156 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 19150 2456 19156 2468
rect 19208 2456 19214 2508
rect 19705 2499 19763 2505
rect 19705 2465 19717 2499
rect 19751 2496 19763 2499
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19751 2468 19993 2496
rect 19751 2465 19763 2468
rect 19705 2459 19763 2465
rect 19981 2465 19993 2468
rect 20027 2496 20039 2499
rect 20070 2496 20076 2508
rect 20027 2468 20076 2496
rect 20027 2465 20039 2468
rect 19981 2459 20039 2465
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 17954 2428 17960 2440
rect 14292 2400 14955 2428
rect 15212 2400 17960 2428
rect 9674 2360 9680 2372
rect 6196 2332 6960 2360
rect 7300 2332 8248 2360
rect 8312 2332 9680 2360
rect 6932 2304 6960 2332
rect 8220 2304 8248 2332
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 10502 2360 10508 2372
rect 9815 2332 10508 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 10502 2320 10508 2332
rect 10560 2360 10566 2372
rect 15212 2360 15240 2400
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 20162 2428 20168 2440
rect 20123 2400 20168 2428
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 10560 2332 15240 2360
rect 10560 2320 10566 2332
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 16209 2363 16267 2369
rect 16209 2360 16221 2363
rect 15528 2332 16221 2360
rect 15528 2320 15534 2332
rect 16209 2329 16221 2332
rect 16255 2329 16267 2363
rect 16209 2323 16267 2329
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 17313 2363 17371 2369
rect 17313 2360 17325 2363
rect 16448 2332 17325 2360
rect 16448 2320 16454 2332
rect 17313 2329 17325 2332
rect 17359 2329 17371 2363
rect 17313 2323 17371 2329
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 18509 2363 18567 2369
rect 18509 2360 18521 2363
rect 17460 2332 18521 2360
rect 17460 2320 17466 2332
rect 18509 2329 18521 2332
rect 18555 2329 18567 2363
rect 18509 2323 18567 2329
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 3620 2264 5457 2292
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 6914 2292 6920 2304
rect 6875 2264 6920 2292
rect 5445 2255 5503 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 8260 2264 8309 2292
rect 8260 2252 8266 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 8665 2295 8723 2301
rect 8665 2261 8677 2295
rect 8711 2292 8723 2295
rect 10778 2292 10784 2304
rect 8711 2264 10784 2292
rect 8711 2261 8723 2264
rect 8665 2255 8723 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 12069 2295 12127 2301
rect 12069 2261 12081 2295
rect 12115 2292 12127 2295
rect 12434 2292 12440 2304
rect 12115 2264 12440 2292
rect 12115 2261 12127 2264
rect 12069 2255 12127 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 12894 2292 12900 2304
rect 12851 2264 12900 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 13909 2295 13967 2301
rect 13909 2292 13921 2295
rect 13780 2264 13921 2292
rect 13780 2252 13786 2264
rect 13909 2261 13921 2264
rect 13955 2261 13967 2295
rect 13909 2255 13967 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 14240 2264 14473 2292
rect 14240 2252 14246 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 14642 2252 14648 2304
rect 14700 2292 14706 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14700 2264 15025 2292
rect 14700 2252 14706 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 15102 2252 15108 2304
rect 15160 2292 15166 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15160 2264 15669 2292
rect 15160 2252 15166 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 15930 2252 15936 2304
rect 15988 2292 15994 2304
rect 16761 2295 16819 2301
rect 16761 2292 16773 2295
rect 15988 2264 16773 2292
rect 15988 2252 15994 2264
rect 16761 2261 16773 2264
rect 16807 2261 16819 2295
rect 16761 2255 16819 2261
rect 16850 2252 16856 2304
rect 16908 2292 16914 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 16908 2264 17877 2292
rect 16908 2252 16914 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 19058 2292 19064 2304
rect 19019 2264 19064 2292
rect 17865 2255 17923 2261
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 11054 2088 11060 2100
rect 8260 2060 11060 2088
rect 8260 2048 8266 2060
rect 11054 2048 11060 2060
rect 11112 2048 11118 2100
rect 11790 2048 11796 2100
rect 11848 2088 11854 2100
rect 20162 2088 20168 2100
rect 11848 2060 20168 2088
rect 11848 2048 11854 2060
rect 20162 2048 20168 2060
rect 20220 2048 20226 2100
rect 1486 1980 1492 2032
rect 1544 2020 1550 2032
rect 7006 2020 7012 2032
rect 1544 1992 7012 2020
rect 1544 1980 1550 1992
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
rect 10778 1980 10784 2032
rect 10836 2020 10842 2032
rect 17862 2020 17868 2032
rect 10836 1992 17868 2020
rect 10836 1980 10842 1992
rect 17862 1980 17868 1992
rect 17920 1980 17926 2032
rect 6914 1912 6920 1964
rect 6972 1952 6978 1964
rect 16298 1952 16304 1964
rect 6972 1924 16304 1952
rect 6972 1912 6978 1924
rect 16298 1912 16304 1924
rect 16356 1912 16362 1964
rect 9122 1776 9128 1828
rect 9180 1816 9186 1828
rect 19610 1816 19616 1828
rect 9180 1788 19616 1816
rect 9180 1776 9186 1788
rect 19610 1776 19616 1788
rect 19668 1776 19674 1828
rect 18138 1368 18144 1420
rect 18196 1408 18202 1420
rect 19058 1408 19064 1420
rect 18196 1380 19064 1408
rect 18196 1368 18202 1380
rect 19058 1368 19064 1380
rect 19116 1368 19122 1420
rect 1946 1300 1952 1352
rect 2004 1340 2010 1352
rect 2682 1340 2688 1352
rect 2004 1312 2688 1340
rect 2004 1300 2010 1312
rect 2682 1300 2688 1312
rect 2740 1300 2746 1352
<< via1 >>
rect 4068 20680 4120 20732
rect 5172 20680 5224 20732
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 3148 20043 3200 20052
rect 3148 20009 3157 20043
rect 3157 20009 3191 20043
rect 3191 20009 3200 20043
rect 3148 20000 3200 20009
rect 5540 19864 5592 19916
rect 3148 19796 3200 19848
rect 2872 19728 2924 19780
rect 4988 19728 5040 19780
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 3056 19660 3108 19712
rect 5632 19660 5684 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 1860 19252 1912 19304
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 4988 19320 5040 19372
rect 3148 19295 3200 19304
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 4068 19184 4120 19236
rect 9036 19252 9088 19304
rect 5540 19227 5592 19236
rect 5540 19193 5549 19227
rect 5549 19193 5583 19227
rect 5583 19193 5592 19227
rect 5540 19184 5592 19193
rect 6276 19184 6328 19236
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2964 19116 3016 19168
rect 3148 19116 3200 19168
rect 3516 19116 3568 19168
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 5908 19159 5960 19168
rect 5908 19125 5917 19159
rect 5917 19125 5951 19159
rect 5951 19125 5960 19159
rect 5908 19116 5960 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 3240 18912 3292 18964
rect 4068 18912 4120 18964
rect 1860 18844 1912 18896
rect 3056 18844 3108 18896
rect 3332 18844 3384 18896
rect 4712 18844 4764 18896
rect 2320 18640 2372 18692
rect 3608 18708 3660 18760
rect 9404 18708 9456 18760
rect 3884 18640 3936 18692
rect 8944 18640 8996 18692
rect 3792 18572 3844 18624
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 4804 18572 4856 18624
rect 5908 18572 5960 18624
rect 7472 18572 7524 18624
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2780 18368 2832 18420
rect 5080 18368 5132 18420
rect 6552 18368 6604 18420
rect 2136 18300 2188 18352
rect 6276 18300 6328 18352
rect 2964 18232 3016 18284
rect 3056 18232 3108 18284
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 2412 18164 2464 18216
rect 7472 18164 7524 18216
rect 9220 18207 9272 18216
rect 3424 18096 3476 18148
rect 1400 18028 1452 18080
rect 2688 18028 2740 18080
rect 3332 18071 3384 18080
rect 3332 18037 3341 18071
rect 3341 18037 3375 18071
rect 3375 18037 3384 18071
rect 3332 18028 3384 18037
rect 3976 18071 4028 18080
rect 3976 18037 3985 18071
rect 3985 18037 4019 18071
rect 4019 18037 4028 18071
rect 3976 18028 4028 18037
rect 4160 18096 4212 18148
rect 5632 18096 5684 18148
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 9864 18164 9916 18216
rect 6276 18028 6328 18080
rect 8208 18028 8260 18080
rect 8300 18028 8352 18080
rect 10140 18028 10192 18080
rect 10324 18028 10376 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 2320 17824 2372 17876
rect 2504 17824 2556 17876
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 3884 17756 3936 17808
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 2872 17688 2924 17740
rect 5540 17620 5592 17672
rect 2596 17552 2648 17604
rect 3516 17552 3568 17604
rect 11796 17756 11848 17808
rect 10232 17731 10284 17740
rect 10232 17697 10241 17731
rect 10241 17697 10275 17731
rect 10275 17697 10284 17731
rect 10232 17688 10284 17697
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 11152 17620 11204 17672
rect 8208 17552 8260 17604
rect 9128 17552 9180 17604
rect 13268 17620 13320 17672
rect 12440 17552 12492 17604
rect 2228 17484 2280 17536
rect 2688 17484 2740 17536
rect 3608 17484 3660 17536
rect 4712 17484 4764 17536
rect 6092 17527 6144 17536
rect 6092 17493 6101 17527
rect 6101 17493 6135 17527
rect 6135 17493 6144 17527
rect 6092 17484 6144 17493
rect 6828 17484 6880 17536
rect 7472 17527 7524 17536
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 8760 17484 8812 17493
rect 12716 17527 12768 17536
rect 12716 17493 12725 17527
rect 12725 17493 12759 17527
rect 12759 17493 12768 17527
rect 12716 17484 12768 17493
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1860 17323 1912 17332
rect 1860 17289 1869 17323
rect 1869 17289 1903 17323
rect 1903 17289 1912 17323
rect 1860 17280 1912 17289
rect 6460 17280 6512 17332
rect 10232 17280 10284 17332
rect 11152 17280 11204 17332
rect 11612 17323 11664 17332
rect 11612 17289 11621 17323
rect 11621 17289 11655 17323
rect 11655 17289 11664 17323
rect 11612 17280 11664 17289
rect 2320 17212 2372 17264
rect 1768 17144 1820 17196
rect 4160 17144 4212 17196
rect 6828 17212 6880 17264
rect 13820 17255 13872 17264
rect 13820 17221 13829 17255
rect 13829 17221 13863 17255
rect 13863 17221 13872 17255
rect 13820 17212 13872 17221
rect 17960 17212 18012 17264
rect 1676 17119 1728 17128
rect 1676 17085 1685 17119
rect 1685 17085 1719 17119
rect 1719 17085 1728 17119
rect 1676 17076 1728 17085
rect 2044 17076 2096 17128
rect 3148 17076 3200 17128
rect 4068 17076 4120 17128
rect 6276 17076 6328 17128
rect 6644 17076 6696 17128
rect 9680 17076 9732 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 12716 17119 12768 17128
rect 12716 17085 12750 17119
rect 12750 17085 12768 17119
rect 12716 17076 12768 17085
rect 3700 17008 3752 17060
rect 4160 17008 4212 17060
rect 4712 17008 4764 17060
rect 10140 17008 10192 17060
rect 2964 16940 3016 16992
rect 3516 16940 3568 16992
rect 3792 16983 3844 16992
rect 3792 16949 3801 16983
rect 3801 16949 3835 16983
rect 3835 16949 3844 16983
rect 3792 16940 3844 16949
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 5632 16940 5684 16949
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 8576 16983 8628 16992
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 9588 16940 9640 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2964 16736 3016 16788
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 3792 16779 3844 16788
rect 3792 16745 3801 16779
rect 3801 16745 3835 16779
rect 3835 16745 3844 16779
rect 3792 16736 3844 16745
rect 4712 16736 4764 16788
rect 6828 16736 6880 16788
rect 8300 16779 8352 16788
rect 8300 16745 8309 16779
rect 8309 16745 8343 16779
rect 8343 16745 8352 16779
rect 8300 16736 8352 16745
rect 8760 16779 8812 16788
rect 8760 16745 8769 16779
rect 8769 16745 8803 16779
rect 8803 16745 8812 16779
rect 8760 16736 8812 16745
rect 9772 16736 9824 16788
rect 10140 16736 10192 16788
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 11704 16736 11756 16788
rect 3424 16668 3476 16720
rect 3056 16643 3108 16652
rect 3056 16609 3065 16643
rect 3065 16609 3099 16643
rect 3099 16609 3108 16643
rect 3056 16600 3108 16609
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 2964 16532 3016 16584
rect 4896 16600 4948 16652
rect 5632 16668 5684 16720
rect 7380 16668 7432 16720
rect 9128 16668 9180 16720
rect 9680 16668 9732 16720
rect 7472 16600 7524 16652
rect 8576 16600 8628 16652
rect 9312 16600 9364 16652
rect 9956 16643 10008 16652
rect 9956 16609 9990 16643
rect 9990 16609 10008 16643
rect 9956 16600 10008 16609
rect 11612 16643 11664 16652
rect 11612 16609 11646 16643
rect 11646 16609 11664 16643
rect 11612 16600 11664 16609
rect 13360 16643 13412 16652
rect 13360 16609 13369 16643
rect 13369 16609 13403 16643
rect 13403 16609 13412 16643
rect 13360 16600 13412 16609
rect 13728 16600 13780 16652
rect 9404 16507 9456 16516
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 4804 16396 4856 16448
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 7472 16396 7524 16405
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 9956 16396 10008 16448
rect 13820 16532 13872 16584
rect 12716 16507 12768 16516
rect 12716 16473 12725 16507
rect 12725 16473 12759 16507
rect 12759 16473 12768 16507
rect 12716 16464 12768 16473
rect 12440 16396 12492 16448
rect 13084 16396 13136 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1768 16235 1820 16244
rect 1768 16201 1777 16235
rect 1777 16201 1811 16235
rect 1811 16201 1820 16235
rect 1768 16192 1820 16201
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 3516 16192 3568 16244
rect 2044 16056 2096 16108
rect 4252 16192 4304 16244
rect 6092 16192 6144 16244
rect 3700 16124 3752 16176
rect 3792 16031 3844 16040
rect 2320 15920 2372 15972
rect 3792 15997 3801 16031
rect 3801 15997 3835 16031
rect 3835 15997 3844 16031
rect 3792 15988 3844 15997
rect 4160 16056 4212 16108
rect 4896 16056 4948 16108
rect 6092 16099 6144 16108
rect 6092 16065 6101 16099
rect 6101 16065 6135 16099
rect 6135 16065 6144 16099
rect 6092 16056 6144 16065
rect 6828 16056 6880 16108
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 9128 16192 9180 16244
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 9772 16192 9824 16201
rect 10324 16192 10376 16244
rect 11612 16192 11664 16244
rect 13820 16192 13872 16244
rect 9956 16124 10008 16176
rect 9588 16056 9640 16108
rect 10508 16056 10560 16108
rect 11060 16056 11112 16108
rect 13360 16056 13412 16108
rect 6000 16031 6052 16040
rect 6000 15997 6009 16031
rect 6009 15997 6043 16031
rect 6043 15997 6052 16031
rect 6000 15988 6052 15997
rect 5724 15920 5776 15972
rect 7472 15920 7524 15972
rect 11152 15963 11204 15972
rect 11152 15929 11161 15963
rect 11161 15929 11195 15963
rect 11195 15929 11204 15963
rect 11152 15920 11204 15929
rect 4436 15852 4488 15904
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 7564 15852 7616 15904
rect 9404 15852 9456 15904
rect 10692 15852 10744 15904
rect 12348 15852 12400 15904
rect 13728 15852 13780 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 1584 15512 1636 15564
rect 3148 15648 3200 15700
rect 3700 15648 3752 15700
rect 4896 15648 4948 15700
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 6000 15691 6052 15700
rect 6000 15657 6009 15691
rect 6009 15657 6043 15691
rect 6043 15657 6052 15691
rect 6000 15648 6052 15657
rect 2320 15623 2372 15632
rect 2320 15589 2329 15623
rect 2329 15589 2363 15623
rect 2363 15589 2372 15623
rect 2320 15580 2372 15589
rect 2872 15580 2924 15632
rect 3424 15580 3476 15632
rect 4252 15580 4304 15632
rect 4436 15580 4488 15632
rect 4712 15580 4764 15632
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 11152 15691 11204 15700
rect 11152 15657 11161 15691
rect 11161 15657 11195 15691
rect 11195 15657 11204 15691
rect 11152 15648 11204 15657
rect 13728 15648 13780 15700
rect 8668 15623 8720 15632
rect 8668 15589 8677 15623
rect 8677 15589 8711 15623
rect 8711 15589 8720 15623
rect 8668 15580 8720 15589
rect 3976 15512 4028 15564
rect 6920 15555 6972 15564
rect 6920 15521 6954 15555
rect 6954 15521 6972 15555
rect 6920 15512 6972 15521
rect 8760 15555 8812 15564
rect 8760 15521 8769 15555
rect 8769 15521 8803 15555
rect 8803 15521 8812 15555
rect 8760 15512 8812 15521
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 10416 15512 10468 15564
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 8852 15487 8904 15496
rect 8852 15453 8861 15487
rect 8861 15453 8895 15487
rect 8895 15453 8904 15487
rect 8852 15444 8904 15453
rect 9956 15444 10008 15496
rect 10968 15444 11020 15496
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12716 15512 12768 15564
rect 3516 15351 3568 15360
rect 3516 15317 3525 15351
rect 3525 15317 3559 15351
rect 3559 15317 3568 15351
rect 3516 15308 3568 15317
rect 4988 15308 5040 15360
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 13084 15308 13136 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 1676 15147 1728 15156
rect 1676 15113 1685 15147
rect 1685 15113 1719 15147
rect 1719 15113 1728 15147
rect 1676 15104 1728 15113
rect 1584 14968 1636 15020
rect 4068 15104 4120 15156
rect 4712 15104 4764 15156
rect 5448 15104 5500 15156
rect 5632 15104 5684 15156
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 8668 15104 8720 15113
rect 8760 15104 8812 15156
rect 10508 15147 10560 15156
rect 4252 15079 4304 15088
rect 4252 15045 4261 15079
rect 4261 15045 4295 15079
rect 4295 15045 4304 15079
rect 4252 15036 4304 15045
rect 10508 15113 10517 15147
rect 10517 15113 10551 15147
rect 10551 15113 10560 15147
rect 10508 15104 10560 15113
rect 10600 15104 10652 15156
rect 11888 15104 11940 15156
rect 13268 15104 13320 15156
rect 3976 14968 4028 15020
rect 3516 14900 3568 14952
rect 6920 14968 6972 15020
rect 8208 14968 8260 15020
rect 5080 14832 5132 14884
rect 8300 14900 8352 14952
rect 9128 14943 9180 14952
rect 9128 14909 9137 14943
rect 9137 14909 9171 14943
rect 9171 14909 9180 14943
rect 9128 14900 9180 14909
rect 9956 14900 10008 14952
rect 10508 14968 10560 15020
rect 10968 14900 11020 14952
rect 2872 14764 2924 14816
rect 3332 14764 3384 14816
rect 4804 14764 4856 14816
rect 5356 14764 5408 14816
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 7656 14764 7708 14773
rect 8484 14764 8536 14816
rect 10600 14764 10652 14816
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 3148 14603 3200 14612
rect 3148 14569 3157 14603
rect 3157 14569 3191 14603
rect 3191 14569 3200 14603
rect 3148 14560 3200 14569
rect 4252 14560 4304 14612
rect 4988 14560 5040 14612
rect 5172 14560 5224 14612
rect 2136 14492 2188 14544
rect 3516 14492 3568 14544
rect 8208 14560 8260 14612
rect 10048 14560 10100 14612
rect 10784 14560 10836 14612
rect 10968 14560 11020 14612
rect 13268 14560 13320 14612
rect 6368 14492 6420 14544
rect 8760 14492 8812 14544
rect 10416 14492 10468 14544
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 2412 14424 2464 14476
rect 3792 14424 3844 14476
rect 3884 14356 3936 14408
rect 11060 14424 11112 14476
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 6644 14356 6696 14408
rect 10324 14399 10376 14408
rect 4712 14220 4764 14272
rect 6644 14220 6696 14272
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 11796 14356 11848 14408
rect 11336 14288 11388 14340
rect 14464 14288 14516 14340
rect 7380 14220 7432 14272
rect 8392 14263 8444 14272
rect 8392 14229 8401 14263
rect 8401 14229 8435 14263
rect 8435 14229 8444 14263
rect 8392 14220 8444 14229
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 10140 14263 10192 14272
rect 10140 14229 10149 14263
rect 10149 14229 10183 14263
rect 10183 14229 10192 14263
rect 10140 14220 10192 14229
rect 10232 14220 10284 14272
rect 13728 14220 13780 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 2964 14016 3016 14068
rect 4712 14016 4764 14068
rect 6552 14016 6604 14068
rect 7380 14016 7432 14068
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 8760 14059 8812 14068
rect 8760 14025 8769 14059
rect 8769 14025 8803 14059
rect 8803 14025 8812 14059
rect 8760 14016 8812 14025
rect 1952 13880 2004 13932
rect 2504 13880 2556 13932
rect 2872 13880 2924 13932
rect 3608 13880 3660 13932
rect 4252 13880 4304 13932
rect 4896 13880 4948 13932
rect 7288 13880 7340 13932
rect 8944 13948 8996 14000
rect 9496 13948 9548 14000
rect 8300 13880 8352 13932
rect 8576 13880 8628 13932
rect 3884 13855 3936 13864
rect 3884 13821 3893 13855
rect 3893 13821 3927 13855
rect 3927 13821 3936 13855
rect 3884 13812 3936 13821
rect 2872 13744 2924 13796
rect 6644 13812 6696 13864
rect 7104 13812 7156 13864
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 5540 13744 5592 13796
rect 8300 13744 8352 13796
rect 10232 13948 10284 14000
rect 10508 14016 10560 14068
rect 13268 14016 13320 14068
rect 14280 14016 14332 14068
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 15476 14016 15528 14068
rect 13360 13991 13412 14000
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 13360 13957 13369 13991
rect 13369 13957 13403 13991
rect 13403 13957 13412 13991
rect 13360 13948 13412 13957
rect 10140 13812 10192 13864
rect 4068 13676 4120 13728
rect 5172 13676 5224 13728
rect 6828 13676 6880 13728
rect 8484 13676 8536 13728
rect 8668 13676 8720 13728
rect 9956 13744 10008 13796
rect 10324 13744 10376 13796
rect 11980 13744 12032 13796
rect 12440 13744 12492 13796
rect 13084 13744 13136 13796
rect 16396 13744 16448 13796
rect 9772 13676 9824 13728
rect 10416 13676 10468 13728
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 13728 13676 13780 13728
rect 15200 13676 15252 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2780 13472 2832 13524
rect 3700 13472 3752 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 5540 13472 5592 13524
rect 5908 13472 5960 13524
rect 8576 13472 8628 13524
rect 10140 13472 10192 13524
rect 11060 13472 11112 13524
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 12900 13515 12952 13524
rect 12900 13481 12909 13515
rect 12909 13481 12943 13515
rect 12943 13481 12952 13515
rect 12900 13472 12952 13481
rect 14280 13472 14332 13524
rect 15292 13472 15344 13524
rect 15476 13515 15528 13524
rect 15476 13481 15485 13515
rect 15485 13481 15519 13515
rect 15519 13481 15528 13515
rect 15476 13472 15528 13481
rect 2136 13404 2188 13456
rect 1676 13379 1728 13388
rect 1676 13345 1685 13379
rect 1685 13345 1719 13379
rect 1719 13345 1728 13379
rect 1676 13336 1728 13345
rect 3148 13404 3200 13456
rect 9404 13404 9456 13456
rect 10048 13447 10100 13456
rect 10048 13413 10082 13447
rect 10082 13413 10100 13447
rect 10048 13404 10100 13413
rect 10968 13404 11020 13456
rect 11980 13404 12032 13456
rect 5908 13336 5960 13388
rect 7012 13336 7064 13388
rect 7380 13336 7432 13388
rect 4712 13268 4764 13320
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 4252 13200 4304 13252
rect 5816 13268 5868 13320
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 8484 13336 8536 13388
rect 12992 13336 13044 13388
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 8392 13200 8444 13252
rect 4160 13132 4212 13184
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 4804 13132 4856 13184
rect 8484 13132 8536 13184
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 8944 13175 8996 13184
rect 8944 13141 8953 13175
rect 8953 13141 8987 13175
rect 8987 13141 8996 13175
rect 8944 13132 8996 13141
rect 10784 13200 10836 13252
rect 12256 13200 12308 13252
rect 17316 13200 17368 13252
rect 11612 13132 11664 13184
rect 15200 13132 15252 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 4252 12928 4304 12980
rect 5172 12928 5224 12980
rect 5264 12928 5316 12980
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 2504 12724 2556 12776
rect 3608 12792 3660 12844
rect 3884 12724 3936 12776
rect 4804 12724 4856 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 6644 12792 6696 12844
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 8576 12860 8628 12912
rect 10968 12928 11020 12980
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 13452 12928 13504 12980
rect 15292 12928 15344 12980
rect 8208 12724 8260 12776
rect 8484 12724 8536 12776
rect 8944 12724 8996 12776
rect 9772 12724 9824 12776
rect 10876 12792 10928 12844
rect 2688 12656 2740 12708
rect 3056 12656 3108 12708
rect 1768 12588 1820 12640
rect 4896 12656 4948 12708
rect 3608 12588 3660 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 4436 12588 4488 12640
rect 4988 12588 5040 12640
rect 10508 12656 10560 12708
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 5908 12631 5960 12640
rect 5908 12597 5917 12631
rect 5917 12597 5951 12631
rect 5951 12597 5960 12631
rect 5908 12588 5960 12597
rect 6092 12588 6144 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7288 12588 7340 12640
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 8300 12588 8352 12640
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 11980 12588 12032 12640
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 13176 12588 13228 12640
rect 15200 12588 15252 12640
rect 15844 12588 15896 12640
rect 16396 12631 16448 12640
rect 16396 12597 16405 12631
rect 16405 12597 16439 12631
rect 16439 12597 16448 12631
rect 16396 12588 16448 12597
rect 17408 12588 17460 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 2228 12384 2280 12436
rect 4252 12384 4304 12436
rect 4436 12427 4488 12436
rect 4436 12393 4445 12427
rect 4445 12393 4479 12427
rect 4479 12393 4488 12427
rect 4436 12384 4488 12393
rect 4620 12384 4672 12436
rect 6644 12427 6696 12436
rect 4712 12316 4764 12368
rect 5448 12316 5500 12368
rect 6644 12393 6653 12427
rect 6653 12393 6687 12427
rect 6687 12393 6696 12427
rect 6644 12384 6696 12393
rect 7012 12359 7064 12368
rect 7012 12325 7021 12359
rect 7021 12325 7055 12359
rect 7055 12325 7064 12359
rect 7012 12316 7064 12325
rect 8668 12316 8720 12368
rect 9864 12384 9916 12436
rect 10048 12427 10100 12436
rect 10048 12393 10057 12427
rect 10057 12393 10091 12427
rect 10091 12393 10100 12427
rect 10048 12384 10100 12393
rect 10876 12384 10928 12436
rect 11060 12384 11112 12436
rect 12624 12384 12676 12436
rect 12716 12384 12768 12436
rect 15476 12384 15528 12436
rect 20812 12384 20864 12436
rect 9956 12316 10008 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 1952 12248 2004 12300
rect 3608 12248 3660 12300
rect 4896 12248 4948 12300
rect 8300 12248 8352 12300
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 4620 12223 4672 12232
rect 3516 12180 3568 12189
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 4712 12180 4764 12232
rect 5264 12223 5316 12232
rect 5264 12189 5273 12223
rect 5273 12189 5307 12223
rect 5307 12189 5316 12223
rect 5264 12180 5316 12189
rect 6828 12180 6880 12232
rect 8208 12180 8260 12232
rect 9864 12248 9916 12300
rect 10232 12316 10284 12368
rect 11152 12248 11204 12300
rect 15568 12248 15620 12300
rect 9128 12180 9180 12232
rect 10048 12180 10100 12232
rect 10140 12180 10192 12232
rect 10508 12180 10560 12232
rect 11704 12180 11756 12232
rect 12808 12180 12860 12232
rect 3056 12044 3108 12096
rect 3516 12044 3568 12096
rect 4712 12044 4764 12096
rect 4896 12044 4948 12096
rect 11612 12112 11664 12164
rect 12072 12112 12124 12164
rect 8208 12044 8260 12096
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 9772 12044 9824 12096
rect 10968 12044 11020 12096
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 11796 12044 11848 12096
rect 12440 12044 12492 12096
rect 12532 12044 12584 12096
rect 14280 12155 14332 12164
rect 14280 12121 14289 12155
rect 14289 12121 14323 12155
rect 14323 12121 14332 12155
rect 14280 12112 14332 12121
rect 15844 12112 15896 12164
rect 16488 12112 16540 12164
rect 19064 12155 19116 12164
rect 19064 12121 19073 12155
rect 19073 12121 19107 12155
rect 19107 12121 19116 12155
rect 19064 12112 19116 12121
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 13820 12044 13872 12096
rect 15384 12044 15436 12096
rect 16396 12044 16448 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1768 11883 1820 11892
rect 1768 11849 1777 11883
rect 1777 11849 1811 11883
rect 1811 11849 1820 11883
rect 1768 11840 1820 11849
rect 4252 11840 4304 11892
rect 5448 11840 5500 11892
rect 7104 11883 7156 11892
rect 7104 11849 7113 11883
rect 7113 11849 7147 11883
rect 7147 11849 7156 11883
rect 7104 11840 7156 11849
rect 7840 11840 7892 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 6276 11772 6328 11824
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 9128 11704 9180 11756
rect 10232 11840 10284 11892
rect 9772 11772 9824 11824
rect 13544 11840 13596 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 11244 11772 11296 11824
rect 11704 11772 11756 11824
rect 12624 11772 12676 11824
rect 2964 11636 3016 11688
rect 3240 11636 3292 11688
rect 5172 11636 5224 11688
rect 6828 11636 6880 11688
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 7932 11636 7984 11688
rect 11060 11636 11112 11688
rect 12072 11636 12124 11688
rect 13728 11636 13780 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 19616 11679 19668 11688
rect 19616 11645 19625 11679
rect 19625 11645 19659 11679
rect 19659 11645 19668 11679
rect 19616 11636 19668 11645
rect 3608 11611 3660 11620
rect 3608 11577 3642 11611
rect 3642 11577 3660 11611
rect 3608 11568 3660 11577
rect 4068 11568 4120 11620
rect 4252 11568 4304 11620
rect 5356 11611 5408 11620
rect 5356 11577 5390 11611
rect 5390 11577 5408 11611
rect 5356 11568 5408 11577
rect 7840 11611 7892 11620
rect 7840 11577 7849 11611
rect 7849 11577 7883 11611
rect 7883 11577 7892 11611
rect 7840 11568 7892 11577
rect 8392 11611 8444 11620
rect 2136 11500 2188 11552
rect 2412 11500 2464 11552
rect 2780 11500 2832 11552
rect 3424 11500 3476 11552
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 8392 11577 8401 11611
rect 8401 11577 8435 11611
rect 8435 11577 8444 11611
rect 8392 11568 8444 11577
rect 12348 11568 12400 11620
rect 13636 11568 13688 11620
rect 15384 11568 15436 11620
rect 16396 11568 16448 11620
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 9404 11543 9456 11552
rect 8760 11500 8812 11509
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10784 11500 10836 11552
rect 10876 11500 10928 11552
rect 12072 11543 12124 11552
rect 12072 11509 12081 11543
rect 12081 11509 12115 11543
rect 12115 11509 12124 11543
rect 12072 11500 12124 11509
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 15200 11500 15252 11552
rect 16212 11500 16264 11552
rect 16488 11500 16540 11552
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 19248 11500 19300 11509
rect 20352 11500 20404 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2504 11296 2556 11348
rect 3056 11296 3108 11348
rect 3608 11296 3660 11348
rect 5080 11296 5132 11348
rect 7012 11296 7064 11348
rect 9404 11296 9456 11348
rect 12072 11296 12124 11348
rect 15568 11296 15620 11348
rect 16488 11296 16540 11348
rect 2320 11228 2372 11280
rect 4160 11228 4212 11280
rect 5356 11228 5408 11280
rect 5632 11271 5684 11280
rect 5632 11237 5641 11271
rect 5641 11237 5675 11271
rect 5675 11237 5684 11271
rect 5632 11228 5684 11237
rect 6828 11228 6880 11280
rect 8116 11228 8168 11280
rect 9128 11228 9180 11280
rect 9680 11228 9732 11280
rect 9956 11271 10008 11280
rect 9956 11237 9990 11271
rect 9990 11237 10008 11271
rect 9956 11228 10008 11237
rect 1492 11092 1544 11144
rect 3240 11160 3292 11212
rect 3792 11160 3844 11212
rect 4988 11160 5040 11212
rect 7380 11160 7432 11212
rect 8208 11160 8260 11212
rect 4160 11092 4212 11144
rect 6184 11135 6236 11144
rect 5448 11024 5500 11076
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 9128 11092 9180 11144
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 10784 11160 10836 11212
rect 12348 11160 12400 11212
rect 13728 11160 13780 11212
rect 15384 11160 15436 11212
rect 17592 11160 17644 11212
rect 18512 11203 18564 11212
rect 18512 11169 18521 11203
rect 18521 11169 18555 11203
rect 18555 11169 18564 11203
rect 18512 11160 18564 11169
rect 13912 11092 13964 11144
rect 15292 11092 15344 11144
rect 16396 11092 16448 11144
rect 19432 11092 19484 11144
rect 11060 11067 11112 11076
rect 11060 11033 11069 11067
rect 11069 11033 11103 11067
rect 11103 11033 11112 11067
rect 11060 11024 11112 11033
rect 12440 11024 12492 11076
rect 13360 11067 13412 11076
rect 13360 11033 13369 11067
rect 13369 11033 13403 11067
rect 13403 11033 13412 11067
rect 13360 11024 13412 11033
rect 14372 11067 14424 11076
rect 14372 11033 14381 11067
rect 14381 11033 14415 11067
rect 14415 11033 14424 11067
rect 14372 11024 14424 11033
rect 16028 11024 16080 11076
rect 16580 11024 16632 11076
rect 18604 11024 18656 11076
rect 19064 11024 19116 11076
rect 1768 10956 1820 11008
rect 1952 10956 2004 11008
rect 3056 10956 3108 11008
rect 3700 10956 3752 11008
rect 9588 10956 9640 11008
rect 9680 10956 9732 11008
rect 10784 10956 10836 11008
rect 13544 10956 13596 11008
rect 14004 10999 14056 11008
rect 14004 10965 14013 10999
rect 14013 10965 14047 10999
rect 14047 10965 14056 10999
rect 14004 10956 14056 10965
rect 15660 10956 15712 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2412 10752 2464 10804
rect 3240 10752 3292 10804
rect 2964 10684 3016 10736
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 2596 10616 2648 10668
rect 2872 10548 2924 10600
rect 3976 10548 4028 10600
rect 6184 10752 6236 10804
rect 7748 10752 7800 10804
rect 10232 10795 10284 10804
rect 8300 10684 8352 10736
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 9128 10548 9180 10600
rect 10232 10761 10241 10795
rect 10241 10761 10275 10795
rect 10275 10761 10284 10795
rect 10232 10752 10284 10761
rect 13360 10752 13412 10804
rect 16212 10752 16264 10804
rect 9956 10727 10008 10736
rect 9956 10693 9965 10727
rect 9965 10693 9999 10727
rect 9999 10693 10008 10727
rect 9956 10684 10008 10693
rect 13084 10684 13136 10736
rect 14464 10684 14516 10736
rect 17408 10752 17460 10804
rect 17960 10684 18012 10736
rect 18512 10684 18564 10736
rect 19432 10727 19484 10736
rect 19432 10693 19441 10727
rect 19441 10693 19475 10727
rect 19475 10693 19484 10727
rect 19432 10684 19484 10693
rect 14188 10616 14240 10668
rect 17592 10659 17644 10668
rect 17592 10625 17601 10659
rect 17601 10625 17635 10659
rect 17635 10625 17644 10659
rect 17592 10616 17644 10625
rect 10508 10548 10560 10600
rect 10600 10548 10652 10600
rect 11612 10548 11664 10600
rect 3792 10480 3844 10532
rect 4988 10523 5040 10532
rect 4988 10489 5022 10523
rect 5022 10489 5040 10523
rect 4988 10480 5040 10489
rect 5356 10480 5408 10532
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 3516 10412 3568 10421
rect 6000 10412 6052 10464
rect 7472 10480 7524 10532
rect 10048 10480 10100 10532
rect 7748 10412 7800 10464
rect 8208 10412 8260 10464
rect 9128 10412 9180 10464
rect 9496 10412 9548 10464
rect 9680 10412 9732 10464
rect 10784 10480 10836 10532
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 11336 10412 11388 10464
rect 14004 10548 14056 10600
rect 15016 10548 15068 10600
rect 18144 10591 18196 10600
rect 18144 10557 18153 10591
rect 18153 10557 18187 10591
rect 18187 10557 18196 10591
rect 18144 10548 18196 10557
rect 12624 10480 12676 10532
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 12992 10412 13044 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 13728 10412 13780 10464
rect 16672 10412 16724 10464
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 18972 10412 19024 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2136 10251 2188 10260
rect 2136 10217 2145 10251
rect 2145 10217 2179 10251
rect 2179 10217 2188 10251
rect 2136 10208 2188 10217
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 3516 10208 3568 10260
rect 3976 10208 4028 10260
rect 6000 10208 6052 10260
rect 7288 10208 7340 10260
rect 8576 10208 8628 10260
rect 3056 10140 3108 10192
rect 4712 10072 4764 10124
rect 5540 10072 5592 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 2688 10047 2740 10056
rect 2688 10013 2697 10047
rect 2697 10013 2731 10047
rect 2731 10013 2740 10047
rect 2688 10004 2740 10013
rect 3516 10004 3568 10056
rect 3700 10004 3752 10056
rect 7196 10072 7248 10124
rect 11796 10208 11848 10260
rect 12992 10208 13044 10260
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 17960 10208 18012 10260
rect 18604 10208 18656 10260
rect 19432 10208 19484 10260
rect 20444 10208 20496 10260
rect 8852 10004 8904 10056
rect 17592 10140 17644 10192
rect 17868 10140 17920 10192
rect 10968 10072 11020 10124
rect 11888 10072 11940 10124
rect 12440 10115 12492 10124
rect 12440 10081 12474 10115
rect 12474 10081 12492 10115
rect 12440 10072 12492 10081
rect 13268 10072 13320 10124
rect 11244 10004 11296 10056
rect 1768 9868 1820 9920
rect 4988 9868 5040 9920
rect 9036 9936 9088 9988
rect 12072 9936 12124 9988
rect 6092 9868 6144 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 8668 9868 8720 9920
rect 9128 9911 9180 9920
rect 9128 9877 9137 9911
rect 9137 9877 9171 9911
rect 9171 9877 9180 9911
rect 9128 9868 9180 9877
rect 9772 9868 9824 9920
rect 9956 9911 10008 9920
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 9956 9868 10008 9877
rect 10324 9868 10376 9920
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 13084 9868 13136 9920
rect 13728 10004 13780 10056
rect 14004 10004 14056 10056
rect 13360 9868 13412 9920
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 14280 9868 14332 9920
rect 15936 9936 15988 9988
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 16580 9911 16632 9920
rect 16580 9877 16589 9911
rect 16589 9877 16623 9911
rect 16623 9877 16632 9911
rect 16580 9868 16632 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2504 9664 2556 9716
rect 2596 9664 2648 9716
rect 7472 9664 7524 9716
rect 1768 9639 1820 9648
rect 1768 9605 1777 9639
rect 1777 9605 1811 9639
rect 1811 9605 1820 9639
rect 1768 9596 1820 9605
rect 2044 9596 2096 9648
rect 3792 9596 3844 9648
rect 5540 9596 5592 9648
rect 5632 9639 5684 9648
rect 5632 9605 5641 9639
rect 5641 9605 5675 9639
rect 5675 9605 5684 9639
rect 5632 9596 5684 9605
rect 6000 9596 6052 9648
rect 7196 9639 7248 9648
rect 7196 9605 7205 9639
rect 7205 9605 7239 9639
rect 7239 9605 7248 9639
rect 7196 9596 7248 9605
rect 16580 9664 16632 9716
rect 17960 9664 18012 9716
rect 19156 9664 19208 9716
rect 20444 9707 20496 9716
rect 20444 9673 20453 9707
rect 20453 9673 20487 9707
rect 20487 9673 20496 9707
rect 20444 9664 20496 9673
rect 2964 9571 3016 9580
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 4068 9528 4120 9580
rect 4712 9528 4764 9580
rect 5356 9528 5408 9580
rect 1308 9460 1360 9512
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 7840 9528 7892 9580
rect 8576 9528 8628 9580
rect 8300 9460 8352 9512
rect 8760 9460 8812 9512
rect 1216 9324 1268 9376
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 3240 9324 3292 9376
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 5908 9392 5960 9444
rect 7104 9392 7156 9444
rect 9680 9528 9732 9580
rect 10968 9528 11020 9580
rect 12440 9528 12492 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 15752 9596 15804 9648
rect 16948 9596 17000 9648
rect 20812 9639 20864 9648
rect 20812 9605 20821 9639
rect 20821 9605 20855 9639
rect 20855 9605 20864 9639
rect 20812 9596 20864 9605
rect 11152 9460 11204 9512
rect 11520 9460 11572 9512
rect 5448 9324 5500 9376
rect 6184 9324 6236 9376
rect 7748 9324 7800 9376
rect 9220 9324 9272 9376
rect 9404 9324 9456 9376
rect 10600 9392 10652 9444
rect 13820 9460 13872 9512
rect 12808 9435 12860 9444
rect 9772 9324 9824 9376
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 15016 9528 15068 9580
rect 18604 9528 18656 9580
rect 14188 9503 14240 9512
rect 14188 9469 14222 9503
rect 14222 9469 14240 9503
rect 14188 9460 14240 9469
rect 14648 9460 14700 9512
rect 16212 9460 16264 9512
rect 11336 9324 11388 9376
rect 12716 9324 12768 9376
rect 14372 9324 14424 9376
rect 14556 9324 14608 9376
rect 15936 9324 15988 9376
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 17224 9324 17276 9376
rect 20076 9367 20128 9376
rect 20076 9333 20085 9367
rect 20085 9333 20119 9367
rect 20119 9333 20128 9367
rect 20076 9324 20128 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2964 9052 3016 9104
rect 3792 9120 3844 9172
rect 5264 9120 5316 9172
rect 5632 9120 5684 9172
rect 7380 9120 7432 9172
rect 5356 9052 5408 9104
rect 6736 9052 6788 9104
rect 8300 9120 8352 9172
rect 9312 9163 9364 9172
rect 9312 9129 9321 9163
rect 9321 9129 9355 9163
rect 9355 9129 9364 9163
rect 9312 9120 9364 9129
rect 12624 9120 12676 9172
rect 12716 9120 12768 9172
rect 1676 8984 1728 9036
rect 3700 8984 3752 9036
rect 4804 9027 4856 9036
rect 4804 8993 4813 9027
rect 4813 8993 4847 9027
rect 4847 8993 4856 9027
rect 4804 8984 4856 8993
rect 6552 9027 6604 9036
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 3240 8916 3292 8968
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 5540 8916 5592 8968
rect 9036 9052 9088 9104
rect 10232 9052 10284 9104
rect 10968 9052 11020 9104
rect 12992 9052 13044 9104
rect 13268 9052 13320 9104
rect 14188 9120 14240 9172
rect 15108 9120 15160 9172
rect 19156 9120 19208 9172
rect 8300 8984 8352 9036
rect 11704 8984 11756 9036
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 13452 8984 13504 9036
rect 13820 9027 13872 9036
rect 13820 8993 13854 9027
rect 13854 8993 13872 9027
rect 13820 8984 13872 8993
rect 17132 9052 17184 9104
rect 17868 9052 17920 9104
rect 20720 9052 20772 9104
rect 14556 8984 14608 9036
rect 16856 8984 16908 9036
rect 3332 8848 3384 8900
rect 6092 8848 6144 8900
rect 6184 8848 6236 8900
rect 3516 8780 3568 8832
rect 5080 8780 5132 8832
rect 5908 8780 5960 8832
rect 8576 8916 8628 8968
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 8760 8848 8812 8900
rect 11428 8916 11480 8968
rect 15568 8916 15620 8968
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 17776 8916 17828 8968
rect 10968 8848 11020 8900
rect 10784 8780 10836 8832
rect 10876 8780 10928 8832
rect 11520 8848 11572 8900
rect 11704 8891 11756 8900
rect 11704 8857 11713 8891
rect 11713 8857 11747 8891
rect 11747 8857 11756 8891
rect 11704 8848 11756 8857
rect 15016 8848 15068 8900
rect 18604 8848 18656 8900
rect 13544 8780 13596 8832
rect 16580 8823 16632 8832
rect 16580 8789 16589 8823
rect 16589 8789 16623 8823
rect 16623 8789 16632 8823
rect 16580 8780 16632 8789
rect 18512 8780 18564 8832
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 18788 8780 18840 8832
rect 20076 8780 20128 8832
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2412 8576 2464 8628
rect 3332 8576 3384 8628
rect 3424 8576 3476 8628
rect 5264 8619 5316 8628
rect 2596 8508 2648 8560
rect 3792 8508 3844 8560
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 5540 8576 5592 8628
rect 6000 8576 6052 8628
rect 6736 8576 6788 8628
rect 6460 8508 6512 8560
rect 6184 8483 6236 8492
rect 2964 8372 3016 8424
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 7932 8576 7984 8628
rect 11152 8576 11204 8628
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 12072 8576 12124 8628
rect 13452 8576 13504 8628
rect 15016 8576 15068 8628
rect 8300 8508 8352 8560
rect 8576 8508 8628 8560
rect 9312 8508 9364 8560
rect 6184 8440 6236 8449
rect 3700 8372 3752 8424
rect 5172 8372 5224 8424
rect 6460 8372 6512 8424
rect 7104 8415 7156 8424
rect 7104 8381 7138 8415
rect 7138 8381 7156 8415
rect 3792 8347 3844 8356
rect 3792 8313 3801 8347
rect 3801 8313 3835 8347
rect 3835 8313 3844 8347
rect 3792 8304 3844 8313
rect 4252 8304 4304 8356
rect 7104 8372 7156 8381
rect 8576 8372 8628 8424
rect 9220 8440 9272 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 9956 8372 10008 8424
rect 10600 8372 10652 8424
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 13820 8508 13872 8560
rect 14280 8508 14332 8560
rect 15200 8508 15252 8560
rect 15568 8619 15620 8628
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 15660 8576 15712 8628
rect 20720 8576 20772 8628
rect 21180 8619 21232 8628
rect 21180 8585 21189 8619
rect 21189 8585 21223 8619
rect 21223 8585 21232 8619
rect 21180 8576 21232 8585
rect 19156 8508 19208 8560
rect 12808 8440 12860 8492
rect 14096 8440 14148 8492
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 13452 8372 13504 8424
rect 14372 8372 14424 8424
rect 14832 8372 14884 8424
rect 9680 8304 9732 8356
rect 9864 8304 9916 8356
rect 11060 8347 11112 8356
rect 11060 8313 11069 8347
rect 11069 8313 11103 8347
rect 11103 8313 11112 8347
rect 11060 8304 11112 8313
rect 12532 8304 12584 8356
rect 16856 8372 16908 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17868 8440 17920 8492
rect 18880 8372 18932 8424
rect 1584 8236 1636 8288
rect 3240 8236 3292 8288
rect 4896 8236 4948 8288
rect 5632 8236 5684 8288
rect 6000 8236 6052 8288
rect 6460 8236 6512 8288
rect 7196 8236 7248 8288
rect 7380 8236 7432 8288
rect 8208 8236 8260 8288
rect 8760 8236 8812 8288
rect 9036 8236 9088 8288
rect 13268 8236 13320 8288
rect 14096 8236 14148 8288
rect 16948 8304 17000 8356
rect 18052 8304 18104 8356
rect 18696 8304 18748 8356
rect 19340 8347 19392 8356
rect 19340 8313 19349 8347
rect 19349 8313 19383 8347
rect 19383 8313 19392 8347
rect 19340 8304 19392 8313
rect 15016 8279 15068 8288
rect 15016 8245 15025 8279
rect 15025 8245 15059 8279
rect 15059 8245 15068 8279
rect 15016 8236 15068 8245
rect 15476 8236 15528 8288
rect 17316 8236 17368 8288
rect 18328 8279 18380 8288
rect 18328 8245 18337 8279
rect 18337 8245 18371 8279
rect 18371 8245 18380 8279
rect 18328 8236 18380 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 2964 8032 3016 8084
rect 3792 8032 3844 8084
rect 4252 8032 4304 8084
rect 4712 8032 4764 8084
rect 4896 8032 4948 8084
rect 3976 7964 4028 8016
rect 6184 7964 6236 8016
rect 1952 7939 2004 7948
rect 1952 7905 1986 7939
rect 1986 7905 2004 7939
rect 1952 7896 2004 7905
rect 3700 7896 3752 7948
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5172 7828 5224 7880
rect 3056 7760 3108 7812
rect 4804 7760 4856 7812
rect 3608 7692 3660 7744
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 4712 7692 4764 7744
rect 5172 7692 5224 7744
rect 6460 7692 6512 7744
rect 6920 8032 6972 8084
rect 8852 8075 8904 8084
rect 8852 8041 8861 8075
rect 8861 8041 8895 8075
rect 8895 8041 8904 8075
rect 8852 8032 8904 8041
rect 7196 7964 7248 8016
rect 14280 8032 14332 8084
rect 15108 8032 15160 8084
rect 15752 8032 15804 8084
rect 16672 8032 16724 8084
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 17500 8032 17552 8084
rect 18696 8032 18748 8084
rect 20720 8032 20772 8084
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 9036 7896 9088 7948
rect 7472 7828 7524 7880
rect 15476 7964 15528 8016
rect 9220 7896 9272 7948
rect 10508 7896 10560 7948
rect 12072 7896 12124 7948
rect 14188 7896 14240 7948
rect 16580 7964 16632 8016
rect 15844 7896 15896 7948
rect 16672 7896 16724 7948
rect 9680 7828 9732 7880
rect 12808 7828 12860 7880
rect 15752 7828 15804 7880
rect 9036 7760 9088 7812
rect 9588 7760 9640 7812
rect 9864 7760 9916 7812
rect 7196 7692 7248 7744
rect 7288 7692 7340 7744
rect 7748 7692 7800 7744
rect 8024 7692 8076 7744
rect 9128 7692 9180 7744
rect 11796 7692 11848 7744
rect 14096 7760 14148 7812
rect 15108 7760 15160 7812
rect 15292 7760 15344 7812
rect 15568 7760 15620 7812
rect 16948 7828 17000 7880
rect 17040 7760 17092 7812
rect 12716 7692 12768 7744
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 13084 7692 13136 7744
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 15936 7692 15988 7744
rect 17776 7692 17828 7744
rect 19524 7735 19576 7744
rect 19524 7701 19533 7735
rect 19533 7701 19567 7735
rect 19567 7701 19576 7735
rect 19524 7692 19576 7701
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 20168 7735 20220 7744
rect 20168 7701 20177 7735
rect 20177 7701 20211 7735
rect 20211 7701 20220 7735
rect 20168 7692 20220 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 3148 7488 3200 7540
rect 4896 7488 4948 7540
rect 4436 7420 4488 7472
rect 4620 7420 4672 7472
rect 5264 7488 5316 7540
rect 5816 7488 5868 7540
rect 6736 7488 6788 7540
rect 9036 7531 9088 7540
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 3516 7352 3568 7404
rect 5080 7352 5132 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 6000 7420 6052 7472
rect 7472 7420 7524 7472
rect 6828 7352 6880 7404
rect 9036 7497 9045 7531
rect 9045 7497 9079 7531
rect 9079 7497 9088 7531
rect 9036 7488 9088 7497
rect 9128 7488 9180 7540
rect 12716 7488 12768 7540
rect 10508 7420 10560 7472
rect 11888 7420 11940 7472
rect 12164 7420 12216 7472
rect 12348 7420 12400 7472
rect 12624 7420 12676 7472
rect 3700 7284 3752 7336
rect 9220 7352 9272 7404
rect 12072 7352 12124 7404
rect 16396 7488 16448 7540
rect 16488 7488 16540 7540
rect 18788 7488 18840 7540
rect 15476 7420 15528 7472
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 13268 7352 13320 7404
rect 12808 7327 12860 7336
rect 1768 7148 1820 7200
rect 3332 7216 3384 7268
rect 3976 7216 4028 7268
rect 5080 7216 5132 7268
rect 3148 7148 3200 7200
rect 5356 7148 5408 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7932 7259 7984 7268
rect 7932 7225 7966 7259
rect 7966 7225 7984 7259
rect 7932 7216 7984 7225
rect 8024 7216 8076 7268
rect 9312 7216 9364 7268
rect 9404 7216 9456 7268
rect 9588 7259 9640 7268
rect 9588 7225 9611 7259
rect 9611 7225 9640 7259
rect 9588 7216 9640 7225
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 13544 7284 13596 7336
rect 14188 7327 14240 7336
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 15200 7352 15252 7404
rect 16028 7352 16080 7404
rect 17316 7352 17368 7404
rect 17960 7352 18012 7404
rect 10508 7148 10560 7200
rect 11244 7148 11296 7200
rect 11704 7148 11756 7200
rect 13820 7148 13872 7200
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 14556 7216 14608 7268
rect 19156 7284 19208 7336
rect 16488 7148 16540 7200
rect 18236 7191 18288 7200
rect 18236 7157 18245 7191
rect 18245 7157 18279 7191
rect 18279 7157 18288 7191
rect 18236 7148 18288 7157
rect 19708 7191 19760 7200
rect 19708 7157 19717 7191
rect 19717 7157 19751 7191
rect 19751 7157 19760 7191
rect 19708 7148 19760 7157
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 1952 6944 2004 6996
rect 3792 6944 3844 6996
rect 4068 6944 4120 6996
rect 9956 6944 10008 6996
rect 10968 6944 11020 6996
rect 11612 6944 11664 6996
rect 11796 6944 11848 6996
rect 11888 6944 11940 6996
rect 17224 6944 17276 6996
rect 17316 6944 17368 6996
rect 17868 6944 17920 6996
rect 18236 6944 18288 6996
rect 3516 6876 3568 6928
rect 3976 6876 4028 6928
rect 11244 6876 11296 6928
rect 1952 6808 2004 6860
rect 4068 6808 4120 6860
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 4804 6808 4856 6860
rect 6828 6808 6880 6860
rect 7472 6808 7524 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9864 6808 9916 6860
rect 10140 6808 10192 6860
rect 11612 6851 11664 6860
rect 11612 6817 11646 6851
rect 11646 6817 11664 6851
rect 11612 6808 11664 6817
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5356 6740 5408 6792
rect 6920 6740 6972 6792
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 9036 6740 9088 6792
rect 9312 6740 9364 6792
rect 2412 6672 2464 6724
rect 3884 6672 3936 6724
rect 5172 6672 5224 6724
rect 5724 6672 5776 6724
rect 6644 6672 6696 6724
rect 10416 6672 10468 6724
rect 2688 6604 2740 6656
rect 2872 6604 2924 6656
rect 5816 6604 5868 6656
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 7380 6604 7432 6656
rect 8208 6604 8260 6656
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 10968 6740 11020 6792
rect 12532 6876 12584 6928
rect 12440 6808 12492 6860
rect 15200 6876 15252 6928
rect 15568 6876 15620 6928
rect 16028 6876 16080 6928
rect 13544 6808 13596 6860
rect 14004 6808 14056 6860
rect 14096 6808 14148 6860
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 12532 6672 12584 6724
rect 16856 6808 16908 6860
rect 18696 6808 18748 6860
rect 18880 6808 18932 6860
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 18420 6783 18472 6792
rect 16028 6740 16080 6749
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 19156 6740 19208 6792
rect 19340 6740 19392 6792
rect 20812 6740 20864 6792
rect 13084 6604 13136 6656
rect 14556 6604 14608 6656
rect 17500 6604 17552 6656
rect 18512 6672 18564 6724
rect 18604 6604 18656 6656
rect 19156 6647 19208 6656
rect 19156 6613 19165 6647
rect 19165 6613 19199 6647
rect 19199 6613 19208 6647
rect 19156 6604 19208 6613
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 20168 6604 20220 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2412 6400 2464 6452
rect 3516 6400 3568 6452
rect 4068 6400 4120 6452
rect 13452 6400 13504 6452
rect 5172 6332 5224 6384
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 6920 6264 6972 6316
rect 7104 6264 7156 6316
rect 9404 6332 9456 6384
rect 10048 6375 10100 6384
rect 10048 6341 10057 6375
rect 10057 6341 10091 6375
rect 10091 6341 10100 6375
rect 10048 6332 10100 6341
rect 1400 6196 1452 6248
rect 1860 6196 1912 6248
rect 3148 6128 3200 6180
rect 5264 6196 5316 6248
rect 5632 6196 5684 6248
rect 5816 6196 5868 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 9588 6264 9640 6316
rect 9956 6264 10008 6316
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 4068 6060 4120 6112
rect 7012 6128 7064 6180
rect 7380 6128 7432 6180
rect 7748 6128 7800 6180
rect 6368 6060 6420 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 6920 6060 6972 6112
rect 7472 6060 7524 6112
rect 10416 6196 10468 6248
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 8668 6128 8720 6180
rect 9220 6060 9272 6112
rect 9588 6060 9640 6112
rect 11244 6128 11296 6180
rect 12532 6196 12584 6248
rect 19156 6400 19208 6452
rect 19340 6443 19392 6452
rect 19340 6409 19349 6443
rect 19349 6409 19383 6443
rect 19383 6409 19392 6443
rect 19340 6400 19392 6409
rect 14004 6264 14056 6316
rect 15016 6264 15068 6316
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 16856 6307 16908 6316
rect 15844 6264 15896 6273
rect 13728 6196 13780 6248
rect 15384 6196 15436 6248
rect 16396 6196 16448 6248
rect 16488 6196 16540 6248
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 17316 6264 17368 6316
rect 17500 6264 17552 6316
rect 18604 6264 18656 6316
rect 17684 6196 17736 6248
rect 18880 6196 18932 6248
rect 12716 6171 12768 6180
rect 12716 6137 12750 6171
rect 12750 6137 12768 6171
rect 12716 6128 12768 6137
rect 12992 6128 13044 6180
rect 14280 6128 14332 6180
rect 15936 6128 15988 6180
rect 11888 6060 11940 6112
rect 12164 6060 12216 6112
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 15108 6060 15160 6112
rect 16856 6128 16908 6180
rect 16672 6103 16724 6112
rect 16672 6069 16681 6103
rect 16681 6069 16715 6103
rect 16715 6069 16724 6103
rect 18052 6128 18104 6180
rect 16672 6060 16724 6069
rect 17500 6060 17552 6112
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 17776 6060 17828 6112
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2504 5856 2556 5908
rect 3976 5856 4028 5908
rect 6552 5856 6604 5908
rect 7104 5856 7156 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 9772 5856 9824 5908
rect 3884 5788 3936 5840
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 3056 5720 3108 5772
rect 4252 5720 4304 5772
rect 4896 5720 4948 5772
rect 2320 5652 2372 5704
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 2412 5584 2464 5636
rect 3332 5652 3384 5704
rect 4068 5652 4120 5704
rect 4160 5652 4212 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 5172 5652 5224 5704
rect 2504 5516 2556 5568
rect 3148 5584 3200 5636
rect 3608 5516 3660 5568
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 7288 5788 7340 5840
rect 5632 5720 5684 5772
rect 6092 5720 6144 5772
rect 6920 5720 6972 5772
rect 7104 5720 7156 5772
rect 8392 5788 8444 5840
rect 8576 5788 8628 5840
rect 11152 5856 11204 5908
rect 11244 5856 11296 5908
rect 12808 5856 12860 5908
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13268 5856 13320 5908
rect 13636 5856 13688 5908
rect 14004 5856 14056 5908
rect 11796 5831 11848 5840
rect 11796 5797 11805 5831
rect 11805 5797 11839 5831
rect 11839 5797 11848 5831
rect 11796 5788 11848 5797
rect 12716 5788 12768 5840
rect 13084 5788 13136 5840
rect 7748 5720 7800 5772
rect 9772 5720 9824 5772
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 8300 5652 8352 5704
rect 9680 5652 9732 5704
rect 9956 5720 10008 5772
rect 10416 5720 10468 5772
rect 10048 5584 10100 5636
rect 10508 5652 10560 5704
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 13544 5720 13596 5772
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 15016 5788 15068 5840
rect 16580 5788 16632 5840
rect 17500 5788 17552 5840
rect 17776 5788 17828 5840
rect 18696 5831 18748 5840
rect 18696 5797 18705 5831
rect 18705 5797 18739 5831
rect 18739 5797 18748 5831
rect 18696 5788 18748 5797
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 16488 5720 16540 5772
rect 17408 5720 17460 5772
rect 17684 5720 17736 5772
rect 19524 5720 19576 5772
rect 12992 5652 13044 5704
rect 13728 5652 13780 5704
rect 14096 5652 14148 5704
rect 12900 5584 12952 5636
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 18880 5652 18932 5704
rect 8576 5559 8628 5568
rect 8576 5525 8585 5559
rect 8585 5525 8619 5559
rect 8619 5525 8628 5559
rect 9312 5559 9364 5568
rect 8576 5516 8628 5525
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 11612 5516 11664 5568
rect 13268 5516 13320 5568
rect 15384 5516 15436 5568
rect 17868 5584 17920 5636
rect 19340 5584 19392 5636
rect 18604 5516 18656 5568
rect 19524 5516 19576 5568
rect 19892 5516 19944 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 3424 5312 3476 5364
rect 4896 5312 4948 5364
rect 4160 5244 4212 5296
rect 4712 5176 4764 5228
rect 13820 5312 13872 5364
rect 14648 5312 14700 5364
rect 15016 5312 15068 5364
rect 17408 5355 17460 5364
rect 6644 5176 6696 5228
rect 6920 5176 6972 5228
rect 7748 5176 7800 5228
rect 10968 5244 11020 5296
rect 11612 5219 11664 5228
rect 2504 5040 2556 5092
rect 2596 5040 2648 5092
rect 5724 5108 5776 5160
rect 6368 5108 6420 5160
rect 8392 5108 8444 5160
rect 11612 5185 11621 5219
rect 11621 5185 11655 5219
rect 11655 5185 11664 5219
rect 11612 5176 11664 5185
rect 4896 5040 4948 5092
rect 7012 5040 7064 5092
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2412 4972 2464 5024
rect 2872 4972 2924 5024
rect 3056 4972 3108 5024
rect 3976 4972 4028 5024
rect 5356 4972 5408 5024
rect 7104 4972 7156 5024
rect 7288 4972 7340 5024
rect 9588 5108 9640 5160
rect 9772 5151 9824 5160
rect 9772 5117 9806 5151
rect 9806 5117 9824 5151
rect 9772 5108 9824 5117
rect 12256 5108 12308 5160
rect 12716 5176 12768 5228
rect 12624 5108 12676 5160
rect 14004 5151 14056 5160
rect 14004 5117 14013 5151
rect 14013 5117 14047 5151
rect 14047 5117 14056 5151
rect 14004 5108 14056 5117
rect 14464 5176 14516 5228
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 18696 5312 18748 5364
rect 19340 5355 19392 5364
rect 19340 5321 19349 5355
rect 19349 5321 19383 5355
rect 19383 5321 19392 5355
rect 19340 5312 19392 5321
rect 17132 5244 17184 5296
rect 20536 5176 20588 5228
rect 16028 5151 16080 5160
rect 16028 5117 16037 5151
rect 16037 5117 16071 5151
rect 16071 5117 16080 5151
rect 16028 5108 16080 5117
rect 8208 4972 8260 5024
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 9956 5040 10008 5092
rect 10508 5040 10560 5092
rect 10784 4972 10836 5024
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 11244 4972 11296 5024
rect 12256 4972 12308 5024
rect 14372 5040 14424 5092
rect 16856 5040 16908 5092
rect 16212 4972 16264 5024
rect 16580 4972 16632 5024
rect 16672 4972 16724 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18420 4972 18472 5024
rect 19340 4972 19392 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 4068 4768 4120 4820
rect 5632 4768 5684 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 6828 4768 6880 4820
rect 8392 4768 8444 4820
rect 9588 4768 9640 4820
rect 10048 4811 10100 4820
rect 10048 4777 10057 4811
rect 10057 4777 10091 4811
rect 10091 4777 10100 4811
rect 10048 4768 10100 4777
rect 10508 4768 10560 4820
rect 3608 4700 3660 4752
rect 1492 4632 1544 4684
rect 3516 4632 3568 4684
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 2504 4564 2556 4616
rect 3332 4564 3384 4616
rect 3792 4564 3844 4616
rect 2780 4539 2832 4548
rect 2780 4505 2789 4539
rect 2789 4505 2823 4539
rect 2823 4505 2832 4539
rect 2780 4496 2832 4505
rect 2964 4496 3016 4548
rect 5356 4564 5408 4616
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 7104 4700 7156 4752
rect 6552 4632 6604 4684
rect 6000 4564 6052 4616
rect 6092 4564 6144 4616
rect 6460 4564 6512 4616
rect 7012 4632 7064 4684
rect 8576 4632 8628 4684
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 8208 4564 8260 4616
rect 10968 4743 11020 4752
rect 10968 4709 11002 4743
rect 11002 4709 11020 4743
rect 10968 4700 11020 4709
rect 11152 4768 11204 4820
rect 14188 4768 14240 4820
rect 14464 4811 14516 4820
rect 14464 4777 14473 4811
rect 14473 4777 14507 4811
rect 14507 4777 14516 4811
rect 14464 4768 14516 4777
rect 15568 4768 15620 4820
rect 16396 4768 16448 4820
rect 18052 4768 18104 4820
rect 18144 4768 18196 4820
rect 18512 4768 18564 4820
rect 18696 4768 18748 4820
rect 20536 4811 20588 4820
rect 20536 4777 20545 4811
rect 20545 4777 20579 4811
rect 20579 4777 20588 4811
rect 20536 4768 20588 4777
rect 11980 4632 12032 4684
rect 16580 4700 16632 4752
rect 17132 4700 17184 4752
rect 19432 4743 19484 4752
rect 19432 4709 19466 4743
rect 19466 4709 19484 4743
rect 19432 4700 19484 4709
rect 14004 4607 14056 4616
rect 4068 4496 4120 4548
rect 8760 4539 8812 4548
rect 8760 4505 8769 4539
rect 8769 4505 8803 4539
rect 8803 4505 8812 4539
rect 8760 4496 8812 4505
rect 2228 4428 2280 4480
rect 3976 4428 4028 4480
rect 6828 4428 6880 4480
rect 8576 4428 8628 4480
rect 9036 4428 9088 4480
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 14648 4564 14700 4616
rect 15384 4632 15436 4684
rect 15936 4632 15988 4684
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 18696 4632 18748 4684
rect 17408 4564 17460 4616
rect 12072 4539 12124 4548
rect 12072 4505 12081 4539
rect 12081 4505 12115 4539
rect 12115 4505 12124 4539
rect 12072 4496 12124 4505
rect 14096 4496 14148 4548
rect 16856 4496 16908 4548
rect 18420 4496 18472 4548
rect 13636 4428 13688 4480
rect 13820 4428 13872 4480
rect 15108 4428 15160 4480
rect 16948 4471 17000 4480
rect 16948 4437 16957 4471
rect 16957 4437 16991 4471
rect 16991 4437 17000 4471
rect 16948 4428 17000 4437
rect 17224 4428 17276 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 3424 4224 3476 4276
rect 4896 4224 4948 4276
rect 5080 4224 5132 4276
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 1860 4088 1912 4140
rect 6184 4224 6236 4276
rect 7196 4224 7248 4276
rect 7932 4224 7984 4276
rect 9036 4224 9088 4276
rect 16212 4224 16264 4276
rect 16396 4224 16448 4276
rect 16580 4224 16632 4276
rect 19432 4267 19484 4276
rect 19432 4233 19441 4267
rect 19441 4233 19475 4267
rect 19475 4233 19484 4267
rect 19432 4224 19484 4233
rect 11428 4156 11480 4208
rect 11612 4156 11664 4208
rect 11796 4156 11848 4208
rect 12532 4156 12584 4208
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 9036 4088 9088 4140
rect 7840 4020 7892 4072
rect 8576 4020 8628 4072
rect 8760 4020 8812 4072
rect 9312 4020 9364 4072
rect 9956 4020 10008 4072
rect 10876 4088 10928 4140
rect 12072 4088 12124 4140
rect 15936 4156 15988 4208
rect 17776 4156 17828 4208
rect 14648 4131 14700 4140
rect 14648 4097 14657 4131
rect 14657 4097 14691 4131
rect 14691 4097 14700 4131
rect 14648 4088 14700 4097
rect 16672 4088 16724 4140
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 17592 4088 17644 4140
rect 13636 4020 13688 4072
rect 2504 3952 2556 4004
rect 3792 3952 3844 4004
rect 3976 3952 4028 4004
rect 2320 3884 2372 3936
rect 4896 3884 4948 3936
rect 5816 3952 5868 4004
rect 6552 3952 6604 4004
rect 8300 3952 8352 4004
rect 8944 3952 8996 4004
rect 10784 3952 10836 4004
rect 10968 3952 11020 4004
rect 16672 3995 16724 4004
rect 5356 3884 5408 3936
rect 9128 3884 9180 3936
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 10508 3884 10560 3936
rect 10876 3884 10928 3936
rect 11796 3884 11848 3936
rect 14556 3884 14608 3936
rect 16672 3961 16681 3995
rect 16681 3961 16715 3995
rect 16715 3961 16724 3995
rect 16672 3952 16724 3961
rect 17224 3884 17276 3936
rect 17868 3884 17920 3936
rect 19248 4020 19300 4072
rect 19892 4020 19944 4072
rect 18420 3952 18472 4004
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 18328 3884 18380 3936
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 4528 3680 4580 3732
rect 6552 3680 6604 3732
rect 9680 3680 9732 3732
rect 9956 3680 10008 3732
rect 10048 3680 10100 3732
rect 11428 3680 11480 3732
rect 1676 3612 1728 3664
rect 3792 3612 3844 3664
rect 6000 3612 6052 3664
rect 7748 3612 7800 3664
rect 8208 3655 8260 3664
rect 8208 3621 8220 3655
rect 8220 3621 8260 3655
rect 8208 3612 8260 3621
rect 8576 3612 8628 3664
rect 11796 3612 11848 3664
rect 1768 3587 1820 3596
rect 1768 3553 1802 3587
rect 1802 3553 1820 3587
rect 1768 3544 1820 3553
rect 3240 3587 3292 3596
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 4712 3544 4764 3596
rect 6828 3544 6880 3596
rect 8760 3544 8812 3596
rect 11980 3544 12032 3596
rect 15292 3680 15344 3732
rect 17132 3680 17184 3732
rect 17316 3680 17368 3732
rect 17776 3680 17828 3732
rect 18604 3680 18656 3732
rect 19064 3680 19116 3732
rect 19432 3680 19484 3732
rect 12624 3612 12676 3664
rect 13176 3612 13228 3664
rect 14004 3612 14056 3664
rect 13820 3544 13872 3596
rect 4068 3476 4120 3528
rect 9312 3476 9364 3528
rect 10968 3476 11020 3528
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 13636 3519 13688 3528
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 18236 3612 18288 3664
rect 18696 3612 18748 3664
rect 14280 3544 14332 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 13636 3476 13688 3485
rect 14648 3519 14700 3528
rect 2504 3340 2556 3392
rect 3240 3340 3292 3392
rect 5356 3408 5408 3460
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 6184 3340 6236 3392
rect 7748 3408 7800 3460
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 8300 3340 8352 3392
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 10876 3340 10928 3392
rect 11704 3340 11756 3392
rect 12164 3340 12216 3392
rect 14372 3408 14424 3460
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 16396 3544 16448 3596
rect 17040 3544 17092 3596
rect 17224 3544 17276 3596
rect 16120 3476 16172 3528
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 15936 3408 15988 3460
rect 18420 3408 18472 3460
rect 19984 3451 20036 3460
rect 19984 3417 19993 3451
rect 19993 3417 20027 3451
rect 20027 3417 20036 3451
rect 19984 3408 20036 3417
rect 14096 3340 14148 3392
rect 17960 3340 18012 3392
rect 19248 3383 19300 3392
rect 19248 3349 19257 3383
rect 19257 3349 19291 3383
rect 19291 3349 19300 3383
rect 19248 3340 19300 3349
rect 19616 3383 19668 3392
rect 19616 3349 19625 3383
rect 19625 3349 19659 3383
rect 19659 3349 19668 3383
rect 19616 3340 19668 3349
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 4068 3136 4120 3188
rect 10140 3179 10192 3188
rect 1768 3068 1820 3120
rect 4436 3068 4488 3120
rect 5540 3068 5592 3120
rect 7196 3068 7248 3120
rect 7472 3068 7524 3120
rect 8668 3068 8720 3120
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 13452 3136 13504 3188
rect 14004 3179 14056 3188
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 14556 3136 14608 3188
rect 15108 3136 15160 3188
rect 17684 3136 17736 3188
rect 11152 3068 11204 3120
rect 11796 3068 11848 3120
rect 11888 3068 11940 3120
rect 20812 3068 20864 3120
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 3608 3000 3660 3052
rect 5724 3000 5776 3052
rect 7748 3000 7800 3052
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 10968 3000 11020 3052
rect 1032 2932 1084 2984
rect 3424 2932 3476 2984
rect 4620 2932 4672 2984
rect 5080 2932 5132 2984
rect 572 2864 624 2916
rect 8576 2932 8628 2984
rect 8760 2975 8812 2984
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8760 2932 8812 2941
rect 9772 2932 9824 2984
rect 204 2796 256 2848
rect 4436 2839 4488 2848
rect 4436 2805 4445 2839
rect 4445 2805 4479 2839
rect 4479 2805 4488 2839
rect 4436 2796 4488 2805
rect 5540 2796 5592 2848
rect 6000 2796 6052 2848
rect 7288 2796 7340 2848
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 7472 2796 7524 2805
rect 8392 2864 8444 2916
rect 9312 2864 9364 2916
rect 11888 2864 11940 2916
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 15936 3000 15988 3052
rect 16580 3000 16632 3052
rect 16856 3000 16908 3052
rect 13268 2932 13320 2984
rect 14188 2932 14240 2984
rect 14556 2975 14608 2984
rect 14556 2941 14565 2975
rect 14565 2941 14599 2975
rect 14599 2941 14608 2975
rect 14556 2932 14608 2941
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 15752 2975 15804 2984
rect 15752 2941 15761 2975
rect 15761 2941 15795 2975
rect 15795 2941 15804 2975
rect 15752 2932 15804 2941
rect 16948 2932 17000 2984
rect 17776 2932 17828 2984
rect 18604 2975 18656 2984
rect 18604 2941 18613 2975
rect 18613 2941 18647 2975
rect 18647 2941 18656 2975
rect 18604 2932 18656 2941
rect 20076 3000 20128 3052
rect 22560 3000 22612 3052
rect 19800 2932 19852 2984
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 12716 2907 12768 2916
rect 12716 2873 12725 2907
rect 12725 2873 12759 2907
rect 12759 2873 12768 2907
rect 12716 2864 12768 2873
rect 13360 2864 13412 2916
rect 13912 2864 13964 2916
rect 14096 2864 14148 2916
rect 15936 2864 15988 2916
rect 17316 2864 17368 2916
rect 18144 2864 18196 2916
rect 9680 2796 9732 2848
rect 10600 2796 10652 2848
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11060 2796 11112 2848
rect 11152 2796 11204 2848
rect 12348 2796 12400 2848
rect 17684 2796 17736 2848
rect 18604 2796 18656 2848
rect 22100 2864 22152 2916
rect 21640 2796 21692 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2504 2592 2556 2644
rect 2688 2592 2740 2644
rect 3976 2592 4028 2644
rect 6092 2592 6144 2644
rect 7380 2592 7432 2644
rect 8300 2592 8352 2644
rect 10600 2592 10652 2644
rect 11060 2592 11112 2644
rect 11888 2592 11940 2644
rect 12072 2592 12124 2644
rect 12624 2592 12676 2644
rect 2964 2524 3016 2576
rect 2780 2456 2832 2508
rect 3884 2524 3936 2576
rect 4436 2524 4488 2576
rect 5540 2524 5592 2576
rect 3792 2456 3844 2508
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 2780 2252 2832 2304
rect 7012 2524 7064 2576
rect 7104 2456 7156 2508
rect 9956 2524 10008 2576
rect 7748 2388 7800 2440
rect 8208 2456 8260 2508
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9680 2456 9732 2508
rect 10048 2456 10100 2508
rect 12072 2456 12124 2508
rect 13452 2524 13504 2576
rect 10140 2388 10192 2440
rect 11060 2388 11112 2440
rect 12164 2388 12216 2440
rect 12716 2456 12768 2508
rect 13820 2592 13872 2644
rect 20904 2592 20956 2644
rect 19248 2524 19300 2576
rect 13912 2456 13964 2508
rect 14464 2456 14516 2508
rect 15200 2456 15252 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 16672 2456 16724 2508
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 17592 2456 17644 2508
rect 17776 2456 17828 2508
rect 18788 2456 18840 2508
rect 19156 2456 19208 2508
rect 20076 2456 20128 2508
rect 9680 2320 9732 2372
rect 10508 2320 10560 2372
rect 17960 2388 18012 2440
rect 20168 2431 20220 2440
rect 20168 2397 20177 2431
rect 20177 2397 20211 2431
rect 20211 2397 20220 2431
rect 20168 2388 20220 2397
rect 15476 2320 15528 2372
rect 16396 2320 16448 2372
rect 17408 2320 17460 2372
rect 6920 2295 6972 2304
rect 6920 2261 6929 2295
rect 6929 2261 6963 2295
rect 6963 2261 6972 2295
rect 6920 2252 6972 2261
rect 8208 2252 8260 2304
rect 10784 2252 10836 2304
rect 12440 2252 12492 2304
rect 12900 2252 12952 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 13728 2252 13780 2304
rect 14188 2252 14240 2304
rect 14648 2252 14700 2304
rect 15108 2252 15160 2304
rect 15936 2252 15988 2304
rect 16856 2252 16908 2304
rect 19064 2295 19116 2304
rect 19064 2261 19073 2295
rect 19073 2261 19107 2295
rect 19107 2261 19116 2295
rect 19064 2252 19116 2261
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 8208 2048 8260 2100
rect 11060 2048 11112 2100
rect 11796 2048 11848 2100
rect 20168 2048 20220 2100
rect 1492 1980 1544 2032
rect 7012 1980 7064 2032
rect 10784 1980 10836 2032
rect 17868 1980 17920 2032
rect 6920 1912 6972 1964
rect 16304 1912 16356 1964
rect 9128 1776 9180 1828
rect 19616 1776 19668 1828
rect 18144 1368 18196 1420
rect 19064 1368 19116 1420
rect 1952 1300 2004 1352
rect 2688 1300 2740 1352
<< metal2 >>
rect 4066 22536 4122 22545
rect 4066 22471 4122 22480
rect 3146 22128 3202 22137
rect 3146 22063 3202 22072
rect 2778 21176 2834 21185
rect 2778 21111 2834 21120
rect 2792 20058 2820 21111
rect 2870 20632 2926 20641
rect 2870 20567 2926 20576
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 1950 19816 2006 19825
rect 2884 19786 2912 20567
rect 2962 20224 3018 20233
rect 2962 20159 3018 20168
rect 1950 19751 2006 19760
rect 2872 19780 2924 19786
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 12306 1440 18022
rect 1596 15570 1624 19110
rect 1688 17134 1716 19654
rect 1964 19514 1992 19751
rect 2872 19722 2924 19728
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2778 19272 2834 19281
rect 1872 18902 1900 19246
rect 2332 19145 2360 19246
rect 2778 19207 2834 19216
rect 2318 19136 2374 19145
rect 2318 19071 2374 19080
rect 1860 18896 1912 18902
rect 1860 18838 1912 18844
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 1964 18426 1992 18799
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 2136 18352 2188 18358
rect 1858 18320 1914 18329
rect 2136 18294 2188 18300
rect 1858 18255 1914 18264
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1780 17202 1808 17682
rect 1872 17338 1900 18255
rect 1950 17912 2006 17921
rect 1950 17847 1952 17856
rect 2004 17847 2006 17856
rect 1952 17818 2004 17824
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1950 16960 2006 16969
rect 1950 16895 2006 16904
rect 1964 16794 1992 16895
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1766 16552 1822 16561
rect 1766 16487 1822 16496
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1688 16096 1716 16390
rect 1780 16250 1808 16487
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 2056 16114 2084 17070
rect 2044 16108 2096 16114
rect 1688 16068 1808 16096
rect 1674 16008 1730 16017
rect 1674 15943 1730 15952
rect 1688 15706 1716 15943
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1674 15600 1730 15609
rect 1584 15564 1636 15570
rect 1674 15535 1730 15544
rect 1584 15506 1636 15512
rect 1596 15026 1624 15506
rect 1688 15162 1716 15535
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1582 13288 1638 13297
rect 1582 13223 1638 13232
rect 1596 12442 1624 13223
rect 1688 12730 1716 13330
rect 1780 13138 1808 16068
rect 2044 16050 2096 16056
rect 1858 14648 1914 14657
rect 1858 14583 1860 14592
rect 1912 14583 1914 14592
rect 1860 14554 1912 14560
rect 2148 14550 2176 18294
rect 2332 18222 2360 18634
rect 2792 18426 2820 19207
rect 2976 19174 3004 20159
rect 3160 20058 3188 22063
rect 3238 21584 3294 21593
rect 3238 21519 3294 21528
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 3068 18902 3096 19654
rect 3160 19310 3188 19790
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3056 18896 3108 18902
rect 3056 18838 3108 18844
rect 3160 18442 3188 19110
rect 3252 18970 3280 21519
rect 4080 20738 4108 22471
rect 4068 20732 4120 20738
rect 4068 20674 4120 20680
rect 5172 20732 5224 20738
rect 5172 20674 5224 20680
rect 4988 19780 5040 19786
rect 4988 19722 5040 19728
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 5000 19378 5028 19722
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 3516 19168 3568 19174
rect 3330 19136 3386 19145
rect 3516 19110 3568 19116
rect 3330 19071 3386 19080
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3344 18902 3372 19071
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3528 18578 3556 19110
rect 4080 18970 4108 19178
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4724 18902 4752 19110
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 3608 18760 3660 18766
rect 3660 18708 3924 18714
rect 3608 18702 3924 18708
rect 3620 18698 3924 18702
rect 3620 18692 3936 18698
rect 3620 18686 3884 18692
rect 3884 18634 3936 18640
rect 3792 18624 3844 18630
rect 3528 18550 3648 18578
rect 3792 18566 3844 18572
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2976 18414 3188 18442
rect 2976 18290 3004 18414
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 2332 17882 2360 18158
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2240 14600 2268 17478
rect 2332 17270 2360 17682
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2332 15638 2360 15914
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 2240 14572 2360 14600
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 1950 14104 2006 14113
rect 1950 14039 1952 14048
rect 2004 14039 2006 14048
rect 1952 14010 2004 14016
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1780 13110 1900 13138
rect 1688 12702 1808 12730
rect 1780 12646 1808 12702
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1780 11898 1808 12582
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10674 1532 11086
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1780 9926 1808 10950
rect 1872 10826 1900 13110
rect 1964 12782 1992 13874
rect 2148 13462 2176 14486
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 2240 12442 2268 14418
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1964 11014 1992 12242
rect 2332 11762 2360 14572
rect 2424 14482 2452 18158
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2516 13938 2544 17818
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2410 12880 2466 12889
rect 2410 12815 2466 12824
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2332 11665 2360 11698
rect 2318 11656 2374 11665
rect 2318 11591 2374 11600
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1872 10798 1992 10826
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 9654 1808 9862
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 1216 9376 1268 9382
rect 1216 9318 1268 9324
rect 1032 2984 1084 2990
rect 1032 2926 1084 2932
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 800 244 2790
rect 584 800 612 2858
rect 1044 800 1072 2926
rect 1228 2009 1256 9318
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1057 1348 9454
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6254 1440 6734
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1504 4146 1532 4626
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1492 2032 1544 2038
rect 1492 1974 1544 1980
rect 1306 1048 1362 1057
rect 1306 983 1362 992
rect 1504 800 1532 1974
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1596 241 1624 8230
rect 1688 7886 1716 8978
rect 1964 7954 1992 10798
rect 2148 10266 2176 11494
rect 2332 11286 2360 11591
rect 2424 11558 2452 12815
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2516 11354 2544 12718
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2320 11280 2372 11286
rect 2372 11240 2452 11268
rect 2320 11222 2372 11228
rect 2424 10810 2452 11240
rect 2502 11248 2558 11257
rect 2502 11183 2558 11192
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2516 10266 2544 11183
rect 2608 10674 2636 17546
rect 2700 17542 2728 18022
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 12714 2728 17478
rect 2884 15638 2912 17682
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2976 16794 3004 16934
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 3068 16658 3096 18226
rect 3160 17134 3188 18414
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3238 17368 3294 17377
rect 3238 17303 3294 17312
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3146 16960 3202 16969
rect 3146 16895 3202 16904
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2976 16250 3004 16526
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3160 15706 3188 16895
rect 3252 16794 3280 17303
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 2872 15632 2924 15638
rect 2924 15592 3004 15620
rect 2872 15574 2924 15580
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 13938 2912 14758
rect 2976 14074 3004 15592
rect 3146 15056 3202 15065
rect 3146 14991 3202 15000
rect 3160 14618 3188 14991
rect 3344 14822 3372 18022
rect 3436 16726 3464 18090
rect 3620 17626 3648 18550
rect 3516 17604 3568 17610
rect 3620 17598 3740 17626
rect 3516 17546 3568 17552
rect 3528 16998 3556 17546
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3436 15638 3464 16662
rect 3528 16250 3556 16934
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 14958 3556 15302
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3528 14550 3556 14894
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3620 13938 3648 17478
rect 3712 17066 3740 17598
rect 3804 17105 3832 18566
rect 4160 18148 4212 18154
rect 4160 18090 4212 18096
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 3790 17096 3846 17105
rect 3700 17060 3752 17066
rect 3790 17031 3846 17040
rect 3700 17002 3752 17008
rect 3712 16182 3740 17002
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3804 16794 3832 16934
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 3804 16046 3832 16730
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2792 13530 2820 13631
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2596 10668 2648 10674
rect 2648 10628 2728 10656
rect 2596 10610 2648 10616
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2516 9722 2544 10202
rect 2700 10062 2728 10628
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2608 9722 2636 9998
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 3670 1716 7822
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1780 6322 1808 7142
rect 1964 7002 1992 7890
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 4146 1900 6190
rect 1964 5914 1992 6802
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3126 1808 3538
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 2056 2961 2084 9590
rect 2318 9344 2374 9353
rect 2318 9279 2374 9288
rect 2134 9072 2190 9081
rect 2134 9007 2190 9016
rect 2042 2952 2098 2961
rect 2042 2887 2098 2896
rect 2148 2825 2176 9007
rect 2332 5710 2360 9279
rect 2410 9208 2466 9217
rect 2410 9143 2466 9152
rect 2424 8634 2452 9143
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2608 8566 2636 9658
rect 2686 9616 2742 9625
rect 2686 9551 2742 9560
rect 2700 9382 2728 9551
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2792 7970 2820 11494
rect 2884 10606 2912 13738
rect 3712 13530 3740 15642
rect 3896 14498 3924 17750
rect 3988 15570 4016 18022
rect 4172 17202 4200 18090
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16658 4108 17070
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 4080 15502 4108 16594
rect 4172 16114 4200 17002
rect 4264 16250 4292 18566
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4724 17066 4752 17478
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4724 16794 4752 17002
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4816 16674 4844 18566
rect 4724 16646 4844 16674
rect 4896 16652 4948 16658
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4448 15638 4476 15846
rect 4724 15638 4752 16646
rect 4896 16594 4948 16600
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 15910 4844 16390
rect 4908 16114 4936 16594
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 15162 4108 15438
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4264 15094 4292 15574
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3804 14482 3924 14498
rect 3792 14476 3924 14482
rect 3844 14470 3924 14476
rect 3792 14418 3844 14424
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3896 13870 3924 14350
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2962 12336 3018 12345
rect 2962 12271 3018 12280
rect 2976 11801 3004 12271
rect 3068 12102 3096 12650
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2962 11792 3018 11801
rect 2962 11727 3018 11736
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2976 10742 3004 11630
rect 3068 11354 3096 12038
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 3068 10198 3096 10950
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2870 9480 2926 9489
rect 2870 9415 2926 9424
rect 2700 7942 2820 7970
rect 2502 7848 2558 7857
rect 2502 7783 2558 7792
rect 2516 7410 2544 7783
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2424 6458 2452 6666
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2424 5642 2452 6394
rect 2516 5914 2544 7346
rect 2700 6882 2728 7942
rect 2700 6854 2820 6882
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2700 5658 2728 6598
rect 2792 5778 2820 6854
rect 2884 6662 2912 9415
rect 2976 9110 3004 9522
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2976 8430 3004 9046
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2976 8090 3004 8366
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 3068 7546 3096 7754
rect 3160 7546 3188 13398
rect 3988 12866 4016 14962
rect 4264 14618 4292 15030
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4264 13938 4292 14554
rect 4724 14414 4752 15098
rect 4816 14822 4844 15846
rect 4908 15706 4936 16050
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 5000 15366 5028 19314
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5092 14890 5120 18362
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4712 14408 4764 14414
rect 4764 14368 4844 14396
rect 4712 14350 4764 14356
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4724 14074 4752 14214
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 3608 12844 3660 12850
rect 3436 12804 3608 12832
rect 3436 12238 3464 12804
rect 3608 12786 3660 12792
rect 3804 12838 4016 12866
rect 3698 12744 3754 12753
rect 3698 12679 3754 12688
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3620 12306 3648 12582
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3252 11218 3280 11630
rect 3436 11558 3464 12174
rect 3528 12102 3556 12174
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3620 11626 3648 12242
rect 3712 11801 3740 12679
rect 3698 11792 3754 11801
rect 3698 11727 3754 11736
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3620 11354 3648 11562
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3804 11218 3832 12838
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3252 10810 3280 11154
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3712 10849 3740 10950
rect 3698 10840 3754 10849
rect 3240 10804 3292 10810
rect 3698 10775 3754 10784
rect 3240 10746 3292 10752
rect 3804 10538 3832 11154
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 10266 3556 10406
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3424 9512 3476 9518
rect 3528 9489 3556 9998
rect 3424 9454 3476 9460
rect 3514 9480 3570 9489
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 8974 3280 9318
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8294 3280 8910
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 8634 3372 8842
rect 3436 8634 3464 9454
rect 3514 9415 3570 9424
rect 3528 8838 3556 9415
rect 3712 9042 3740 9998
rect 3804 9654 3832 10474
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3804 9178 3832 9590
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3712 8430 3740 8978
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3422 8256 3478 8265
rect 3422 8191 3478 8200
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3436 7313 3464 8191
rect 3712 7954 3740 8366
rect 3804 8362 3832 8502
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 8090 3832 8298
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3146 7304 3202 7313
rect 3422 7304 3478 7313
rect 3146 7239 3202 7248
rect 3332 7268 3384 7274
rect 3160 7206 3188 7239
rect 3422 7239 3478 7248
rect 3332 7210 3384 7216
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2872 5704 2924 5710
rect 2412 5636 2464 5642
rect 2700 5630 2820 5658
rect 2872 5646 2924 5652
rect 2412 5578 2464 5584
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2516 5098 2544 5510
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2240 4865 2268 4966
rect 2226 4856 2282 4865
rect 2226 4791 2228 4800
rect 2280 4791 2282 4800
rect 2228 4762 2280 4768
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2134 2816 2190 2825
rect 2134 2751 2190 2760
rect 1952 1352 2004 1358
rect 1952 1294 2004 1300
rect 1964 800 1992 1294
rect 1582 232 1638 241
rect 1582 167 1638 176
rect 1950 0 2006 800
rect 2240 649 2268 4422
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 800 2360 3878
rect 2424 2553 2452 4966
rect 2516 4622 2544 5034
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2516 4010 2544 4558
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2516 3398 2544 3946
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 2650 2544 3334
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2410 2544 2466 2553
rect 2410 2479 2466 2488
rect 2608 1601 2636 5034
rect 2792 4706 2820 5630
rect 2884 5030 2912 5646
rect 3068 5030 3096 5714
rect 3160 5642 3188 6122
rect 3344 5710 3372 7210
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3436 5370 3464 7239
rect 3528 6934 3556 7346
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3528 6458 3556 6870
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3620 5953 3648 7686
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3606 5944 3662 5953
rect 3606 5879 3662 5888
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3146 5128 3202 5137
rect 3146 5063 3202 5072
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2700 4678 2820 4706
rect 2700 3482 2728 4678
rect 2778 4584 2834 4593
rect 2778 4519 2780 4528
rect 2832 4519 2834 4528
rect 2964 4548 3016 4554
rect 2780 4490 2832 4496
rect 2964 4490 3016 4496
rect 2778 4040 2834 4049
rect 2778 3975 2834 3984
rect 2792 3482 2820 3975
rect 2700 3454 2820 3482
rect 2778 2680 2834 2689
rect 2688 2644 2740 2650
rect 2778 2615 2834 2624
rect 2688 2586 2740 2592
rect 2594 1592 2650 1601
rect 2594 1527 2650 1536
rect 2700 1358 2728 2586
rect 2792 2514 2820 2615
rect 2976 2582 3004 4490
rect 3068 3505 3096 4966
rect 3160 4826 3188 5063
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3620 4758 3648 5510
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3332 4616 3384 4622
rect 3238 4584 3294 4593
rect 3332 4558 3384 4564
rect 3238 4519 3294 4528
rect 3252 3602 3280 4519
rect 3344 4282 3372 4558
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3054 3496 3110 3505
rect 3054 3431 3110 3440
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 2310 2820 2450
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 2792 800 2820 2246
rect 3252 800 3280 3334
rect 3436 2990 3464 4218
rect 3528 4185 3556 4626
rect 3514 4176 3570 4185
rect 3514 4111 3570 4120
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3620 3058 3648 4014
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3528 2446 3556 2994
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3712 800 3740 7278
rect 3804 7002 3832 7686
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3896 6730 3924 12718
rect 4080 11626 4108 13670
rect 4724 13326 4752 14010
rect 4816 13920 4844 14368
rect 4896 13932 4948 13938
rect 4816 13892 4896 13920
rect 4896 13874 4948 13880
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4172 11286 4200 13126
rect 4264 12986 4292 13194
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4264 12442 4292 12582
rect 4448 12442 4476 12582
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4264 11898 4292 12378
rect 4632 12238 4660 12378
rect 4724 12374 4752 13126
rect 4816 12782 4844 13126
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4908 12714 4936 13874
rect 5000 13025 5028 14554
rect 4986 13016 5042 13025
rect 4986 12951 5042 12960
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 5000 12646 5028 12951
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 12102 4752 12174
rect 4908 12102 4936 12242
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 10266 4016 10542
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 3974 10024 4030 10033
rect 3974 9959 4030 9968
rect 3988 8945 4016 9959
rect 4080 9586 4108 10095
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3974 8936 4030 8945
rect 3974 8871 4030 8880
rect 4172 8514 4200 11086
rect 4080 8486 4200 8514
rect 4080 8242 4108 8486
rect 4264 8362 4292 11562
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4724 10130 4752 11494
rect 4802 11384 4858 11393
rect 4802 11319 4858 11328
rect 4816 10577 4844 11319
rect 4802 10568 4858 10577
rect 4802 10503 4858 10512
rect 4802 10432 4858 10441
rect 4802 10367 4858 10376
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4724 9586 4752 10066
rect 4816 10033 4844 10367
rect 4802 10024 4858 10033
rect 4802 9959 4858 9968
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4908 9058 4936 12038
rect 5000 11218 5028 12582
rect 5092 11354 5120 14826
rect 5184 14618 5212 20674
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5552 19242 5580 19858
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5644 18154 5672 19654
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 6276 19236 6328 19242
rect 6276 19178 6328 19184
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18630 5948 19110
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 6288 18358 6316 19178
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6276 18352 6328 18358
rect 6276 18294 6328 18300
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5460 15162 5488 15642
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13530 5212 13670
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5184 12986 5212 13466
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12986 5304 13262
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5276 12238 5304 12582
rect 5264 12232 5316 12238
rect 5184 12192 5264 12220
rect 5184 11694 5212 12192
rect 5264 12174 5316 12180
rect 5368 11744 5396 14758
rect 5552 13802 5580 17614
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5644 16726 5672 16934
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5644 15162 5672 16662
rect 6012 16046 6040 16934
rect 6104 16250 6132 17478
rect 6288 17134 6316 18022
rect 6564 17354 6592 18362
rect 7484 18222 7512 18566
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7484 17542 7512 18158
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17610 8248 18022
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 6472 17338 6592 17354
rect 6460 17332 6592 17338
rect 6512 17326 6592 17332
rect 6460 17274 6512 17280
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6104 16114 6132 16186
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13530 5580 13738
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5448 12776 5500 12782
rect 5446 12744 5448 12753
rect 5500 12744 5502 12753
rect 5446 12679 5502 12688
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5460 11898 5488 12310
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5276 11716 5396 11744
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 9926 5028 10474
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5170 9888 5226 9897
rect 5170 9823 5226 9832
rect 4988 9376 5040 9382
rect 5184 9364 5212 9823
rect 5276 9625 5304 11716
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 11286 5396 11562
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5368 10538 5396 11222
rect 5460 11082 5488 11834
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5262 9616 5318 9625
rect 5368 9586 5396 10474
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5552 9654 5580 10066
rect 5644 9654 5672 11222
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5262 9551 5318 9560
rect 5356 9580 5408 9586
rect 5040 9336 5212 9364
rect 4988 9318 5040 9324
rect 4804 9036 4856 9042
rect 4908 9030 5028 9058
rect 4804 8978 4856 8984
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4816 8242 4844 8978
rect 4080 8214 4200 8242
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3988 7274 4016 7958
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 3988 6934 4016 7103
rect 4080 7002 4108 7511
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 4066 6760 4122 6769
rect 3884 6724 3936 6730
rect 4066 6695 4122 6704
rect 3884 6666 3936 6672
rect 4080 6458 4108 6695
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 6236 4200 8214
rect 4724 8214 4844 8242
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4724 8090 4752 8214
rect 4908 8090 4936 8230
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4264 6440 4292 8026
rect 4894 7984 4950 7993
rect 4894 7919 4950 7928
rect 4908 7886 4936 7919
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4712 7744 4764 7750
rect 4816 7721 4844 7754
rect 4712 7686 4764 7692
rect 4802 7712 4858 7721
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4620 7472 4672 7478
rect 4724 7449 4752 7686
rect 4802 7647 4858 7656
rect 4710 7440 4766 7449
rect 4672 7420 4710 7426
rect 4620 7414 4710 7420
rect 4448 7041 4476 7414
rect 4632 7398 4710 7414
rect 4710 7375 4766 7384
rect 4434 7032 4490 7041
rect 4434 6967 4490 6976
rect 4448 6866 4476 6967
rect 4816 6866 4844 7647
rect 4908 7546 4936 7822
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4712 6792 4764 6798
rect 4710 6760 4712 6769
rect 4764 6760 4766 6769
rect 4710 6695 4766 6704
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4264 6412 4476 6440
rect 3882 6216 3938 6225
rect 4172 6208 4292 6236
rect 3882 6151 3938 6160
rect 3896 5846 3924 6151
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3988 5914 4016 6054
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3884 5840 3936 5846
rect 4080 5817 4108 6054
rect 3884 5782 3936 5788
rect 4066 5808 4122 5817
rect 4264 5778 4292 6208
rect 4066 5743 4122 5752
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4068 5704 4120 5710
rect 3974 5672 4030 5681
rect 4068 5646 4120 5652
rect 4160 5704 4212 5710
rect 4448 5658 4476 6412
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4160 5646 4212 5652
rect 3974 5607 4030 5616
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 4826 3832 5510
rect 3988 5030 4016 5607
rect 4080 5574 4108 5646
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4172 5302 4200 5646
rect 4264 5630 4476 5658
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4160 5296 4212 5302
rect 4066 5264 4122 5273
rect 4160 5238 4212 5244
rect 4066 5199 4122 5208
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3804 4622 3832 4762
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3804 4010 3832 4558
rect 3988 4486 4016 4966
rect 4080 4826 4108 5199
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 4080 4321 4108 4490
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3882 3632 3938 3641
rect 3804 2514 3832 3606
rect 3882 3567 3938 3576
rect 3896 2582 3924 3567
rect 3988 2650 4016 3946
rect 4080 3738 4108 4111
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 3194 4108 3470
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4172 3074 4200 5238
rect 4080 3046 4200 3074
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 4080 800 4108 3046
rect 4264 1442 4292 5630
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5234 4752 5646
rect 4908 5370 4936 5714
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4908 4282 4936 5034
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3777 4936 3878
rect 4894 3768 4950 3777
rect 4528 3732 4580 3738
rect 4894 3703 4950 3712
rect 4528 3674 4580 3680
rect 4540 3641 4568 3674
rect 4526 3632 4582 3641
rect 4526 3567 4582 3576
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4436 3120 4488 3126
rect 4724 3108 4752 3538
rect 4488 3097 4752 3108
rect 4488 3088 4766 3097
rect 4488 3080 4710 3088
rect 4436 3062 4488 3068
rect 4710 3023 4766 3032
rect 4620 2984 4672 2990
rect 4618 2952 4620 2961
rect 4672 2952 4674 2961
rect 4618 2887 4674 2896
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4448 2582 4476 2790
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1414 4568 1442
rect 4540 800 4568 1414
rect 5000 800 5028 9030
rect 5184 9024 5212 9336
rect 5276 9178 5304 9551
rect 5356 9522 5408 9528
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5368 9110 5396 9522
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5184 8996 5304 9024
rect 5080 8968 5132 8974
rect 5132 8928 5212 8956
rect 5080 8910 5132 8916
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 7410 5120 8774
rect 5184 8430 5212 8928
rect 5276 8786 5304 8996
rect 5276 8758 5396 8786
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5184 7886 5212 8366
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5092 7274 5120 7346
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5184 6730 5212 7686
rect 5276 7546 5304 8570
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 5184 5710 5212 6326
rect 5276 6254 5304 7482
rect 5368 7206 5396 8758
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 6798 5396 7142
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4622 5396 4966
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4457 5396 4558
rect 5354 4448 5410 4457
rect 5354 4383 5410 4392
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5092 2990 5120 4218
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3466 5396 3878
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5264 3392 5316 3398
rect 5262 3360 5264 3369
rect 5316 3360 5318 3369
rect 5262 3295 5318 3304
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5460 800 5488 9318
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8634 5580 8910
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5644 8294 5672 9114
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5630 7576 5686 7585
rect 5630 7511 5686 7520
rect 5644 7410 5672 7511
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5736 7290 5764 15914
rect 6012 15706 6040 15982
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5920 13394 5948 13466
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5828 7546 5856 13262
rect 5908 12640 5960 12646
rect 5906 12608 5908 12617
rect 6092 12640 6144 12646
rect 5960 12608 5962 12617
rect 6092 12582 6144 12588
rect 5906 12543 5962 12552
rect 6104 10690 6132 12582
rect 6288 11830 6316 17070
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6380 13326 6408 14486
rect 6564 14074 6592 17326
rect 6840 17270 6868 17478
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6656 15502 6684 17070
rect 6840 16794 6868 17206
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6840 16114 6868 16730
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7392 16114 7420 16662
rect 7484 16658 7512 17478
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7484 15978 7512 16390
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6656 14414 6684 15438
rect 6932 15026 6960 15506
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6656 13870 6684 14214
rect 7392 14074 7420 14214
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6656 12850 6684 13806
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6458 12608 6514 12617
rect 6458 12543 6514 12552
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10810 6224 11086
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6104 10662 6316 10690
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 10266 6040 10406
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6012 9654 6040 10202
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5920 8838 5948 9386
rect 5998 8936 6054 8945
rect 6104 8906 6132 9862
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 8906 6224 9318
rect 5998 8871 6054 8880
rect 6092 8900 6144 8906
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5552 7262 5764 7290
rect 5552 3126 5580 7262
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5644 5817 5672 6190
rect 5630 5808 5686 5817
rect 5630 5743 5632 5752
rect 5684 5743 5686 5752
rect 5632 5714 5684 5720
rect 5644 5683 5672 5714
rect 5736 5166 5764 6666
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 6254 5856 6598
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5644 4078 5672 4762
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5736 3924 5764 4626
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5828 4185 5856 4558
rect 5814 4176 5870 4185
rect 5814 4111 5870 4120
rect 5828 4010 5856 4111
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5644 3896 5764 3924
rect 5644 3482 5672 3896
rect 5644 3454 5764 3482
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5736 3058 5764 3454
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2582 5580 2790
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5920 800 5948 8774
rect 6012 8634 6040 8871
rect 6092 8842 6144 8848
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7478 6040 8230
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 6104 5778 6132 8842
rect 6196 8673 6224 8842
rect 6182 8664 6238 8673
rect 6182 8599 6238 8608
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6196 8022 6224 8434
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6196 7585 6224 7958
rect 6182 7576 6238 7585
rect 6182 7511 6238 7520
rect 6182 6896 6238 6905
rect 6182 6831 6238 6840
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6012 3670 6040 4558
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6012 2854 6040 3606
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6104 2650 6132 4558
rect 6196 4282 6224 6831
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6196 3398 6224 4218
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6288 800 6316 10662
rect 6366 9616 6422 9625
rect 6366 9551 6422 9560
rect 6380 6905 6408 9551
rect 6472 8566 6500 12543
rect 6656 12442 6684 12786
rect 6840 12646 6868 13670
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 7024 12374 7052 13330
rect 7116 12753 7144 13806
rect 7102 12744 7158 12753
rect 7102 12679 7158 12688
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11694 6868 12174
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 7024 11529 7052 12310
rect 7116 11898 7144 12679
rect 7300 12646 7328 13874
rect 7392 13394 7420 14010
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7286 12064 7342 12073
rect 7286 11999 7342 12008
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7300 11778 7328 11999
rect 7208 11750 7328 11778
rect 7010 11520 7066 11529
rect 7010 11455 7066 11464
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6840 11121 6868 11222
rect 6826 11112 6882 11121
rect 6826 11047 6882 11056
rect 6734 9208 6790 9217
rect 6734 9143 6790 9152
rect 6748 9110 6776 9143
rect 6736 9104 6788 9110
rect 6550 9072 6606 9081
rect 6736 9046 6788 9052
rect 6550 9007 6552 9016
rect 6604 9007 6606 9016
rect 6552 8978 6604 8984
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6472 8294 6500 8366
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6564 7868 6592 8978
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6748 8344 6776 8570
rect 6748 8316 6868 8344
rect 6840 8242 6868 8316
rect 6472 7840 6592 7868
rect 6656 8214 6868 8242
rect 6472 7750 6500 7840
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6366 6896 6422 6905
rect 6366 6831 6422 6840
rect 6656 6730 6684 8214
rect 6826 8120 6882 8129
rect 6826 8055 6882 8064
rect 6920 8084 6972 8090
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5166 6408 6054
rect 6642 5944 6698 5953
rect 6552 5908 6604 5914
rect 6642 5879 6698 5888
rect 6552 5850 6604 5856
rect 6458 5536 6514 5545
rect 6458 5471 6514 5480
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6380 4729 6408 4762
rect 6366 4720 6422 4729
rect 6366 4655 6422 4664
rect 6472 4622 6500 5471
rect 6564 4690 6592 5850
rect 6656 5681 6684 5879
rect 6642 5672 6698 5681
rect 6642 5607 6698 5616
rect 6656 5234 6684 5607
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6564 4010 6592 4626
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6564 3738 6592 3946
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6748 800 6776 7482
rect 6840 7410 6868 8055
rect 6920 8026 6972 8032
rect 6932 7721 6960 8026
rect 6918 7712 6974 7721
rect 6918 7647 6974 7656
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6932 6882 6960 7647
rect 6840 6866 6960 6882
rect 6828 6860 6960 6866
rect 6880 6854 6960 6860
rect 6828 6802 6880 6808
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7024 6746 7052 11290
rect 7208 10130 7236 11750
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7300 10266 7328 11630
rect 7392 11218 7420 13330
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7484 10690 7512 15914
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7392 10662 7512 10690
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7208 9654 7236 10066
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7116 8430 7144 9386
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 8022 7236 8230
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7300 7954 7328 10202
rect 7392 9353 7420 10662
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7484 9722 7512 10474
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7378 9344 7434 9353
rect 7378 9279 7434 9288
rect 7392 9178 7420 9279
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7102 7848 7158 7857
rect 7286 7848 7342 7857
rect 7102 7783 7158 7792
rect 7208 7806 7286 7834
rect 7116 7313 7144 7783
rect 7208 7750 7236 7806
rect 7286 7783 7342 7792
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7102 7304 7158 7313
rect 7102 7239 7158 7248
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6932 6322 6960 6734
rect 7024 6718 7144 6746
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6826 6216 6882 6225
rect 7024 6186 7052 6598
rect 7116 6322 7144 6718
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6826 6151 6882 6160
rect 7012 6180 7064 6186
rect 6840 6118 6868 6151
rect 7012 6122 7064 6128
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6920 6112 6972 6118
rect 6972 6060 7052 6066
rect 6920 6054 7052 6060
rect 6932 6038 7052 6054
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6826 5264 6882 5273
rect 6932 5234 6960 5714
rect 6826 5199 6882 5208
rect 6920 5228 6972 5234
rect 6840 4826 6868 5199
rect 6920 5170 6972 5176
rect 7024 5098 7052 6038
rect 7116 5914 7144 6258
rect 7208 6254 7236 7142
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7300 6168 7328 7686
rect 7392 6662 7420 8230
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7484 7478 7512 7822
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7380 6180 7432 6186
rect 7300 6140 7380 6168
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7116 5778 7144 5850
rect 7300 5846 7328 6140
rect 7380 6122 7432 6128
rect 7484 6118 7512 6802
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7288 5840 7340 5846
rect 7194 5808 7250 5817
rect 7104 5772 7156 5778
rect 7288 5782 7340 5788
rect 7194 5743 7250 5752
rect 7104 5714 7156 5720
rect 7208 5710 7236 5743
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6840 4486 6868 4762
rect 7116 4758 7144 4966
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 7024 4196 7052 4626
rect 7208 4282 7236 5646
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 6932 4168 7052 4196
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6840 3602 6868 4082
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6932 2689 6960 4168
rect 7102 3768 7158 3777
rect 7102 3703 7158 3712
rect 6918 2680 6974 2689
rect 6918 2615 6974 2624
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6932 1970 6960 2246
rect 7024 2038 7052 2518
rect 7116 2514 7144 3703
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 7208 800 7236 3062
rect 7300 2961 7328 4966
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3126 7512 3334
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7286 2952 7342 2961
rect 7286 2887 7342 2896
rect 7484 2854 7512 3062
rect 7288 2848 7340 2854
rect 7472 2848 7524 2854
rect 7340 2796 7420 2802
rect 7288 2790 7420 2796
rect 7472 2790 7524 2796
rect 7300 2774 7420 2790
rect 7392 2650 7420 2774
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7392 2553 7420 2586
rect 7378 2544 7434 2553
rect 7378 2479 7434 2488
rect 7576 1442 7604 15846
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15026 8248 16934
rect 8312 16794 8340 18022
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8588 16658 8616 16934
rect 8772 16794 8800 17478
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8680 15162 8708 15574
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8772 15162 8800 15506
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7668 1578 7696 14758
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14618 8248 14962
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8312 14074 8340 14894
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8312 13802 8340 13874
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8404 13258 8432 14214
rect 8496 13870 8524 14758
rect 8864 14634 8892 15438
rect 8772 14606 8892 14634
rect 8772 14550 8800 14606
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8772 14278 8800 14486
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 14074 8800 14214
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8956 14006 8984 18634
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13394 8524 13670
rect 8588 13530 8616 13874
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8114 13016 8170 13025
rect 8114 12951 8170 12960
rect 8128 12628 8156 12951
rect 8404 12850 8432 13194
rect 8680 13190 8708 13670
rect 8484 13184 8536 13190
rect 8668 13184 8720 13190
rect 8536 13132 8616 13138
rect 8484 13126 8616 13132
rect 8668 13126 8720 13132
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8496 13110 8616 13126
rect 8588 12918 8616 13110
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8208 12776 8260 12782
rect 8484 12776 8536 12782
rect 8260 12736 8340 12764
rect 8208 12718 8260 12724
rect 8312 12646 8340 12736
rect 8484 12718 8536 12724
rect 8208 12640 8260 12646
rect 8128 12600 8208 12628
rect 8208 12582 8260 12588
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8220 12238 8248 12582
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7852 11626 7880 11834
rect 7932 11688 7984 11694
rect 7930 11656 7932 11665
rect 7984 11656 7986 11665
rect 7840 11620 7892 11626
rect 7760 11580 7840 11608
rect 7760 10810 7788 11580
rect 7930 11591 7986 11600
rect 7840 11562 7892 11568
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 8128 10554 8156 11222
rect 8220 11218 8248 12038
rect 8312 11665 8340 12242
rect 8298 11656 8354 11665
rect 8298 11591 8354 11600
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 10674 8248 11154
rect 8300 10736 8352 10742
rect 8404 10724 8432 11562
rect 8352 10696 8432 10724
rect 8300 10678 8352 10684
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8128 10526 8248 10554
rect 8220 10470 8248 10526
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7760 9908 7788 10406
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7840 9920 7892 9926
rect 7760 9888 7840 9908
rect 7892 9888 7894 9897
rect 7760 9880 7838 9888
rect 7838 9823 7894 9832
rect 7838 9616 7894 9625
rect 7838 9551 7840 9560
rect 7892 9551 7894 9560
rect 7840 9522 7892 9528
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 9058 7788 9318
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7760 9030 7972 9058
rect 7944 8634 7972 9030
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8220 8294 8248 10406
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 9178 8340 9454
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8566 8340 8978
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8496 8072 8524 12718
rect 8680 12481 8708 13126
rect 8956 12782 8984 13126
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8666 12472 8722 12481
rect 8666 12407 8722 12416
rect 8680 12374 8708 12407
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 9048 11898 9076 19246
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 18222 9260 18566
rect 9416 18290 9444 18702
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9876 17882 9904 18158
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9140 16726 9168 17546
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9140 16250 9168 16662
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9140 14958 9168 16186
rect 9324 15706 9352 16594
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 15910 9444 16458
rect 9600 16114 9628 16934
rect 9692 16726 9720 17070
rect 10152 17066 10180 18022
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10244 17338 10272 17682
rect 10336 17678 10364 18022
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 10152 16794 10180 17002
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9692 16590 9720 16662
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9784 16250 9812 16730
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9968 16454 9996 16594
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9968 16182 9996 16390
rect 10336 16250 10364 17614
rect 11164 17338 11192 17614
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 11072 16114 11100 16730
rect 11624 16658 11652 17274
rect 11716 16794 11744 18022
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11624 16250 11652 16594
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9968 14958 9996 15438
rect 9128 14952 9180 14958
rect 9956 14952 10008 14958
rect 9180 14912 9536 14940
rect 9128 14894 9180 14900
rect 9508 14006 9536 14912
rect 9956 14894 10008 14900
rect 10060 14618 10088 15506
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10428 14550 10456 15506
rect 10520 15162 10548 16050
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15366 10732 15846
rect 11164 15706 11192 15914
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10612 15042 10640 15098
rect 10520 15026 10640 15042
rect 10508 15020 10640 15026
rect 10560 15014 10640 15020
rect 10508 14962 10560 14968
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9416 13790 9720 13818
rect 9416 13462 9444 13790
rect 9692 13569 9720 13790
rect 9772 13728 9824 13734
rect 9770 13696 9772 13705
rect 9824 13696 9826 13705
rect 9770 13631 9826 13640
rect 9678 13560 9734 13569
rect 9678 13495 9734 13504
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9770 13424 9826 13433
rect 9770 13359 9826 13368
rect 9784 13326 9812 13359
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12782 9812 13262
rect 9772 12776 9824 12782
rect 9126 12744 9182 12753
rect 9772 12718 9824 12724
rect 9126 12679 9182 12688
rect 9140 12238 9168 12679
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8574 10432 8630 10441
rect 8574 10367 8630 10376
rect 8588 10266 8616 10367
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8588 8974 8616 9522
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8566 8616 8910
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8576 8424 8628 8430
rect 8574 8392 8576 8401
rect 8628 8392 8630 8401
rect 8574 8327 8630 8336
rect 8404 8044 8524 8072
rect 8298 7984 8354 7993
rect 8298 7919 8354 7928
rect 7748 7744 7800 7750
rect 8024 7744 8076 7750
rect 7748 7686 7800 7692
rect 8022 7712 8024 7721
rect 8076 7712 8078 7721
rect 7760 7256 7788 7686
rect 8022 7647 8078 7656
rect 7932 7268 7984 7274
rect 7760 7228 7932 7256
rect 7760 6798 7788 7228
rect 8024 7268 8076 7274
rect 7984 7228 8024 7256
rect 7932 7210 7984 7216
rect 8024 7210 8076 7216
rect 8312 7177 8340 7919
rect 8404 7868 8432 8044
rect 8404 7840 8524 7868
rect 8298 7168 8354 7177
rect 7820 7100 8116 7120
rect 8298 7103 8354 7112
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7760 5778 7788 6122
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7760 4808 7788 5170
rect 8220 5114 8248 6598
rect 8392 5840 8444 5846
rect 8298 5808 8354 5817
rect 8392 5782 8444 5788
rect 8298 5743 8354 5752
rect 8312 5710 8340 5743
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8404 5166 8432 5782
rect 8392 5160 8444 5166
rect 8220 5086 8340 5114
rect 8392 5102 8444 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7760 4780 7972 4808
rect 7944 4622 7972 4780
rect 8220 4622 8248 4966
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7746 4448 7802 4457
rect 7746 4383 7802 4392
rect 7760 3670 7788 4383
rect 7852 4078 7880 4558
rect 7944 4282 7972 4558
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 8312 4010 8340 5086
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8404 4826 8432 4966
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7760 3058 7788 3402
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7760 2446 7788 2994
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 2514 8248 3606
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8390 3360 8446 3369
rect 8312 3058 8340 3334
rect 8390 3295 8446 3304
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8312 2650 8340 2994
rect 8404 2922 8432 3295
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 2106 8248 2246
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 7668 1550 8064 1578
rect 7576 1414 7696 1442
rect 7668 800 7696 1414
rect 8036 800 8064 1550
rect 8496 800 8524 7840
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 5846 8616 6598
rect 8680 6186 8708 9862
rect 8772 9518 8800 11494
rect 9140 11286 9168 11698
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9140 11150 9168 11222
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 10606 9168 11086
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 9034 10024 9090 10033
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8772 8294 8800 8842
rect 8864 8401 8892 9998
rect 9034 9959 9036 9968
rect 9088 9959 9090 9968
rect 9036 9930 9088 9936
rect 9140 9926 9168 10406
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9036 9104 9088 9110
rect 9088 9064 9168 9092
rect 9036 9046 9088 9052
rect 9034 8800 9090 8809
rect 9034 8735 9090 8744
rect 8850 8392 8906 8401
rect 8850 8327 8906 8336
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8864 8090 8892 8327
rect 9048 8294 9076 8735
rect 9140 8480 9168 9064
rect 9232 8922 9260 9318
rect 9324 9178 9352 12582
rect 9876 12442 9904 13874
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9968 13433 9996 13738
rect 10060 13462 10088 13874
rect 10152 13870 10180 14214
rect 10244 14006 10272 14214
rect 10232 14000 10284 14006
rect 10336 13977 10364 14350
rect 10428 14090 10456 14486
rect 10612 14385 10640 14758
rect 10598 14376 10654 14385
rect 10598 14311 10654 14320
rect 10428 14074 10548 14090
rect 10428 14068 10560 14074
rect 10428 14062 10508 14068
rect 10508 14010 10560 14016
rect 10232 13942 10284 13948
rect 10322 13968 10378 13977
rect 10322 13903 10378 13912
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10152 13530 10180 13806
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10048 13456 10100 13462
rect 9954 13424 10010 13433
rect 10048 13398 10100 13404
rect 9954 13359 10010 13368
rect 9968 12566 10272 12594
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9968 12374 9996 12566
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9416 11558 9444 12038
rect 9784 11830 9812 12038
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9678 11520 9734 11529
rect 9416 11354 9444 11494
rect 9678 11455 9734 11464
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9692 11286 9720 11455
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9680 11144 9732 11150
rect 9784 11098 9812 11766
rect 9732 11092 9812 11098
rect 9680 11086 9812 11092
rect 9692 11070 9812 11086
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9232 8894 9352 8922
rect 9324 8566 9352 8894
rect 9416 8673 9444 9318
rect 9402 8664 9458 8673
rect 9402 8599 9458 8608
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9220 8492 9272 8498
rect 9140 8452 9220 8480
rect 9220 8434 9272 8440
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 9048 7954 9260 7970
rect 9036 7948 9272 7954
rect 9088 7942 9220 7948
rect 9036 7890 9088 7896
rect 9220 7890 9272 7896
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9048 7546 9076 7754
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7546 9168 7686
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8574 5672 8630 5681
rect 8680 5658 8708 6122
rect 8956 5914 8984 6802
rect 9048 6798 9076 7482
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9232 6118 9260 7346
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9324 6798 9352 7210
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9416 6390 9444 7210
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8630 5630 8708 5658
rect 8574 5607 8630 5616
rect 8588 5574 8616 5607
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8588 4486 8616 4626
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8576 4480 8628 4486
rect 8574 4448 8576 4457
rect 8628 4448 8630 4457
rect 8574 4383 8630 4392
rect 8772 4078 8800 4490
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9048 4282 9076 4422
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9048 4146 9076 4218
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9324 4078 9352 5510
rect 9508 4842 9536 10406
rect 9600 9568 9628 10950
rect 9692 10470 9720 10950
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9784 9926 9812 11070
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9680 9580 9732 9586
rect 9600 9540 9680 9568
rect 9680 9522 9732 9528
rect 9784 9466 9812 9862
rect 9692 9438 9812 9466
rect 9692 8974 9720 9438
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 8968 9732 8974
rect 9784 8945 9812 9318
rect 9680 8910 9732 8916
rect 9770 8936 9826 8945
rect 9692 8362 9720 8910
rect 9770 8871 9826 8880
rect 9876 8362 9904 12242
rect 10060 12238 10088 12378
rect 10244 12374 10272 12566
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10046 11384 10102 11393
rect 10046 11319 10102 11328
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9968 10742 9996 11222
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 10060 10538 10088 11319
rect 10152 10690 10180 12174
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10244 10810 10272 11834
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10152 10662 10272 10690
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 8945 9996 9862
rect 10244 9194 10272 10662
rect 10336 9926 10364 13738
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10152 9166 10272 9194
rect 9954 8936 10010 8945
rect 9954 8871 10010 8880
rect 9954 8664 10010 8673
rect 9954 8599 10010 8608
rect 9968 8430 9996 8599
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9692 7886 9720 8298
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9876 7818 9904 8298
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9600 7274 9628 7754
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 6118 9628 6258
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9770 6080 9826 6089
rect 9600 5166 9628 6054
rect 9770 6015 9826 6024
rect 9678 5944 9734 5953
rect 9784 5914 9812 6015
rect 9678 5879 9734 5888
rect 9772 5908 9824 5914
rect 9692 5710 9720 5879
rect 9772 5850 9824 5856
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9784 5166 9812 5714
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9416 4814 9536 4842
rect 9600 4826 9628 5102
rect 9588 4820 9640 4826
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 8588 3670 8616 4014
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8666 3224 8722 3233
rect 8666 3159 8722 3168
rect 8680 3126 8708 3159
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8772 2990 8800 3538
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8588 2825 8616 2926
rect 8574 2816 8630 2825
rect 8574 2751 8630 2760
rect 8956 800 8984 3946
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 2446 9168 3878
rect 9324 3534 9352 4014
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 2922 9352 3470
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9140 1834 9168 2382
rect 9128 1828 9180 1834
rect 9128 1770 9180 1776
rect 9416 800 9444 4814
rect 9588 4762 9640 4768
rect 9586 4720 9642 4729
rect 9586 4655 9642 4664
rect 9600 4321 9628 4655
rect 9586 4312 9642 4321
rect 9586 4247 9642 4256
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9692 2854 9720 3674
rect 9784 2990 9812 3878
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9680 2848 9732 2854
rect 9876 2836 9904 6802
rect 9968 6322 9996 6938
rect 10152 6866 10180 9166
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10244 8498 10272 9046
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10140 6860 10192 6866
rect 10428 6848 10456 13670
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10520 12238 10548 12650
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10506 10704 10562 10713
rect 10506 10639 10562 10648
rect 10520 10606 10548 10639
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10612 10441 10640 10542
rect 10598 10432 10654 10441
rect 10598 10367 10654 10376
rect 10612 9450 10640 10367
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10520 7478 10548 7890
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10140 6802 10192 6808
rect 10244 6820 10456 6848
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9956 5772 10008 5778
rect 10060 5760 10088 6326
rect 10008 5732 10088 5760
rect 9956 5714 10008 5720
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9954 5128 10010 5137
rect 9954 5063 9956 5072
rect 10008 5063 10010 5072
rect 9956 5034 10008 5040
rect 10060 4826 10088 5578
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3738 9996 4014
rect 10060 3738 10088 4762
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9680 2790 9732 2796
rect 9784 2808 9904 2836
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9692 2378 9720 2450
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9784 800 9812 2808
rect 9968 2582 9996 3334
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10060 2514 10088 3674
rect 10152 3194 10180 6598
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10152 2446 10180 3130
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10244 800 10272 6820
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6254 10456 6666
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10428 3233 10456 5714
rect 10520 5710 10548 7142
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10520 4826 10548 5034
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10508 3936 10560 3942
rect 10612 3913 10640 8366
rect 10508 3878 10560 3884
rect 10598 3904 10654 3913
rect 10414 3224 10470 3233
rect 10414 3159 10470 3168
rect 10520 2378 10548 3878
rect 10598 3839 10654 3848
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10612 2650 10640 2790
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 10612 2417 10640 2586
rect 10598 2408 10654 2417
rect 10508 2372 10560 2378
rect 10598 2343 10654 2352
rect 10508 2314 10560 2320
rect 10704 800 10732 15302
rect 10980 14958 11008 15438
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14618 10824 14758
rect 10980 14618 11008 14894
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11072 13938 11100 14418
rect 11808 14414 11836 17750
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12452 17134 12480 17546
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17134 12756 17478
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12452 16454 12480 17070
rect 12728 16522 12756 17070
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11900 15162 11928 15506
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11888 14816 11940 14822
rect 11992 14804 12020 15438
rect 11940 14776 12020 14804
rect 11888 14758 11940 14764
rect 11796 14408 11848 14414
rect 11164 14346 11376 14362
rect 11796 14350 11848 14356
rect 11164 14340 11388 14346
rect 11164 14334 11336 14340
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11072 13530 11100 13874
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10796 12073 10824 13194
rect 10980 12986 11008 13398
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10874 12880 10930 12889
rect 10874 12815 10876 12824
rect 10928 12815 10930 12824
rect 10876 12786 10928 12792
rect 11164 12594 11192 14334
rect 11336 14282 11388 14288
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11624 12986 11652 13126
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 10980 12566 11192 12594
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10782 12064 10838 12073
rect 10782 11999 10838 12008
rect 10888 11558 10916 12378
rect 10980 12102 11008 12566
rect 11058 12472 11114 12481
rect 11058 12407 11060 12416
rect 11112 12407 11114 12416
rect 11610 12472 11666 12481
rect 11900 12458 11928 14758
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11992 13802 12020 14418
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11992 12646 12020 13398
rect 12256 13252 12308 13258
rect 12176 13212 12256 13240
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11900 12430 12020 12458
rect 11610 12407 11666 12416
rect 11060 12378 11112 12384
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 11778 11100 12038
rect 10980 11750 11100 11778
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10796 11218 10824 11494
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10538 10824 10950
rect 10980 10792 11008 11750
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11072 11082 11100 11630
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10980 10764 11100 10792
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 11072 10180 11100 10764
rect 11164 10452 11192 12242
rect 11624 12170 11652 12407
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11716 11830 11744 12174
rect 11796 12096 11848 12102
rect 11848 12056 11928 12084
rect 11796 12038 11848 12044
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11256 11121 11284 11766
rect 11242 11112 11298 11121
rect 11242 11047 11298 11056
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11244 10464 11296 10470
rect 11164 10424 11244 10452
rect 11244 10406 11296 10412
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11072 10152 11192 10180
rect 10968 10124 11020 10130
rect 11020 10084 11100 10112
rect 10968 10066 11020 10072
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 9110 11008 9522
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10782 8936 10838 8945
rect 10980 8906 11008 9046
rect 10782 8871 10838 8880
rect 10968 8900 11020 8906
rect 10796 8838 10824 8871
rect 10968 8842 11020 8848
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10888 8673 10916 8774
rect 10874 8664 10930 8673
rect 10874 8599 10930 8608
rect 10782 8528 10838 8537
rect 10782 8463 10838 8472
rect 10796 5896 10824 8463
rect 10966 8392 11022 8401
rect 11072 8362 11100 10084
rect 11164 9704 11192 10152
rect 11256 10062 11284 10406
rect 11348 10169 11376 10406
rect 11334 10160 11390 10169
rect 11334 10095 11390 10104
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11164 9676 11468 9704
rect 11152 9512 11204 9518
rect 11204 9460 11376 9466
rect 11152 9454 11376 9460
rect 11164 9438 11376 9454
rect 11348 9382 11376 9438
rect 11336 9376 11388 9382
rect 11150 9344 11206 9353
rect 11336 9318 11388 9324
rect 11150 9279 11206 9288
rect 11164 8634 11192 9279
rect 11440 8974 11468 9676
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11532 8906 11560 9454
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8634 11652 10542
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11808 9926 11836 10202
rect 11900 10130 11928 12056
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11796 9920 11848 9926
rect 11794 9888 11796 9897
rect 11848 9888 11850 9897
rect 11794 9823 11850 9832
rect 11702 9616 11758 9625
rect 11702 9551 11758 9560
rect 11716 9042 11744 9551
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 10966 8327 11022 8336
rect 11060 8356 11112 8362
rect 10874 7984 10930 7993
rect 10874 7919 10930 7928
rect 10888 7585 10916 7919
rect 10874 7576 10930 7585
rect 10874 7511 10930 7520
rect 10980 7002 11008 8327
rect 11060 8298 11112 8304
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10980 6798 11008 6938
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10796 5868 10916 5896
rect 10782 5808 10838 5817
rect 10782 5743 10838 5752
rect 10796 5030 10824 5743
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10888 4146 10916 5868
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10980 4758 11008 5238
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11072 4706 11100 8298
rect 11610 7848 11666 7857
rect 11610 7783 11666 7792
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11244 7200 11296 7206
rect 11624 7177 11652 7783
rect 11716 7206 11744 8842
rect 11808 8430 11836 9823
rect 11900 9042 11928 10066
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11886 8256 11942 8265
rect 11886 8191 11942 8200
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11704 7200 11756 7206
rect 11244 7142 11296 7148
rect 11610 7168 11666 7177
rect 11256 6934 11284 7142
rect 11704 7142 11756 7148
rect 11610 7103 11666 7112
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11624 6866 11652 6938
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11150 6080 11206 6089
rect 11150 6015 11206 6024
rect 11164 5914 11192 6015
rect 11256 5914 11284 6122
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11164 5352 11192 5850
rect 11256 5710 11284 5850
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11164 5324 11284 5352
rect 11256 5030 11284 5324
rect 11624 5234 11652 5510
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11164 4826 11192 4966
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11072 4678 11192 4706
rect 10966 4448 11022 4457
rect 10966 4383 11022 4392
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10796 2310 10824 3946
rect 10888 3942 10916 4082
rect 10980 4010 11008 4383
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10888 2854 10916 3334
rect 10980 3058 11008 3470
rect 11058 3224 11114 3233
rect 11058 3159 11114 3168
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11072 2854 11100 3159
rect 11164 3126 11192 4678
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11440 3738 11468 4150
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 10876 2848 10928 2854
rect 10874 2816 10876 2825
rect 11060 2848 11112 2854
rect 10928 2816 10930 2825
rect 11060 2790 11112 2796
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 10874 2751 10930 2760
rect 11072 2650 11100 2790
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 2038 10824 2246
rect 11072 2106 11100 2382
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 10784 2032 10836 2038
rect 10784 1974 10836 1980
rect 11164 800 11192 2790
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11624 800 11652 4150
rect 11716 3398 11744 7142
rect 11808 7002 11836 7686
rect 11900 7585 11928 8191
rect 11886 7576 11942 7585
rect 11886 7511 11942 7520
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11900 7002 11928 7414
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11794 6488 11850 6497
rect 11794 6423 11850 6432
rect 11808 5846 11836 6423
rect 11886 6352 11942 6361
rect 11886 6287 11942 6296
rect 11900 6118 11928 6287
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11992 4842 12020 12430
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11694 12112 12106
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12072 11552 12124 11558
rect 12070 11520 12072 11529
rect 12124 11520 12126 11529
rect 12070 11455 12126 11464
rect 12084 11354 12112 11455
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12072 10464 12124 10470
rect 12070 10432 12072 10441
rect 12124 10432 12126 10441
rect 12070 10367 12126 10376
rect 12176 10305 12204 13212
rect 12256 13194 12308 13200
rect 12360 11744 12388 15846
rect 12728 15570 12756 16458
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 13096 15366 13124 16390
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12438 13968 12494 13977
rect 12438 13903 12494 13912
rect 12452 13802 12480 13903
rect 13096 13802 13124 15302
rect 13280 15162 13308 17614
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 13820 17264 13872 17270
rect 17960 17264 18012 17270
rect 13820 17206 13872 17212
rect 17958 17232 17960 17241
rect 18012 17232 18014 17241
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13372 16114 13400 16594
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13740 15910 13768 16594
rect 13832 16590 13860 17206
rect 17958 17167 18014 17176
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13832 16250 13860 16526
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15706 13768 15846
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13280 14618 13308 15098
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13280 14074 13308 14554
rect 13358 14376 13414 14385
rect 13358 14311 13414 14320
rect 14464 14340 14516 14346
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13372 14006 13400 14311
rect 14464 14282 14516 14288
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12452 12102 12480 13738
rect 12992 13728 13044 13734
rect 12530 13696 12586 13705
rect 12992 13670 13044 13676
rect 12530 13631 12586 13640
rect 12544 13530 12572 13631
rect 12898 13560 12954 13569
rect 12532 13524 12584 13530
rect 12898 13495 12900 13504
rect 12532 13466 12584 13472
rect 12952 13495 12954 13504
rect 12900 13466 12952 13472
rect 13004 13394 13032 13670
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13372 12968 13400 13942
rect 13740 13734 13768 14214
rect 14476 14074 14504 14282
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 14292 13530 14320 14010
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 15212 13190 15240 13670
rect 15488 13530 15516 14010
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 13452 12980 13504 12986
rect 13372 12940 13452 12968
rect 13452 12922 13504 12928
rect 15212 12646 15240 13126
rect 15304 12986 15332 13466
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 12636 12442 12664 12582
rect 12714 12472 12770 12481
rect 12624 12436 12676 12442
rect 12714 12407 12716 12416
rect 12624 12378 12676 12384
rect 12768 12407 12770 12416
rect 12716 12378 12768 12384
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12268 11716 12388 11744
rect 12162 10296 12218 10305
rect 12162 10231 12218 10240
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12084 8634 12112 9930
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12084 7954 12112 8366
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 7410 12112 7890
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12176 6202 12204 7414
rect 12268 7188 12296 11716
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12360 11529 12388 11562
rect 12544 11529 12572 12038
rect 12636 11830 12664 12378
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12346 11520 12402 11529
rect 12346 11455 12402 11464
rect 12530 11520 12586 11529
rect 12530 11455 12586 11464
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12360 7478 12388 11154
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10130 12480 11018
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9586 12480 10066
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12636 9178 12664 10474
rect 12820 9704 12848 12174
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 10742 13124 11494
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10266 13032 10406
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12820 9676 12940 9704
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9178 12756 9318
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12820 8498 12848 9386
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12268 7160 12388 7188
rect 12084 6174 12204 6202
rect 12084 5137 12112 6174
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 5681 12204 6054
rect 12162 5672 12218 5681
rect 12162 5607 12218 5616
rect 12070 5128 12126 5137
rect 12070 5063 12126 5072
rect 11808 4814 12020 4842
rect 11808 4214 11836 4814
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11992 4457 12020 4626
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 11978 4448 12034 4457
rect 11978 4383 12034 4392
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11886 3904 11942 3913
rect 11808 3670 11836 3878
rect 11886 3839 11942 3848
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11900 3482 11928 3839
rect 11992 3602 12020 4383
rect 12084 4146 12112 4490
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12176 4026 12204 5607
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12268 5030 12296 5102
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12084 3998 12204 4026
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 12084 3534 12112 3998
rect 12072 3528 12124 3534
rect 11900 3454 12020 3482
rect 12072 3470 12124 3476
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11808 2106 11836 3062
rect 11900 2922 11928 3062
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11900 2650 11928 2858
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11992 800 12020 3454
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12084 2514 12112 2586
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12176 2446 12204 3334
rect 12360 2854 12388 7160
rect 12544 6934 12572 8298
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 7546 12756 7686
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12532 6928 12584 6934
rect 12636 6905 12664 7414
rect 12820 7342 12848 7822
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12532 6870 12584 6876
rect 12622 6896 12678 6905
rect 12440 6860 12492 6866
rect 12622 6831 12678 6840
rect 12440 6802 12492 6808
rect 12452 6322 12480 6802
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12544 6361 12572 6666
rect 12530 6352 12586 6361
rect 12440 6316 12492 6322
rect 12530 6287 12586 6296
rect 12440 6258 12492 6264
rect 12452 4978 12480 6258
rect 12532 6248 12584 6254
rect 12584 6196 12756 6202
rect 12532 6190 12756 6196
rect 12544 6186 12756 6190
rect 12544 6180 12768 6186
rect 12544 6174 12716 6180
rect 12716 6122 12768 6128
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12716 5840 12768 5846
rect 12820 5817 12848 5850
rect 12716 5782 12768 5788
rect 12806 5808 12862 5817
rect 12622 5672 12678 5681
rect 12622 5607 12678 5616
rect 12636 5166 12664 5607
rect 12728 5234 12756 5782
rect 12806 5743 12862 5752
rect 12912 5642 12940 9676
rect 13004 9586 13032 10202
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13004 9110 13032 9522
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13096 7970 13124 9862
rect 13188 9353 13216 12582
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15488 12442 15516 13466
rect 16408 12646 16436 13738
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13556 11898 13584 12038
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13728 11688 13780 11694
rect 13726 11656 13728 11665
rect 13780 11656 13782 11665
rect 13636 11620 13688 11626
rect 13726 11591 13782 11600
rect 13636 11562 13688 11568
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13372 10810 13400 11018
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 10130 13308 10406
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13174 9344 13230 9353
rect 13174 9279 13230 9288
rect 13280 9110 13308 10066
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13096 7942 13216 7970
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13004 6186 13032 7686
rect 13096 7410 13124 7686
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13004 5914 13032 6122
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13004 5710 13032 5850
rect 13096 5846 13124 6598
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12452 4950 12572 4978
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 12452 2990 12480 4791
rect 12544 4214 12572 4950
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 13188 3670 13216 7942
rect 13280 7410 13308 8230
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13280 5574 13308 5850
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12636 2650 12664 3606
rect 13280 2990 13308 5510
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13372 2922 13400 9862
rect 13464 9489 13492 11494
rect 13648 11257 13676 11562
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13634 11248 13690 11257
rect 13740 11218 13768 11494
rect 13634 11183 13690 11192
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10470 13584 10950
rect 13832 10713 13860 12038
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13818 10704 13874 10713
rect 13818 10639 13874 10648
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13450 9480 13506 9489
rect 13450 9415 13506 9424
rect 13450 9344 13506 9353
rect 13450 9279 13506 9288
rect 13464 9042 13492 9279
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13556 8838 13584 10406
rect 13740 10062 13768 10406
rect 13728 10056 13780 10062
rect 13634 10024 13690 10033
rect 13728 9998 13780 10004
rect 13634 9959 13690 9968
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13464 8430 13492 8570
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 6866 13584 7278
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13450 6624 13506 6633
rect 13450 6559 13506 6568
rect 13464 6458 13492 6559
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13450 6352 13506 6361
rect 13450 6287 13506 6296
rect 13464 3194 13492 6287
rect 13648 5914 13676 9959
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 9353 13860 9454
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8566 13860 8978
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13924 8242 13952 11086
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14016 10606 14044 10950
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13832 8214 13952 8242
rect 13832 7426 13860 8214
rect 13740 7398 13860 7426
rect 13740 7018 13768 7398
rect 14016 7290 14044 9998
rect 14108 8498 14136 11494
rect 14292 11393 14320 12106
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11626 15424 12038
rect 15580 11898 15608 12242
rect 15856 12170 15884 12582
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14278 11384 14334 11393
rect 14684 11376 14980 11396
rect 14278 11319 14334 11328
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 10033 14228 10610
rect 14186 10024 14242 10033
rect 14186 9959 14242 9968
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14200 9518 14228 9862
rect 14292 9625 14320 9862
rect 14278 9616 14334 9625
rect 14278 9551 14334 9560
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 9178 14228 9454
rect 14384 9382 14412 11018
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14280 8560 14332 8566
rect 14186 8528 14242 8537
rect 14096 8492 14148 8498
rect 14280 8502 14332 8508
rect 14186 8463 14188 8472
rect 14096 8434 14148 8440
rect 14240 8463 14242 8472
rect 14188 8434 14240 8440
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14108 7818 14136 8230
rect 14186 8120 14242 8129
rect 14292 8090 14320 8502
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14186 8055 14242 8064
rect 14280 8084 14332 8090
rect 14200 7954 14228 8055
rect 14280 8026 14332 8032
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14186 7712 14242 7721
rect 14186 7647 14242 7656
rect 14200 7342 14228 7647
rect 13832 7262 14044 7290
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14278 7304 14334 7313
rect 13832 7206 13860 7262
rect 14278 7239 14334 7248
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13740 6990 13952 7018
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13740 5953 13768 6190
rect 13726 5944 13782 5953
rect 13636 5908 13688 5914
rect 13726 5879 13782 5888
rect 13636 5850 13688 5856
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13556 5681 13584 5714
rect 13728 5704 13780 5710
rect 13542 5672 13598 5681
rect 13728 5646 13780 5652
rect 13542 5607 13598 5616
rect 13542 4856 13598 4865
rect 13542 4791 13598 4800
rect 13556 4185 13584 4791
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13542 4176 13598 4185
rect 13542 4111 13598 4120
rect 13648 4078 13676 4422
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13542 3632 13598 3641
rect 13542 3567 13598 3576
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12728 2514 12756 2858
rect 13464 2582 13492 3130
rect 13556 3097 13584 3567
rect 13648 3534 13676 4014
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13542 3088 13598 3097
rect 13542 3023 13598 3032
rect 13740 2632 13768 5646
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13832 5273 13860 5306
rect 13818 5264 13874 5273
rect 13818 5199 13874 5208
rect 13820 4480 13872 4486
rect 13924 4457 13952 6990
rect 14016 6866 14044 7142
rect 14292 7041 14320 7239
rect 14278 7032 14334 7041
rect 14278 6967 14334 6976
rect 14094 6896 14150 6905
rect 14004 6860 14056 6866
rect 14094 6831 14096 6840
rect 14004 6802 14056 6808
rect 14148 6831 14150 6840
rect 14096 6802 14148 6808
rect 14016 6322 14044 6802
rect 14278 6624 14334 6633
rect 14278 6559 14334 6568
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14292 6186 14320 6559
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14096 6112 14148 6118
rect 14384 6066 14412 8366
rect 14096 6054 14148 6060
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14016 5166 14044 5850
rect 14108 5710 14136 6054
rect 14200 6038 14412 6066
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 14200 4978 14228 6038
rect 14476 5896 14504 10678
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15028 10266 15056 10542
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14648 9512 14700 9518
rect 14646 9480 14648 9489
rect 14700 9480 14702 9489
rect 14646 9415 14702 9424
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 9042 14596 9318
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15028 9058 15056 9522
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14844 9030 15056 9058
rect 14844 8430 14872 9030
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15028 8634 15056 8842
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 15028 8294 15056 8570
rect 15120 8548 15148 9114
rect 15212 9081 15240 11494
rect 15396 11218 15424 11562
rect 15580 11354 15608 11834
rect 16408 11626 16436 12038
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15198 9072 15254 9081
rect 15198 9007 15254 9016
rect 15200 8560 15252 8566
rect 15120 8520 15200 8548
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15120 8090 15148 8520
rect 15200 8502 15252 8508
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15304 7818 15332 11086
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7274 14596 7686
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14568 6662 14596 7210
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14292 5868 14504 5896
rect 14292 5001 14320 5868
rect 14568 5794 14596 6598
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15028 5846 15056 6258
rect 15120 6118 15148 7754
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15212 6934 15240 7346
rect 15290 7168 15346 7177
rect 15290 7103 15346 7112
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15016 5840 15068 5846
rect 14464 5772 14516 5778
rect 14568 5766 14688 5794
rect 15016 5782 15068 5788
rect 14464 5714 14516 5720
rect 14476 5234 14504 5714
rect 14660 5710 14688 5766
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14660 5370 14688 5646
rect 15014 5536 15070 5545
rect 15120 5522 15148 6054
rect 15070 5494 15148 5522
rect 15014 5471 15070 5480
rect 15028 5370 15056 5471
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14108 4950 14228 4978
rect 14278 4992 14334 5001
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 13820 4422 13872 4428
rect 13910 4448 13966 4457
rect 13832 3602 13860 4422
rect 13910 4383 13966 4392
rect 14016 3670 14044 4558
rect 14108 4554 14136 4950
rect 14278 4927 14334 4936
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 14016 3194 14044 3606
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14108 2922 14136 3334
rect 14200 2990 14228 4762
rect 14384 4706 14412 5034
rect 14476 4826 14504 5170
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15106 4856 15162 4865
rect 14464 4820 14516 4826
rect 15106 4791 15162 4800
rect 14464 4762 14516 4768
rect 14384 4678 14504 4706
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14188 2984 14240 2990
rect 14292 2961 14320 3538
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14384 3194 14412 3402
rect 14476 3369 14504 4678
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14660 4146 14688 4558
rect 15120 4486 15148 4791
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15304 4298 15332 7103
rect 15396 6254 15424 11154
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15672 9897 15700 10950
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15580 8634 15608 8910
rect 15672 8634 15700 9823
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15474 8528 15530 8537
rect 15474 8463 15530 8472
rect 15488 8294 15516 8463
rect 15476 8288 15528 8294
rect 15764 8242 15792 9590
rect 15948 9382 15976 9930
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15476 8230 15528 8236
rect 15672 8214 15792 8242
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15488 7478 15516 7958
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7721 15608 7754
rect 15566 7712 15622 7721
rect 15566 7647 15622 7656
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15580 6934 15608 7647
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 5001 15424 5510
rect 15382 4992 15438 5001
rect 15382 4927 15438 4936
rect 15396 4690 15424 4927
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15212 4270 15332 4298
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3516 14596 3878
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15106 3768 15162 3777
rect 15106 3703 15162 3712
rect 14648 3528 14700 3534
rect 14568 3488 14648 3516
rect 14648 3470 14700 3476
rect 14462 3360 14518 3369
rect 14462 3295 14518 3304
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14188 2926 14240 2932
rect 14278 2952 14334 2961
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 14096 2916 14148 2922
rect 14278 2887 14334 2896
rect 14096 2858 14148 2864
rect 13820 2644 13872 2650
rect 13740 2604 13820 2632
rect 13820 2586 13872 2592
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13924 2514 13952 2858
rect 14476 2514 14504 3295
rect 15120 3194 15148 3703
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14568 2990 14596 3130
rect 14556 2984 14608 2990
rect 14832 2984 14884 2990
rect 14556 2926 14608 2932
rect 14830 2952 14832 2961
rect 14884 2952 14886 2961
rect 14830 2887 14886 2896
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15212 2514 15240 4270
rect 15488 3913 15516 6734
rect 15672 5778 15700 8214
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15764 7886 15792 8026
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15856 7750 15884 7890
rect 15948 7750 15976 9318
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15750 6624 15806 6633
rect 15750 6559 15806 6568
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15580 4826 15608 5170
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15474 3904 15530 3913
rect 15474 3839 15530 3848
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15304 3602 15332 3674
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15488 2514 15516 3839
rect 15764 3346 15792 6559
rect 15856 6322 15884 7686
rect 16040 7410 16068 11018
rect 16224 10810 16252 11494
rect 16408 11150 16436 11562
rect 16500 11558 16528 12106
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 11354 16528 11494
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16592 10826 16620 11018
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16500 10798 16620 10826
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16120 8968 16172 8974
rect 16118 8936 16120 8945
rect 16172 8936 16174 8945
rect 16118 8871 16174 8880
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 16040 6798 16068 6870
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15948 5778 15976 6122
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16040 5166 16068 6734
rect 16224 5386 16252 9454
rect 16132 5358 16252 5386
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16040 5001 16068 5102
rect 16026 4992 16082 5001
rect 16026 4927 16082 4936
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15948 4214 15976 4626
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 16132 3618 16160 5358
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4282 16252 4966
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16040 3590 16160 3618
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15672 3318 15792 3346
rect 15672 3233 15700 3318
rect 15658 3224 15714 3233
rect 15658 3159 15714 3168
rect 15842 3224 15898 3233
rect 15842 3159 15898 3168
rect 15752 2984 15804 2990
rect 15856 2972 15884 3159
rect 15948 3058 15976 3402
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15804 2944 15884 2972
rect 15752 2926 15804 2932
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 15948 2825 15976 2858
rect 15934 2816 15990 2825
rect 15934 2751 15990 2760
rect 16040 2553 16068 3590
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16132 3233 16160 3470
rect 16118 3224 16174 3233
rect 16118 3159 16174 3168
rect 16026 2544 16082 2553
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15476 2508 15528 2514
rect 16026 2479 16082 2488
rect 15476 2450 15528 2456
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 12452 800 12480 2246
rect 12912 800 12940 2246
rect 13372 800 13400 2246
rect 13740 800 13768 2246
rect 14200 800 14228 2246
rect 14660 800 14688 2246
rect 15120 800 15148 2246
rect 15488 800 15516 2314
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 15948 800 15976 2246
rect 16316 1970 16344 9862
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 7546 16436 9318
rect 16500 8401 16528 10798
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9722 16620 9862
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16486 8392 16542 8401
rect 16486 8327 16542 8336
rect 16592 8022 16620 8774
rect 16684 8090 16712 10406
rect 16960 9654 16988 10406
rect 17328 10266 17356 13194
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 12102 17448 12582
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 18510 12336 18566 12345
rect 18510 12271 18566 12280
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 10810 17448 12038
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18524 11218 18552 12271
rect 19062 12200 19118 12209
rect 19062 12135 19064 12144
rect 19116 12135 19118 12144
rect 19064 12106 19116 12112
rect 19076 11694 19104 12106
rect 19614 11792 19670 11801
rect 19614 11727 19670 11736
rect 19628 11694 19656 11727
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17604 10674 17632 11154
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18524 10742 18552 11154
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17604 10198 17632 10610
rect 17972 10266 18000 10678
rect 18144 10600 18196 10606
rect 18142 10568 18144 10577
rect 18196 10568 18198 10577
rect 18142 10503 18198 10512
rect 18616 10266 18644 11018
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8430 16896 8978
rect 17144 8430 17172 9046
rect 16856 8424 16908 8430
rect 17132 8424 17184 8430
rect 16856 8366 16908 8372
rect 16946 8392 17002 8401
rect 17132 8366 17184 8372
rect 16946 8327 16948 8336
rect 17000 8327 17002 8336
rect 16948 8298 17000 8304
rect 16762 8120 16818 8129
rect 16672 8084 16724 8090
rect 16762 8055 16818 8064
rect 16672 8026 16724 8032
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16684 7954 16712 8026
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16408 6254 16436 7482
rect 16500 7206 16528 7482
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16670 6488 16726 6497
rect 16670 6423 16726 6432
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16500 6100 16528 6190
rect 16684 6118 16712 6423
rect 16672 6112 16724 6118
rect 16500 6072 16620 6100
rect 16592 5846 16620 6072
rect 16672 6054 16724 6060
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16500 5001 16528 5714
rect 16592 5030 16620 5782
rect 16580 5024 16632 5030
rect 16486 4992 16542 5001
rect 16580 4966 16632 4972
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16486 4927 16542 4936
rect 16684 4842 16712 4966
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16500 4814 16712 4842
rect 16408 4282 16436 4762
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16500 3618 16528 4814
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16592 4282 16620 4694
rect 16776 4321 16804 8055
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16868 6322 16896 6802
rect 16960 6633 16988 7822
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 16946 6624 17002 6633
rect 16946 6559 17002 6568
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16856 6180 16908 6186
rect 17052 6168 17080 7754
rect 17236 7002 17264 9318
rect 17880 9110 17908 10134
rect 17972 9722 18000 10202
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 18616 9586 18644 10202
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17314 8392 17370 8401
rect 17590 8392 17646 8401
rect 17370 8350 17540 8378
rect 17314 8327 17370 8336
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17328 8090 17356 8230
rect 17512 8090 17540 8350
rect 17788 8378 17816 8910
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 17866 8664 17922 8673
rect 18116 8656 18412 8676
rect 17866 8599 17922 8608
rect 17880 8498 17908 8599
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17590 8327 17646 8336
rect 17696 8350 17816 8378
rect 18052 8356 18104 8362
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17328 7002 17356 7346
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17328 6322 17356 6938
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17512 6322 17540 6598
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 16908 6140 17080 6168
rect 16856 6122 16908 6128
rect 16946 5944 17002 5953
rect 16946 5879 17002 5888
rect 16856 5092 16908 5098
rect 16856 5034 16908 5040
rect 16868 4554 16896 5034
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16762 4312 16818 4321
rect 16580 4276 16632 4282
rect 16762 4247 16818 4256
rect 16580 4218 16632 4224
rect 16868 4146 16896 4490
rect 16960 4486 16988 5879
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16672 4140 16724 4146
rect 16408 3602 16528 3618
rect 16396 3596 16528 3602
rect 16448 3590 16528 3596
rect 16592 4100 16672 4128
rect 16396 3538 16448 3544
rect 16592 3058 16620 4100
rect 16672 4082 16724 4088
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16670 4040 16726 4049
rect 16670 3975 16672 3984
rect 16724 3975 16726 3984
rect 16672 3946 16724 3952
rect 16670 3632 16726 3641
rect 16670 3567 16726 3576
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16684 2961 16712 3567
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 3058 16896 3470
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16960 2990 16988 4422
rect 17052 3602 17080 6140
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17512 5846 17540 6054
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17130 5672 17186 5681
rect 17130 5607 17186 5616
rect 17144 5302 17172 5607
rect 17420 5370 17448 5714
rect 17604 5409 17632 8327
rect 17696 6254 17724 8350
rect 18052 8298 18104 8304
rect 17776 7744 17828 7750
rect 18064 7732 18092 8298
rect 18328 8288 18380 8294
rect 18156 8265 18328 8276
rect 18142 8256 18328 8265
rect 18198 8248 18328 8256
rect 18328 8230 18380 8236
rect 18142 8191 18198 8200
rect 18524 7857 18552 8774
rect 18510 7848 18566 7857
rect 18510 7783 18566 7792
rect 17776 7686 17828 7692
rect 17972 7704 18092 7732
rect 17788 6361 17816 7686
rect 17972 7585 18000 7704
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 17958 7576 18014 7585
rect 18116 7568 18412 7588
rect 17958 7511 18014 7520
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17972 7177 18000 7346
rect 18236 7200 18288 7206
rect 17958 7168 18014 7177
rect 18236 7142 18288 7148
rect 17958 7103 18014 7112
rect 18248 7002 18276 7142
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 17774 6352 17830 6361
rect 17774 6287 17830 6296
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17684 6112 17736 6118
rect 17682 6080 17684 6089
rect 17776 6112 17828 6118
rect 17736 6080 17738 6089
rect 17776 6054 17828 6060
rect 17682 6015 17738 6024
rect 17788 5846 17816 6054
rect 17776 5840 17828 5846
rect 17774 5808 17776 5817
rect 17828 5808 17830 5817
rect 17684 5772 17736 5778
rect 17774 5743 17830 5752
rect 17684 5714 17736 5720
rect 17590 5400 17646 5409
rect 17408 5364 17460 5370
rect 17590 5335 17646 5344
rect 17408 5306 17460 5312
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17144 3738 17172 4694
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17236 3942 17264 4422
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17328 3738 17356 4626
rect 17420 4622 17448 5306
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 16948 2984 17000 2990
rect 16670 2952 16726 2961
rect 16948 2926 17000 2932
rect 16670 2887 16726 2896
rect 16684 2514 16712 2887
rect 17144 2514 17172 3674
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17236 3369 17264 3538
rect 17222 3360 17278 3369
rect 17222 3295 17278 3304
rect 17604 2938 17632 4082
rect 17696 3194 17724 5714
rect 17880 5642 17908 6938
rect 18616 6905 18644 8842
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18708 8362 18736 8774
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18708 7528 18736 8026
rect 18800 7993 18828 8774
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18786 7984 18842 7993
rect 18786 7919 18842 7928
rect 18788 7540 18840 7546
rect 18708 7500 18788 7528
rect 18788 7482 18840 7488
rect 17958 6896 18014 6905
rect 17958 6831 18014 6840
rect 18602 6896 18658 6905
rect 18602 6831 18658 6840
rect 18696 6860 18748 6866
rect 17972 6225 18000 6831
rect 18696 6802 18748 6808
rect 18420 6792 18472 6798
rect 18418 6760 18420 6769
rect 18472 6760 18474 6769
rect 18418 6695 18474 6704
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17958 6216 18014 6225
rect 17958 6151 18014 6160
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 18064 5953 18092 6122
rect 18050 5944 18106 5953
rect 18050 5879 18106 5888
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 17788 4214 17816 4966
rect 18052 4820 18104 4826
rect 18144 4820 18196 4826
rect 18104 4780 18144 4808
rect 18052 4762 18104 4768
rect 18144 4762 18196 4768
rect 18432 4706 18460 4966
rect 18524 4826 18552 6666
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18616 6322 18644 6598
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18708 5846 18736 6802
rect 18800 6361 18828 7482
rect 18892 6866 18920 8366
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18892 6497 18920 6802
rect 18878 6488 18934 6497
rect 18878 6423 18934 6432
rect 18786 6352 18842 6361
rect 18786 6287 18842 6296
rect 18880 6248 18932 6254
rect 18800 6208 18880 6236
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18616 4865 18644 5510
rect 18708 5370 18736 5782
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18694 4992 18750 5001
rect 18694 4927 18750 4936
rect 18602 4856 18658 4865
rect 18512 4820 18564 4826
rect 18708 4826 18736 4927
rect 18602 4791 18658 4800
rect 18696 4820 18748 4826
rect 18512 4762 18564 4768
rect 18696 4762 18748 4768
rect 18432 4678 18644 4706
rect 18432 4554 18460 4678
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17788 3738 17816 4150
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 18236 3936 18288 3942
rect 18328 3936 18380 3942
rect 18236 3878 18288 3884
rect 18326 3904 18328 3913
rect 18380 3904 18382 3913
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17328 2922 17632 2938
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 17316 2916 17632 2922
rect 17368 2910 17632 2916
rect 17316 2858 17368 2864
rect 17604 2514 17632 2910
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16408 800 16436 2314
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 800 16896 2246
rect 17420 1170 17448 2314
rect 17328 1142 17448 1170
rect 17328 800 17356 1142
rect 17696 800 17724 2790
rect 17788 2514 17816 2926
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17880 2038 17908 3878
rect 18248 3670 18276 3878
rect 18326 3839 18382 3848
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18432 3466 18460 3946
rect 18616 3738 18644 4678
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18708 3670 18736 4626
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 2446 18000 3334
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18602 3224 18658 3233
rect 18602 3159 18658 3168
rect 18616 2990 18644 3159
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 17960 2440 18012 2446
rect 18156 2417 18184 2858
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 17960 2382 18012 2388
rect 18142 2408 18198 2417
rect 18142 2343 18198 2352
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17868 2032 17920 2038
rect 17868 1974 17920 1980
rect 18144 1420 18196 1426
rect 18144 1362 18196 1368
rect 18156 800 18184 1362
rect 18616 800 18644 2790
rect 18800 2514 18828 6208
rect 18880 6190 18932 6196
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 2825 18920 5646
rect 18878 2816 18934 2825
rect 18878 2751 18934 2760
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 18984 898 19012 10406
rect 19076 3738 19104 11018
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19168 9178 19196 9658
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19168 8566 19196 9114
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19168 6798 19196 7278
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19168 6458 19196 6598
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19154 6352 19210 6361
rect 19154 6287 19210 6296
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19168 2514 19196 6287
rect 19260 4078 19288 11494
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10742 19472 11086
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19444 10266 19472 10678
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20088 8838 20116 9318
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 7041 19380 8298
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 19338 7032 19394 7041
rect 19338 6967 19394 6976
rect 19340 6792 19392 6798
rect 19536 6769 19564 7686
rect 19812 7449 19840 7686
rect 19798 7440 19854 7449
rect 19798 7375 19854 7384
rect 20180 7313 20208 7686
rect 20166 7304 20222 7313
rect 20166 7239 20222 7248
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19340 6734 19392 6740
rect 19522 6760 19578 6769
rect 19352 6458 19380 6734
rect 19522 6695 19578 6704
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19430 5808 19486 5817
rect 19536 5778 19564 6598
rect 19430 5743 19486 5752
rect 19524 5772 19576 5778
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19352 5370 19380 5578
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19352 3641 19380 4966
rect 19444 4758 19472 5743
rect 19524 5714 19576 5720
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19444 4282 19472 4694
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19536 3777 19564 5510
rect 19522 3768 19578 3777
rect 19432 3732 19484 3738
rect 19522 3703 19578 3712
rect 19432 3674 19484 3680
rect 19338 3632 19394 3641
rect 19338 3567 19394 3576
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19260 2582 19288 3334
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19076 1426 19104 2246
rect 19064 1420 19116 1426
rect 19064 1362 19116 1368
rect 18984 870 19104 898
rect 19076 800 19104 870
rect 19444 800 19472 3674
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19628 1834 19656 3334
rect 19720 3097 19748 7142
rect 19892 5568 19944 5574
rect 19812 5528 19892 5556
rect 19706 3088 19762 3097
rect 19706 3023 19762 3032
rect 19812 2990 19840 5528
rect 19892 5510 19944 5516
rect 20088 4185 20116 7142
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20180 5273 20208 6598
rect 20166 5264 20222 5273
rect 20166 5199 20222 5208
rect 20074 4176 20130 4185
rect 20074 4111 20130 4120
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19616 1828 19668 1834
rect 19616 1770 19668 1776
rect 19904 800 19932 4014
rect 19982 3496 20038 3505
rect 19982 3431 19984 3440
rect 20036 3431 20038 3440
rect 19984 3402 20036 3408
rect 19996 2990 20024 3402
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 20088 2514 20116 2994
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20180 2106 20208 2382
rect 20168 2100 20220 2106
rect 20168 2042 20220 2048
rect 20364 800 20392 11494
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20456 9722 20484 10202
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20824 9654 20852 12378
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20732 8634 20760 9046
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21192 8634 21220 8774
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 20732 8090 20760 8570
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20548 4826 20576 5170
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20824 4593 20852 6734
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21270 6080 21326 6089
rect 21192 4729 21220 6054
rect 21270 6015 21326 6024
rect 21178 4720 21234 4729
rect 21178 4655 21234 4664
rect 20810 4584 20866 4593
rect 20810 4519 20866 4528
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 20824 800 20852 3062
rect 20916 2650 20944 3878
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21284 898 21312 6015
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21192 870 21312 898
rect 21192 800 21220 870
rect 21652 800 21680 2790
rect 22112 800 22140 2858
rect 22572 800 22600 2994
rect 2226 640 2282 649
rect 2226 575 2282 584
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10690 0 10746 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14186 0 14242 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19890 0 19946 800
rect 20350 0 20406 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
<< via2 >>
rect 4066 22480 4122 22536
rect 3146 22072 3202 22128
rect 2778 21120 2834 21176
rect 2870 20576 2926 20632
rect 1950 19760 2006 19816
rect 2962 20168 3018 20224
rect 2778 19216 2834 19272
rect 2318 19080 2374 19136
rect 1950 18808 2006 18864
rect 1858 18264 1914 18320
rect 1950 17876 2006 17912
rect 1950 17856 1952 17876
rect 1952 17856 2004 17876
rect 2004 17856 2006 17876
rect 1950 16904 2006 16960
rect 1766 16496 1822 16552
rect 1674 15952 1730 16008
rect 1674 15544 1730 15600
rect 1582 13232 1638 13288
rect 1858 14612 1914 14648
rect 1858 14592 1860 14612
rect 1860 14592 1912 14612
rect 1912 14592 1914 14612
rect 3238 21528 3294 21584
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 3330 19080 3386 19136
rect 1950 14068 2006 14104
rect 1950 14048 1952 14068
rect 1952 14048 2004 14068
rect 2004 14048 2006 14068
rect 2410 12824 2466 12880
rect 2318 11600 2374 11656
rect 1214 1944 1270 2000
rect 1306 992 1362 1048
rect 2502 11192 2558 11248
rect 3238 17312 3294 17368
rect 3146 16904 3202 16960
rect 3146 15000 3202 15056
rect 3790 17040 3846 17096
rect 2778 13640 2834 13696
rect 2318 9288 2374 9344
rect 2134 9016 2190 9072
rect 2042 2896 2098 2952
rect 2410 9152 2466 9208
rect 2686 9560 2742 9616
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 2962 12280 3018 12336
rect 2962 11736 3018 11792
rect 2870 9424 2926 9480
rect 2502 7792 2558 7848
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3698 12688 3754 12744
rect 3698 11736 3754 11792
rect 3698 10784 3754 10840
rect 3514 9424 3570 9480
rect 3422 8200 3478 8256
rect 3146 7248 3202 7304
rect 3422 7248 3478 7304
rect 2226 4820 2282 4856
rect 2226 4800 2228 4820
rect 2228 4800 2280 4820
rect 2280 4800 2282 4820
rect 2134 2760 2190 2816
rect 1582 176 1638 232
rect 2410 2488 2466 2544
rect 3606 5888 3662 5944
rect 3146 5072 3202 5128
rect 2778 4548 2834 4584
rect 2778 4528 2780 4548
rect 2780 4528 2832 4548
rect 2832 4528 2834 4548
rect 2778 3984 2834 4040
rect 2778 2624 2834 2680
rect 2594 1536 2650 1592
rect 3238 4528 3294 4584
rect 3054 3440 3110 3496
rect 3514 4120 3570 4176
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4986 12960 5042 13016
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 10104 4122 10160
rect 3974 9968 4030 10024
rect 3974 8880 4030 8936
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4802 11328 4858 11384
rect 4802 10512 4858 10568
rect 4802 10376 4858 10432
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4802 9968 4858 10024
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 5446 12724 5448 12744
rect 5448 12724 5500 12744
rect 5500 12724 5502 12744
rect 5446 12688 5502 12724
rect 5170 9832 5226 9888
rect 5262 9560 5318 9616
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4066 7520 4122 7576
rect 3974 7112 4030 7168
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 4066 6704 4122 6760
rect 4894 7928 4950 7984
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4802 7656 4858 7712
rect 4710 7384 4766 7440
rect 4434 6976 4490 7032
rect 4710 6740 4712 6760
rect 4712 6740 4764 6760
rect 4764 6740 4766 6760
rect 4710 6704 4766 6740
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 3882 6160 3938 6216
rect 4066 5752 4122 5808
rect 3974 5616 4030 5672
rect 4066 5208 4122 5264
rect 4066 4256 4122 4312
rect 4066 4120 4122 4176
rect 3882 3576 3938 3632
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4894 3712 4950 3768
rect 4526 3576 4582 3632
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4710 3032 4766 3088
rect 4618 2932 4620 2952
rect 4620 2932 4672 2952
rect 4672 2932 4674 2952
rect 4618 2896 4674 2932
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5354 4392 5410 4448
rect 5262 3340 5264 3360
rect 5264 3340 5316 3360
rect 5316 3340 5318 3360
rect 5262 3304 5318 3340
rect 5630 7520 5686 7576
rect 5906 12588 5908 12608
rect 5908 12588 5960 12608
rect 5960 12588 5962 12608
rect 5906 12552 5962 12588
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 6458 12552 6514 12608
rect 5998 8880 6054 8936
rect 5630 5772 5686 5808
rect 5630 5752 5632 5772
rect 5632 5752 5684 5772
rect 5684 5752 5686 5772
rect 5814 4120 5870 4176
rect 6182 8608 6238 8664
rect 6182 7520 6238 7576
rect 6182 6840 6238 6896
rect 6366 9560 6422 9616
rect 7102 12688 7158 12744
rect 7286 12008 7342 12064
rect 7010 11464 7066 11520
rect 6826 11056 6882 11112
rect 6734 9152 6790 9208
rect 6550 9036 6606 9072
rect 6550 9016 6552 9036
rect 6552 9016 6604 9036
rect 6604 9016 6606 9036
rect 6366 6840 6422 6896
rect 6826 8064 6882 8120
rect 6642 5888 6698 5944
rect 6458 5480 6514 5536
rect 6366 4664 6422 4720
rect 6642 5616 6698 5672
rect 6918 7656 6974 7712
rect 7378 9288 7434 9344
rect 7102 7792 7158 7848
rect 7286 7792 7342 7848
rect 7102 7248 7158 7304
rect 6826 6160 6882 6216
rect 6826 5208 6882 5264
rect 7194 5752 7250 5808
rect 7102 3712 7158 3768
rect 6918 2624 6974 2680
rect 7286 2896 7342 2952
rect 7378 2488 7434 2544
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 8114 12960 8170 13016
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7930 11636 7932 11656
rect 7932 11636 7984 11656
rect 7984 11636 7986 11656
rect 7930 11600 7986 11636
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8298 11600 8354 11656
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7838 9868 7840 9888
rect 7840 9868 7892 9888
rect 7892 9868 7894 9888
rect 7838 9832 7894 9868
rect 7838 9580 7894 9616
rect 7838 9560 7840 9580
rect 7840 9560 7892 9580
rect 7892 9560 7894 9580
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 8666 12416 8722 12472
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 9770 13676 9772 13696
rect 9772 13676 9824 13696
rect 9824 13676 9826 13696
rect 9770 13640 9826 13676
rect 9678 13504 9734 13560
rect 9770 13368 9826 13424
rect 9126 12688 9182 12744
rect 8574 10376 8630 10432
rect 8574 8372 8576 8392
rect 8576 8372 8628 8392
rect 8628 8372 8630 8392
rect 8574 8336 8630 8372
rect 8298 7928 8354 7984
rect 8022 7692 8024 7712
rect 8024 7692 8076 7712
rect 8076 7692 8078 7712
rect 8022 7656 8078 7692
rect 8298 7112 8354 7168
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8298 5752 8354 5808
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7746 4392 7802 4448
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8390 3304 8446 3360
rect 9034 9988 9090 10024
rect 9034 9968 9036 9988
rect 9036 9968 9088 9988
rect 9088 9968 9090 9988
rect 9034 8744 9090 8800
rect 8850 8336 8906 8392
rect 10598 14320 10654 14376
rect 10322 13912 10378 13968
rect 9954 13368 10010 13424
rect 9678 11464 9734 11520
rect 9402 8608 9458 8664
rect 8574 5616 8630 5672
rect 8574 4428 8576 4448
rect 8576 4428 8628 4448
rect 8628 4428 8630 4448
rect 8574 4392 8630 4428
rect 9770 8880 9826 8936
rect 10046 11328 10102 11384
rect 9954 8880 10010 8936
rect 9954 8608 10010 8664
rect 9770 6024 9826 6080
rect 9678 5888 9734 5944
rect 8666 3168 8722 3224
rect 8574 2760 8630 2816
rect 9586 4664 9642 4720
rect 9586 4256 9642 4312
rect 10506 10648 10562 10704
rect 10598 10376 10654 10432
rect 9954 5092 10010 5128
rect 9954 5072 9956 5092
rect 9956 5072 10008 5092
rect 10008 5072 10010 5092
rect 10414 3168 10470 3224
rect 10598 3848 10654 3904
rect 10598 2352 10654 2408
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 10874 12844 10930 12880
rect 10874 12824 10876 12844
rect 10876 12824 10928 12844
rect 10928 12824 10930 12844
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 10782 12008 10838 12064
rect 11058 12436 11114 12472
rect 11058 12416 11060 12436
rect 11060 12416 11112 12436
rect 11112 12416 11114 12436
rect 11610 12416 11666 12472
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11242 11056 11298 11112
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 10782 8880 10838 8936
rect 10874 8608 10930 8664
rect 10782 8472 10838 8528
rect 10966 8336 11022 8392
rect 11334 10104 11390 10160
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11150 9288 11206 9344
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11794 9868 11796 9888
rect 11796 9868 11848 9888
rect 11848 9868 11850 9888
rect 11794 9832 11850 9868
rect 11702 9560 11758 9616
rect 10874 7928 10930 7984
rect 10874 7520 10930 7576
rect 10782 5752 10838 5808
rect 11610 7792 11666 7848
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11886 8200 11942 8256
rect 11610 7112 11666 7168
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11150 6024 11206 6080
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 10966 4392 11022 4448
rect 11058 3168 11114 3224
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 10874 2796 10876 2816
rect 10876 2796 10928 2816
rect 10928 2796 10930 2816
rect 10874 2760 10930 2796
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 11886 7520 11942 7576
rect 11794 6432 11850 6488
rect 11886 6296 11942 6352
rect 12070 11500 12072 11520
rect 12072 11500 12124 11520
rect 12124 11500 12126 11520
rect 12070 11464 12126 11500
rect 12070 10412 12072 10432
rect 12072 10412 12124 10432
rect 12124 10412 12126 10432
rect 12070 10376 12126 10412
rect 12438 13912 12494 13968
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 17212 17960 17232
rect 17960 17212 18012 17232
rect 18012 17212 18014 17232
rect 17958 17176 18014 17212
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 13358 14320 13414 14376
rect 12530 13640 12586 13696
rect 12898 13524 12954 13560
rect 12898 13504 12900 13524
rect 12900 13504 12952 13524
rect 12952 13504 12954 13524
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 12714 12436 12770 12472
rect 12714 12416 12716 12436
rect 12716 12416 12768 12436
rect 12768 12416 12770 12436
rect 12162 10240 12218 10296
rect 12346 11464 12402 11520
rect 12530 11464 12586 11520
rect 12162 5616 12218 5672
rect 12070 5072 12126 5128
rect 11978 4392 12034 4448
rect 11886 3848 11942 3904
rect 12622 6840 12678 6896
rect 12530 6296 12586 6352
rect 12622 5616 12678 5672
rect 12806 5752 12862 5808
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 13726 11636 13728 11656
rect 13728 11636 13780 11656
rect 13780 11636 13782 11656
rect 13726 11600 13782 11636
rect 13174 9288 13230 9344
rect 12438 4800 12494 4856
rect 13634 11192 13690 11248
rect 13818 10648 13874 10704
rect 13450 9424 13506 9480
rect 13450 9288 13506 9344
rect 13634 9968 13690 10024
rect 13450 6568 13506 6624
rect 13450 6296 13506 6352
rect 13818 9288 13874 9344
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14278 11328 14334 11384
rect 14186 9968 14242 10024
rect 14278 9560 14334 9616
rect 14186 8492 14242 8528
rect 14186 8472 14188 8492
rect 14188 8472 14240 8492
rect 14240 8472 14242 8492
rect 14186 8064 14242 8120
rect 14186 7656 14242 7712
rect 14278 7248 14334 7304
rect 13726 5888 13782 5944
rect 13542 5616 13598 5672
rect 13542 4800 13598 4856
rect 13542 4120 13598 4176
rect 13542 3576 13598 3632
rect 13542 3032 13598 3088
rect 13818 5208 13874 5264
rect 14278 6976 14334 7032
rect 14094 6860 14150 6896
rect 14094 6840 14096 6860
rect 14096 6840 14148 6860
rect 14148 6840 14150 6860
rect 14278 6568 14334 6624
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14646 9460 14648 9480
rect 14648 9460 14700 9480
rect 14700 9460 14702 9480
rect 14646 9424 14702 9460
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 15198 9016 15254 9072
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 15290 7112 15346 7168
rect 15014 5480 15070 5536
rect 13910 4392 13966 4448
rect 14278 4936 14334 4992
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 15106 4800 15162 4856
rect 15658 9832 15714 9888
rect 15474 8472 15530 8528
rect 15566 7656 15622 7712
rect 15382 4936 15438 4992
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 15106 3712 15162 3768
rect 14462 3304 14518 3360
rect 14278 2896 14334 2952
rect 14830 2932 14832 2952
rect 14832 2932 14884 2952
rect 14884 2932 14886 2952
rect 14830 2896 14886 2932
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15750 6568 15806 6624
rect 15474 3848 15530 3904
rect 16118 8916 16120 8936
rect 16120 8916 16172 8936
rect 16172 8916 16174 8936
rect 16118 8880 16174 8916
rect 16026 4936 16082 4992
rect 15658 3168 15714 3224
rect 15842 3168 15898 3224
rect 15934 2760 15990 2816
rect 16118 3168 16174 3224
rect 16026 2488 16082 2544
rect 16486 8336 16542 8392
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18510 12280 18566 12336
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 19062 12164 19118 12200
rect 19062 12144 19064 12164
rect 19064 12144 19116 12164
rect 19116 12144 19118 12164
rect 19614 11736 19670 11792
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18142 10548 18144 10568
rect 18144 10548 18196 10568
rect 18196 10548 18198 10568
rect 18142 10512 18198 10548
rect 16946 8356 17002 8392
rect 16946 8336 16948 8356
rect 16948 8336 17000 8356
rect 17000 8336 17002 8356
rect 16762 8064 16818 8120
rect 16670 6432 16726 6488
rect 16486 4936 16542 4992
rect 16946 6568 17002 6624
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17314 8336 17370 8392
rect 17590 8336 17646 8392
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 17866 8608 17922 8664
rect 16946 5888 17002 5944
rect 16762 4256 16818 4312
rect 16670 4004 16726 4040
rect 16670 3984 16672 4004
rect 16672 3984 16724 4004
rect 16724 3984 16726 4004
rect 16670 3576 16726 3632
rect 17130 5616 17186 5672
rect 18142 8200 18198 8256
rect 18510 7792 18566 7848
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 17958 7520 18014 7576
rect 17958 7112 18014 7168
rect 17774 6296 17830 6352
rect 17682 6060 17684 6080
rect 17684 6060 17736 6080
rect 17736 6060 17738 6080
rect 17682 6024 17738 6060
rect 17774 5788 17776 5808
rect 17776 5788 17828 5808
rect 17828 5788 17830 5808
rect 17774 5752 17830 5788
rect 17590 5344 17646 5400
rect 16670 2896 16726 2952
rect 17222 3304 17278 3360
rect 18786 7928 18842 7984
rect 17958 6840 18014 6896
rect 18602 6840 18658 6896
rect 18418 6740 18420 6760
rect 18420 6740 18472 6760
rect 18472 6740 18474 6760
rect 18418 6704 18474 6740
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17958 6160 18014 6216
rect 18050 5888 18106 5944
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18878 6432 18934 6488
rect 18786 6296 18842 6352
rect 18694 4936 18750 4992
rect 18602 4800 18658 4856
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18326 3884 18328 3904
rect 18328 3884 18380 3904
rect 18380 3884 18382 3904
rect 18326 3848 18382 3884
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18602 3168 18658 3224
rect 18142 2352 18198 2408
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18878 2760 18934 2816
rect 19154 6296 19210 6352
rect 19338 6976 19394 7032
rect 19798 7384 19854 7440
rect 20166 7248 20222 7304
rect 19522 6704 19578 6760
rect 19430 5752 19486 5808
rect 19522 3712 19578 3768
rect 19338 3576 19394 3632
rect 19706 3032 19762 3088
rect 20166 5208 20222 5264
rect 20074 4120 20130 4176
rect 19982 3460 20038 3496
rect 19982 3440 19984 3460
rect 19984 3440 20036 3460
rect 20036 3440 20038 3460
rect 21270 6024 21326 6080
rect 21178 4664 21234 4720
rect 20810 4528 20866 4584
rect 2226 584 2282 640
<< metal3 >>
rect 0 22538 800 22568
rect 4061 22538 4127 22541
rect 0 22536 4127 22538
rect 0 22480 4066 22536
rect 4122 22480 4127 22536
rect 0 22478 4127 22480
rect 0 22448 800 22478
rect 4061 22475 4127 22478
rect 0 22130 800 22160
rect 3141 22130 3207 22133
rect 0 22128 3207 22130
rect 0 22072 3146 22128
rect 3202 22072 3207 22128
rect 0 22070 3207 22072
rect 0 22040 800 22070
rect 3141 22067 3207 22070
rect 0 21586 800 21616
rect 3233 21586 3299 21589
rect 0 21584 3299 21586
rect 0 21528 3238 21584
rect 3294 21528 3299 21584
rect 0 21526 3299 21528
rect 0 21496 800 21526
rect 3233 21523 3299 21526
rect 0 21178 800 21208
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 0 20634 800 20664
rect 2865 20634 2931 20637
rect 0 20632 2931 20634
rect 0 20576 2870 20632
rect 2926 20576 2931 20632
rect 0 20574 2931 20576
rect 0 20544 800 20574
rect 2865 20571 2931 20574
rect 0 20226 800 20256
rect 2957 20226 3023 20229
rect 0 20224 3023 20226
rect 0 20168 2962 20224
rect 3018 20168 3023 20224
rect 0 20166 3023 20168
rect 0 20136 800 20166
rect 2957 20163 3023 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 800 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 800 19758
rect 1945 19755 2011 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 800 19304
rect 2773 19274 2839 19277
rect 0 19272 2839 19274
rect 0 19216 2778 19272
rect 2834 19216 2839 19272
rect 0 19214 2839 19216
rect 0 19184 800 19214
rect 2773 19211 2839 19214
rect 2313 19138 2379 19141
rect 3325 19138 3391 19141
rect 2313 19136 3391 19138
rect 2313 19080 2318 19136
rect 2374 19080 3330 19136
rect 3386 19080 3391 19136
rect 2313 19078 3391 19080
rect 2313 19075 2379 19078
rect 3325 19075 3391 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 800 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 800 18806
rect 1945 18803 2011 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 800 18352
rect 1853 18322 1919 18325
rect 0 18320 1919 18322
rect 0 18264 1858 18320
rect 1914 18264 1919 18320
rect 0 18262 1919 18264
rect 0 18232 800 18262
rect 1853 18259 1919 18262
rect 7808 17984 8128 17985
rect 0 17914 800 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 800 17854
rect 1945 17851 2011 17854
rect 4376 17440 4696 17441
rect 0 17370 800 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 3233 17370 3299 17373
rect 0 17368 3299 17370
rect 0 17312 3238 17368
rect 3294 17312 3299 17368
rect 0 17310 3299 17312
rect 0 17280 800 17310
rect 3233 17307 3299 17310
rect 17953 17234 18019 17237
rect 22000 17234 22800 17264
rect 17953 17232 22800 17234
rect 17953 17176 17958 17232
rect 18014 17176 22800 17232
rect 17953 17174 22800 17176
rect 17953 17171 18019 17174
rect 22000 17144 22800 17174
rect 3785 17098 3851 17101
rect 3742 17096 3851 17098
rect 3742 17040 3790 17096
rect 3846 17040 3851 17096
rect 3742 17035 3851 17040
rect 0 16962 800 16992
rect 1945 16962 2011 16965
rect 0 16960 2011 16962
rect 0 16904 1950 16960
rect 2006 16904 2011 16960
rect 0 16902 2011 16904
rect 0 16872 800 16902
rect 1945 16899 2011 16902
rect 3141 16962 3207 16965
rect 3742 16962 3802 17035
rect 3141 16960 3802 16962
rect 3141 16904 3146 16960
rect 3202 16904 3802 16960
rect 3141 16902 3802 16904
rect 3141 16899 3207 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 0 16554 800 16584
rect 1761 16554 1827 16557
rect 0 16552 1827 16554
rect 0 16496 1766 16552
rect 1822 16496 1827 16552
rect 0 16494 1827 16496
rect 0 16464 800 16494
rect 1761 16491 1827 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 800 16040
rect 1669 16010 1735 16013
rect 0 16008 1735 16010
rect 0 15952 1674 16008
rect 1730 15952 1735 16008
rect 0 15950 1735 15952
rect 0 15920 800 15950
rect 1669 15947 1735 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 800 15632
rect 1669 15602 1735 15605
rect 0 15600 1735 15602
rect 0 15544 1674 15600
rect 1730 15544 1735 15600
rect 0 15542 1735 15544
rect 0 15512 800 15542
rect 1669 15539 1735 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 800 15088
rect 3141 15058 3207 15061
rect 0 15056 3207 15058
rect 0 15000 3146 15056
rect 3202 15000 3207 15056
rect 0 14998 3207 15000
rect 0 14968 800 14998
rect 3141 14995 3207 14998
rect 7808 14720 8128 14721
rect 0 14650 800 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 800 14590
rect 1853 14587 1919 14590
rect 10593 14378 10659 14381
rect 13353 14378 13419 14381
rect 10593 14376 13419 14378
rect 10593 14320 10598 14376
rect 10654 14320 13358 14376
rect 13414 14320 13419 14376
rect 10593 14318 13419 14320
rect 10593 14315 10659 14318
rect 13353 14315 13419 14318
rect 4376 14176 4696 14177
rect 0 14106 800 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1945 14106 2011 14109
rect 0 14104 2011 14106
rect 0 14048 1950 14104
rect 2006 14048 2011 14104
rect 0 14046 2011 14048
rect 0 14016 800 14046
rect 1945 14043 2011 14046
rect 10317 13970 10383 13973
rect 12433 13970 12499 13973
rect 10317 13968 12499 13970
rect 10317 13912 10322 13968
rect 10378 13912 12438 13968
rect 12494 13912 12499 13968
rect 10317 13910 12499 13912
rect 10317 13907 10383 13910
rect 12433 13907 12499 13910
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 9765 13698 9831 13701
rect 12525 13698 12591 13701
rect 9765 13696 12591 13698
rect 9765 13640 9770 13696
rect 9826 13640 12530 13696
rect 12586 13640 12591 13696
rect 9765 13638 12591 13640
rect 9765 13635 9831 13638
rect 12525 13635 12591 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 9673 13562 9739 13565
rect 12893 13562 12959 13565
rect 9673 13560 12959 13562
rect 9673 13504 9678 13560
rect 9734 13504 12898 13560
rect 12954 13504 12959 13560
rect 9673 13502 12959 13504
rect 9673 13499 9739 13502
rect 12893 13499 12959 13502
rect 9765 13426 9831 13429
rect 9949 13426 10015 13429
rect 9765 13424 10015 13426
rect 9765 13368 9770 13424
rect 9826 13368 9954 13424
rect 10010 13368 10015 13424
rect 9765 13366 10015 13368
rect 9765 13363 9831 13366
rect 9949 13363 10015 13366
rect 0 13290 800 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 800 13230
rect 1577 13227 1643 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 4981 13018 5047 13021
rect 8109 13018 8175 13021
rect 4981 13016 8175 13018
rect 4981 12960 4986 13016
rect 5042 12960 8114 13016
rect 8170 12960 8175 13016
rect 4981 12958 8175 12960
rect 4981 12955 5047 12958
rect 8109 12955 8175 12958
rect 2405 12882 2471 12885
rect 10869 12882 10935 12885
rect 2405 12880 10935 12882
rect 2405 12824 2410 12880
rect 2466 12824 10874 12880
rect 10930 12824 10935 12880
rect 2405 12822 10935 12824
rect 2405 12819 2471 12822
rect 10869 12819 10935 12822
rect 0 12746 800 12776
rect 3693 12746 3759 12749
rect 0 12744 3759 12746
rect 0 12688 3698 12744
rect 3754 12688 3759 12744
rect 0 12686 3759 12688
rect 0 12656 800 12686
rect 3693 12683 3759 12686
rect 5441 12746 5507 12749
rect 7097 12746 7163 12749
rect 9121 12746 9187 12749
rect 5441 12744 7163 12746
rect 5441 12688 5446 12744
rect 5502 12688 7102 12744
rect 7158 12688 7163 12744
rect 5441 12686 7163 12688
rect 5441 12683 5507 12686
rect 7097 12683 7163 12686
rect 7238 12744 9187 12746
rect 7238 12688 9126 12744
rect 9182 12688 9187 12744
rect 7238 12686 9187 12688
rect 5901 12610 5967 12613
rect 6453 12610 6519 12613
rect 7238 12610 7298 12686
rect 9121 12683 9187 12686
rect 5901 12608 7298 12610
rect 5901 12552 5906 12608
rect 5962 12552 6458 12608
rect 6514 12552 7298 12608
rect 5901 12550 7298 12552
rect 5901 12547 5967 12550
rect 6453 12547 6519 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 8661 12474 8727 12477
rect 11053 12474 11119 12477
rect 8661 12472 11119 12474
rect 8661 12416 8666 12472
rect 8722 12416 11058 12472
rect 11114 12416 11119 12472
rect 8661 12414 11119 12416
rect 8661 12411 8727 12414
rect 11053 12411 11119 12414
rect 11605 12474 11671 12477
rect 12709 12474 12775 12477
rect 11605 12472 12775 12474
rect 11605 12416 11610 12472
rect 11666 12416 12714 12472
rect 12770 12416 12775 12472
rect 11605 12414 12775 12416
rect 11605 12411 11671 12414
rect 12709 12411 12775 12414
rect 0 12338 800 12368
rect 2957 12338 3023 12341
rect 18505 12338 18571 12341
rect 0 12278 2882 12338
rect 0 12248 800 12278
rect 2822 12202 2882 12278
rect 2957 12336 18571 12338
rect 2957 12280 2962 12336
rect 3018 12280 18510 12336
rect 18566 12280 18571 12336
rect 2957 12278 18571 12280
rect 2957 12275 3023 12278
rect 18505 12275 18571 12278
rect 19057 12202 19123 12205
rect 2822 12200 19123 12202
rect 2822 12144 19062 12200
rect 19118 12144 19123 12200
rect 2822 12142 19123 12144
rect 19057 12139 19123 12142
rect 7281 12066 7347 12069
rect 10777 12066 10843 12069
rect 7281 12064 10843 12066
rect 7281 12008 7286 12064
rect 7342 12008 10782 12064
rect 10838 12008 10843 12064
rect 7281 12006 10843 12008
rect 7281 12003 7347 12006
rect 10777 12003 10843 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 800 11824
rect 2957 11794 3023 11797
rect 0 11792 3023 11794
rect 0 11736 2962 11792
rect 3018 11736 3023 11792
rect 0 11734 3023 11736
rect 0 11704 800 11734
rect 2957 11731 3023 11734
rect 3693 11794 3759 11797
rect 19609 11794 19675 11797
rect 3693 11792 19675 11794
rect 3693 11736 3698 11792
rect 3754 11736 19614 11792
rect 19670 11736 19675 11792
rect 3693 11734 19675 11736
rect 3693 11731 3759 11734
rect 19609 11731 19675 11734
rect 2313 11658 2379 11661
rect 7925 11658 7991 11661
rect 2313 11656 7991 11658
rect 2313 11600 2318 11656
rect 2374 11600 7930 11656
rect 7986 11600 7991 11656
rect 2313 11598 7991 11600
rect 2313 11595 2379 11598
rect 7925 11595 7991 11598
rect 8293 11658 8359 11661
rect 13721 11658 13787 11661
rect 8293 11656 13787 11658
rect 8293 11600 8298 11656
rect 8354 11600 13726 11656
rect 13782 11600 13787 11656
rect 8293 11598 13787 11600
rect 8293 11595 8359 11598
rect 13721 11595 13787 11598
rect 7005 11522 7071 11525
rect 7230 11522 7236 11524
rect 7005 11520 7236 11522
rect 7005 11464 7010 11520
rect 7066 11464 7236 11520
rect 7005 11462 7236 11464
rect 7005 11459 7071 11462
rect 7230 11460 7236 11462
rect 7300 11460 7306 11524
rect 9673 11522 9739 11525
rect 12065 11522 12131 11525
rect 9673 11520 12131 11522
rect 9673 11464 9678 11520
rect 9734 11464 12070 11520
rect 12126 11464 12131 11520
rect 9673 11462 12131 11464
rect 9673 11459 9739 11462
rect 12065 11459 12131 11462
rect 12341 11522 12407 11525
rect 12525 11522 12591 11525
rect 12341 11520 12591 11522
rect 12341 11464 12346 11520
rect 12402 11464 12530 11520
rect 12586 11464 12591 11520
rect 12341 11462 12591 11464
rect 12341 11459 12407 11462
rect 12525 11459 12591 11462
rect 7808 11456 8128 11457
rect 0 11386 800 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 4797 11386 4863 11389
rect 0 11384 4863 11386
rect 0 11328 4802 11384
rect 4858 11328 4863 11384
rect 0 11326 4863 11328
rect 0 11296 800 11326
rect 4797 11323 4863 11326
rect 10041 11386 10107 11389
rect 14273 11386 14339 11389
rect 10041 11384 14339 11386
rect 10041 11328 10046 11384
rect 10102 11328 14278 11384
rect 14334 11328 14339 11384
rect 10041 11326 14339 11328
rect 10041 11323 10107 11326
rect 14273 11323 14339 11326
rect 2497 11250 2563 11253
rect 13629 11250 13695 11253
rect 2497 11248 13695 11250
rect 2497 11192 2502 11248
rect 2558 11192 13634 11248
rect 13690 11192 13695 11248
rect 2497 11190 13695 11192
rect 2497 11187 2563 11190
rect 13629 11187 13695 11190
rect 6821 11114 6887 11117
rect 11237 11114 11303 11117
rect 6821 11112 11303 11114
rect 6821 11056 6826 11112
rect 6882 11056 11242 11112
rect 11298 11056 11303 11112
rect 6821 11054 11303 11056
rect 6821 11051 6887 11054
rect 11237 11051 11303 11054
rect 4376 10912 4696 10913
rect 0 10842 800 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3693 10842 3759 10845
rect 0 10840 3759 10842
rect 0 10784 3698 10840
rect 3754 10784 3759 10840
rect 0 10782 3759 10784
rect 0 10752 800 10782
rect 3693 10779 3759 10782
rect 10501 10706 10567 10709
rect 13813 10706 13879 10709
rect 10501 10704 13879 10706
rect 10501 10648 10506 10704
rect 10562 10648 13818 10704
rect 13874 10648 13879 10704
rect 10501 10646 13879 10648
rect 10501 10643 10567 10646
rect 13813 10643 13879 10646
rect 4797 10570 4863 10573
rect 18137 10570 18203 10573
rect 4797 10568 18203 10570
rect 4797 10512 4802 10568
rect 4858 10512 18142 10568
rect 18198 10512 18203 10568
rect 4797 10510 18203 10512
rect 4797 10507 4863 10510
rect 18137 10507 18203 10510
rect 0 10434 800 10464
rect 4797 10434 4863 10437
rect 0 10432 4863 10434
rect 0 10376 4802 10432
rect 4858 10376 4863 10432
rect 0 10374 4863 10376
rect 0 10344 800 10374
rect 4797 10371 4863 10374
rect 8569 10434 8635 10437
rect 10593 10434 10659 10437
rect 12065 10434 12131 10437
rect 8569 10432 10426 10434
rect 8569 10376 8574 10432
rect 8630 10376 10426 10432
rect 8569 10374 10426 10376
rect 8569 10371 8635 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 10366 10298 10426 10374
rect 10593 10432 12131 10434
rect 10593 10376 10598 10432
rect 10654 10376 12070 10432
rect 12126 10376 12131 10432
rect 10593 10374 12131 10376
rect 10593 10371 10659 10374
rect 12065 10371 12131 10374
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 12157 10298 12223 10301
rect 10366 10296 12223 10298
rect 10366 10240 12162 10296
rect 12218 10240 12223 10296
rect 10366 10238 12223 10240
rect 12157 10235 12223 10238
rect 4061 10162 4127 10165
rect 11329 10162 11395 10165
rect 4061 10160 11395 10162
rect 4061 10104 4066 10160
rect 4122 10104 11334 10160
rect 11390 10104 11395 10160
rect 4061 10102 11395 10104
rect 4061 10099 4127 10102
rect 11329 10099 11395 10102
rect 0 10026 800 10056
rect 3969 10026 4035 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 800 9966
rect 3969 9963 4035 9966
rect 4797 10026 4863 10029
rect 9029 10026 9095 10029
rect 4797 10024 9095 10026
rect 4797 9968 4802 10024
rect 4858 9968 9034 10024
rect 9090 9968 9095 10024
rect 4797 9966 9095 9968
rect 4797 9963 4863 9966
rect 9029 9963 9095 9966
rect 13629 10026 13695 10029
rect 14181 10026 14247 10029
rect 13629 10024 14247 10026
rect 13629 9968 13634 10024
rect 13690 9968 14186 10024
rect 14242 9968 14247 10024
rect 13629 9966 14247 9968
rect 13629 9963 13695 9966
rect 14181 9963 14247 9966
rect 5165 9890 5231 9893
rect 7833 9890 7899 9893
rect 5165 9888 7899 9890
rect 5165 9832 5170 9888
rect 5226 9832 7838 9888
rect 7894 9832 7899 9888
rect 5165 9830 7899 9832
rect 5165 9827 5231 9830
rect 7833 9827 7899 9830
rect 11789 9890 11855 9893
rect 15653 9890 15719 9893
rect 11789 9888 15719 9890
rect 11789 9832 11794 9888
rect 11850 9832 15658 9888
rect 15714 9832 15719 9888
rect 11789 9830 15719 9832
rect 11789 9827 11855 9830
rect 15653 9827 15719 9830
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 2681 9618 2747 9621
rect 5257 9618 5323 9621
rect 2681 9616 5323 9618
rect 2681 9560 2686 9616
rect 2742 9560 5262 9616
rect 5318 9560 5323 9616
rect 2681 9558 5323 9560
rect 2681 9555 2747 9558
rect 5257 9555 5323 9558
rect 6361 9618 6427 9621
rect 7833 9618 7899 9621
rect 6361 9616 7899 9618
rect 6361 9560 6366 9616
rect 6422 9560 7838 9616
rect 7894 9560 7899 9616
rect 6361 9558 7899 9560
rect 6361 9555 6427 9558
rect 7833 9555 7899 9558
rect 11697 9618 11763 9621
rect 14273 9618 14339 9621
rect 11697 9616 14339 9618
rect 11697 9560 11702 9616
rect 11758 9560 14278 9616
rect 14334 9560 14339 9616
rect 11697 9558 14339 9560
rect 11697 9555 11763 9558
rect 14273 9555 14339 9558
rect 0 9482 800 9512
rect 2865 9482 2931 9485
rect 0 9480 2931 9482
rect 0 9424 2870 9480
rect 2926 9424 2931 9480
rect 0 9422 2931 9424
rect 0 9392 800 9422
rect 2865 9419 2931 9422
rect 3509 9482 3575 9485
rect 13445 9482 13511 9485
rect 14641 9482 14707 9485
rect 3509 9480 14707 9482
rect 3509 9424 3514 9480
rect 3570 9424 13450 9480
rect 13506 9424 14646 9480
rect 14702 9424 14707 9480
rect 3509 9422 14707 9424
rect 3509 9419 3575 9422
rect 13445 9419 13511 9422
rect 14641 9419 14707 9422
rect 2313 9346 2379 9349
rect 7373 9346 7439 9349
rect 2313 9344 7439 9346
rect 2313 9288 2318 9344
rect 2374 9288 7378 9344
rect 7434 9288 7439 9344
rect 2313 9286 7439 9288
rect 2313 9283 2379 9286
rect 7373 9283 7439 9286
rect 11145 9346 11211 9349
rect 13169 9346 13235 9349
rect 11145 9344 13235 9346
rect 11145 9288 11150 9344
rect 11206 9288 13174 9344
rect 13230 9288 13235 9344
rect 11145 9286 13235 9288
rect 11145 9283 11211 9286
rect 13169 9283 13235 9286
rect 13445 9346 13511 9349
rect 13813 9346 13879 9349
rect 13445 9344 13879 9346
rect 13445 9288 13450 9344
rect 13506 9288 13818 9344
rect 13874 9288 13879 9344
rect 13445 9286 13879 9288
rect 13445 9283 13511 9286
rect 13813 9283 13879 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 2405 9210 2471 9213
rect 6729 9210 6795 9213
rect 2405 9208 6795 9210
rect 2405 9152 2410 9208
rect 2466 9152 6734 9208
rect 6790 9152 6795 9208
rect 2405 9150 6795 9152
rect 2405 9147 2471 9150
rect 6729 9147 6795 9150
rect 0 9074 800 9104
rect 2129 9074 2195 9077
rect 0 9072 2195 9074
rect 0 9016 2134 9072
rect 2190 9016 2195 9072
rect 0 9014 2195 9016
rect 0 8984 800 9014
rect 2129 9011 2195 9014
rect 6545 9074 6611 9077
rect 15193 9074 15259 9077
rect 6545 9072 15259 9074
rect 6545 9016 6550 9072
rect 6606 9016 15198 9072
rect 15254 9016 15259 9072
rect 6545 9014 15259 9016
rect 6545 9011 6611 9014
rect 15193 9011 15259 9014
rect 3969 8938 4035 8941
rect 5993 8938 6059 8941
rect 7230 8938 7236 8940
rect 3969 8936 4860 8938
rect 3969 8880 3974 8936
rect 4030 8880 4860 8936
rect 3969 8878 4860 8880
rect 3969 8875 4035 8878
rect 4800 8802 4860 8878
rect 5993 8936 7236 8938
rect 5993 8880 5998 8936
rect 6054 8880 7236 8936
rect 5993 8878 7236 8880
rect 5993 8875 6059 8878
rect 7230 8876 7236 8878
rect 7300 8938 7306 8940
rect 9765 8938 9831 8941
rect 9949 8938 10015 8941
rect 7300 8936 10015 8938
rect 7300 8880 9770 8936
rect 9826 8880 9954 8936
rect 10010 8880 10015 8936
rect 7300 8878 10015 8880
rect 7300 8876 7306 8878
rect 9765 8875 9831 8878
rect 9949 8875 10015 8878
rect 10777 8938 10843 8941
rect 16113 8938 16179 8941
rect 10777 8936 16179 8938
rect 10777 8880 10782 8936
rect 10838 8880 16118 8936
rect 16174 8880 16179 8936
rect 10777 8878 16179 8880
rect 10777 8875 10843 8878
rect 16113 8875 16179 8878
rect 9029 8802 9095 8805
rect 4800 8800 9095 8802
rect 4800 8744 9034 8800
rect 9090 8744 9095 8800
rect 4800 8742 9095 8744
rect 9029 8739 9095 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 6177 8668 6243 8669
rect 6126 8604 6132 8668
rect 6196 8666 6243 8668
rect 9397 8666 9463 8669
rect 6196 8664 9463 8666
rect 6238 8608 9402 8664
rect 9458 8608 9463 8664
rect 6196 8606 9463 8608
rect 6196 8604 6243 8606
rect 6177 8603 6243 8604
rect 9397 8603 9463 8606
rect 9949 8666 10015 8669
rect 10869 8666 10935 8669
rect 9949 8664 10935 8666
rect 9949 8608 9954 8664
rect 10010 8608 10874 8664
rect 10930 8608 10935 8664
rect 9949 8606 10935 8608
rect 9949 8603 10015 8606
rect 10869 8603 10935 8606
rect 17534 8604 17540 8668
rect 17604 8666 17610 8668
rect 17861 8666 17927 8669
rect 17604 8664 17927 8666
rect 17604 8608 17866 8664
rect 17922 8608 17927 8664
rect 17604 8606 17927 8608
rect 17604 8604 17610 8606
rect 17861 8603 17927 8606
rect 0 8530 800 8560
rect 10777 8530 10843 8533
rect 0 8528 10843 8530
rect 0 8472 10782 8528
rect 10838 8472 10843 8528
rect 0 8470 10843 8472
rect 0 8440 800 8470
rect 10777 8467 10843 8470
rect 14181 8530 14247 8533
rect 15469 8530 15535 8533
rect 14181 8528 15535 8530
rect 14181 8472 14186 8528
rect 14242 8472 15474 8528
rect 15530 8472 15535 8528
rect 14181 8470 15535 8472
rect 14181 8467 14247 8470
rect 15469 8467 15535 8470
rect 8569 8394 8635 8397
rect 8845 8394 8911 8397
rect 5766 8334 8402 8394
rect 3417 8258 3483 8261
rect 5766 8258 5826 8334
rect 3417 8256 5826 8258
rect 3417 8200 3422 8256
rect 3478 8200 5826 8256
rect 3417 8198 5826 8200
rect 8342 8258 8402 8334
rect 8569 8392 8911 8394
rect 8569 8336 8574 8392
rect 8630 8336 8850 8392
rect 8906 8336 8911 8392
rect 8569 8334 8911 8336
rect 8569 8331 8635 8334
rect 8845 8331 8911 8334
rect 10961 8394 11027 8397
rect 16481 8394 16547 8397
rect 10961 8392 16547 8394
rect 10961 8336 10966 8392
rect 11022 8336 16486 8392
rect 16542 8336 16547 8392
rect 10961 8334 16547 8336
rect 10961 8331 11027 8334
rect 16481 8331 16547 8334
rect 16941 8394 17007 8397
rect 17309 8394 17375 8397
rect 17585 8396 17651 8397
rect 16941 8392 17375 8394
rect 16941 8336 16946 8392
rect 17002 8336 17314 8392
rect 17370 8336 17375 8392
rect 16941 8334 17375 8336
rect 16941 8331 17007 8334
rect 17309 8331 17375 8334
rect 17534 8332 17540 8396
rect 17604 8394 17651 8396
rect 17604 8392 17696 8394
rect 17646 8336 17696 8392
rect 17604 8334 17696 8336
rect 17604 8332 17651 8334
rect 17585 8331 17651 8332
rect 11881 8258 11947 8261
rect 8342 8256 11947 8258
rect 8342 8200 11886 8256
rect 11942 8200 11947 8256
rect 8342 8198 11947 8200
rect 3417 8195 3483 8198
rect 11881 8195 11947 8198
rect 18137 8256 18203 8261
rect 18137 8200 18142 8256
rect 18198 8200 18203 8256
rect 18137 8195 18203 8200
rect 7808 8192 8128 8193
rect 0 8122 800 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 6821 8122 6887 8125
rect 0 8120 6887 8122
rect 0 8064 6826 8120
rect 6882 8064 6887 8120
rect 0 8062 6887 8064
rect 0 8032 800 8062
rect 6821 8059 6887 8062
rect 8334 8060 8340 8124
rect 8404 8122 8410 8124
rect 14181 8122 14247 8125
rect 8404 8120 14247 8122
rect 8404 8064 14186 8120
rect 14242 8064 14247 8120
rect 8404 8062 14247 8064
rect 8404 8060 8410 8062
rect 14181 8059 14247 8062
rect 16757 8122 16823 8125
rect 18140 8122 18200 8195
rect 16757 8120 18200 8122
rect 16757 8064 16762 8120
rect 16818 8064 18200 8120
rect 16757 8062 18200 8064
rect 16757 8059 16823 8062
rect 4889 7986 4955 7989
rect 8293 7986 8359 7989
rect 4889 7984 8359 7986
rect 4889 7928 4894 7984
rect 4950 7928 8298 7984
rect 8354 7928 8359 7984
rect 4889 7926 8359 7928
rect 4889 7923 4955 7926
rect 8293 7923 8359 7926
rect 10869 7986 10935 7989
rect 18781 7986 18847 7989
rect 10869 7984 18847 7986
rect 10869 7928 10874 7984
rect 10930 7928 18786 7984
rect 18842 7928 18847 7984
rect 10869 7926 18847 7928
rect 10869 7923 10935 7926
rect 18781 7923 18847 7926
rect 2497 7850 2563 7853
rect 7097 7850 7163 7853
rect 2497 7848 7163 7850
rect 2497 7792 2502 7848
rect 2558 7792 7102 7848
rect 7158 7792 7163 7848
rect 2497 7790 7163 7792
rect 2497 7787 2563 7790
rect 7097 7787 7163 7790
rect 7281 7850 7347 7853
rect 8334 7850 8340 7852
rect 7281 7848 8340 7850
rect 7281 7792 7286 7848
rect 7342 7792 8340 7848
rect 7281 7790 8340 7792
rect 7281 7787 7347 7790
rect 8334 7788 8340 7790
rect 8404 7788 8410 7852
rect 11605 7850 11671 7853
rect 18505 7850 18571 7853
rect 11605 7848 18571 7850
rect 11605 7792 11610 7848
rect 11666 7792 18510 7848
rect 18566 7792 18571 7848
rect 11605 7790 18571 7792
rect 11605 7787 11671 7790
rect 18505 7787 18571 7790
rect 4797 7714 4863 7717
rect 6913 7714 6979 7717
rect 8017 7714 8083 7717
rect 4797 7712 6378 7714
rect 4797 7656 4802 7712
rect 4858 7656 6378 7712
rect 4797 7654 6378 7656
rect 4797 7651 4863 7654
rect 4376 7648 4696 7649
rect 0 7578 800 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 800 7518
rect 4061 7515 4127 7518
rect 5625 7578 5691 7581
rect 6177 7578 6243 7581
rect 5625 7576 6243 7578
rect 5625 7520 5630 7576
rect 5686 7520 6182 7576
rect 6238 7520 6243 7576
rect 5625 7518 6243 7520
rect 6318 7578 6378 7654
rect 6913 7712 8083 7714
rect 6913 7656 6918 7712
rect 6974 7656 8022 7712
rect 8078 7656 8083 7712
rect 6913 7654 8083 7656
rect 6913 7651 6979 7654
rect 8017 7651 8083 7654
rect 14181 7714 14247 7717
rect 15561 7714 15627 7717
rect 14181 7712 15627 7714
rect 14181 7656 14186 7712
rect 14242 7656 15566 7712
rect 15622 7656 15627 7712
rect 14181 7654 15627 7656
rect 14181 7651 14247 7654
rect 15561 7651 15627 7654
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 10869 7578 10935 7581
rect 6318 7576 10935 7578
rect 6318 7520 10874 7576
rect 10930 7520 10935 7576
rect 6318 7518 10935 7520
rect 5625 7515 5691 7518
rect 6177 7515 6243 7518
rect 10869 7515 10935 7518
rect 11881 7578 11947 7581
rect 17953 7578 18019 7581
rect 11881 7576 18019 7578
rect 11881 7520 11886 7576
rect 11942 7520 17958 7576
rect 18014 7520 18019 7576
rect 11881 7518 18019 7520
rect 11881 7515 11947 7518
rect 17953 7515 18019 7518
rect 4705 7442 4771 7445
rect 19793 7442 19859 7445
rect 4705 7440 19859 7442
rect 4705 7384 4710 7440
rect 4766 7384 19798 7440
rect 19854 7384 19859 7440
rect 4705 7382 19859 7384
rect 4705 7379 4771 7382
rect 19793 7379 19859 7382
rect 3141 7306 3207 7309
rect 3417 7306 3483 7309
rect 3141 7304 3483 7306
rect 3141 7248 3146 7304
rect 3202 7248 3422 7304
rect 3478 7248 3483 7304
rect 3141 7246 3483 7248
rect 3141 7243 3207 7246
rect 3417 7243 3483 7246
rect 7097 7306 7163 7309
rect 14273 7306 14339 7309
rect 20161 7306 20227 7309
rect 7097 7304 14339 7306
rect 7097 7248 7102 7304
rect 7158 7248 14278 7304
rect 14334 7248 14339 7304
rect 7097 7246 14339 7248
rect 7097 7243 7163 7246
rect 14273 7243 14339 7246
rect 14414 7304 20227 7306
rect 14414 7248 20166 7304
rect 20222 7248 20227 7304
rect 14414 7246 20227 7248
rect 0 7170 800 7200
rect 3969 7170 4035 7173
rect 0 7168 4035 7170
rect 0 7112 3974 7168
rect 4030 7112 4035 7168
rect 0 7110 4035 7112
rect 0 7080 800 7110
rect 3969 7107 4035 7110
rect 8293 7170 8359 7173
rect 11605 7170 11671 7173
rect 14414 7170 14474 7246
rect 20161 7243 20227 7246
rect 8293 7168 11671 7170
rect 8293 7112 8298 7168
rect 8354 7112 11610 7168
rect 11666 7112 11671 7168
rect 8293 7110 11671 7112
rect 8293 7107 8359 7110
rect 11605 7107 11671 7110
rect 12206 7110 14474 7170
rect 15285 7170 15351 7173
rect 17953 7170 18019 7173
rect 15285 7168 18019 7170
rect 15285 7112 15290 7168
rect 15346 7112 17958 7168
rect 18014 7112 18019 7168
rect 15285 7110 18019 7112
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 4429 7034 4495 7037
rect 4429 7032 6746 7034
rect 4429 6976 4434 7032
rect 4490 6976 6746 7032
rect 4429 6974 6746 6976
rect 4429 6971 4495 6974
rect 4061 6898 4127 6901
rect 6177 6898 6243 6901
rect 6361 6898 6427 6901
rect 4061 6896 6427 6898
rect 4061 6840 4066 6896
rect 4122 6840 6182 6896
rect 6238 6840 6366 6896
rect 6422 6840 6427 6896
rect 4061 6838 6427 6840
rect 6686 6898 6746 6974
rect 12206 6898 12266 7110
rect 15285 7107 15351 7110
rect 17953 7107 18019 7110
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 14273 7034 14339 7037
rect 19333 7034 19399 7037
rect 14273 7032 14474 7034
rect 14273 6976 14278 7032
rect 14334 6976 14474 7032
rect 14273 6974 14474 6976
rect 14273 6971 14339 6974
rect 6686 6838 12266 6898
rect 12617 6898 12683 6901
rect 14089 6898 14155 6901
rect 12617 6896 14155 6898
rect 12617 6840 12622 6896
rect 12678 6840 14094 6896
rect 14150 6840 14155 6896
rect 12617 6838 14155 6840
rect 14414 6898 14474 6974
rect 15150 7032 19399 7034
rect 15150 6976 19338 7032
rect 19394 6976 19399 7032
rect 15150 6974 19399 6976
rect 15150 6898 15210 6974
rect 19333 6971 19399 6974
rect 14414 6838 15210 6898
rect 17953 6898 18019 6901
rect 18597 6898 18663 6901
rect 17953 6896 18663 6898
rect 17953 6840 17958 6896
rect 18014 6840 18602 6896
rect 18658 6840 18663 6896
rect 17953 6838 18663 6840
rect 4061 6835 4127 6838
rect 6177 6835 6243 6838
rect 6361 6835 6427 6838
rect 12617 6835 12683 6838
rect 14089 6835 14155 6838
rect 17953 6835 18019 6838
rect 18597 6835 18663 6838
rect 0 6762 800 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 800 6702
rect 4061 6699 4127 6702
rect 4705 6762 4771 6765
rect 18413 6762 18479 6765
rect 4705 6760 18479 6762
rect 4705 6704 4710 6760
rect 4766 6704 18418 6760
rect 18474 6704 18479 6760
rect 4705 6702 18479 6704
rect 4705 6699 4771 6702
rect 18413 6699 18479 6702
rect 19517 6764 19583 6765
rect 19517 6760 19564 6764
rect 19628 6762 19634 6764
rect 19517 6704 19522 6760
rect 19517 6700 19564 6704
rect 19628 6702 19674 6762
rect 19628 6700 19634 6702
rect 19517 6699 19583 6700
rect 13445 6626 13511 6629
rect 14273 6626 14339 6629
rect 13445 6624 14339 6626
rect 13445 6568 13450 6624
rect 13506 6568 14278 6624
rect 14334 6568 14339 6624
rect 13445 6566 14339 6568
rect 13445 6563 13511 6566
rect 14273 6563 14339 6566
rect 15745 6626 15811 6629
rect 16941 6626 17007 6629
rect 15745 6624 17007 6626
rect 15745 6568 15750 6624
rect 15806 6568 16946 6624
rect 17002 6568 17007 6624
rect 15745 6566 17007 6568
rect 15745 6563 15811 6566
rect 16941 6563 17007 6566
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 11789 6490 11855 6493
rect 16665 6490 16731 6493
rect 11789 6488 16731 6490
rect 11789 6432 11794 6488
rect 11850 6432 16670 6488
rect 16726 6432 16731 6488
rect 11789 6430 16731 6432
rect 11789 6427 11855 6430
rect 16665 6427 16731 6430
rect 18638 6428 18644 6492
rect 18708 6490 18714 6492
rect 18873 6490 18939 6493
rect 18708 6488 18939 6490
rect 18708 6432 18878 6488
rect 18934 6432 18939 6488
rect 18708 6430 18939 6432
rect 18708 6428 18714 6430
rect 18873 6427 18939 6430
rect 11881 6354 11947 6357
rect 12525 6354 12591 6357
rect 11881 6352 12591 6354
rect 11881 6296 11886 6352
rect 11942 6296 12530 6352
rect 12586 6296 12591 6352
rect 11881 6294 12591 6296
rect 11881 6291 11947 6294
rect 12525 6291 12591 6294
rect 13445 6354 13511 6357
rect 17769 6354 17835 6357
rect 13445 6352 17835 6354
rect 13445 6296 13450 6352
rect 13506 6296 17774 6352
rect 17830 6296 17835 6352
rect 13445 6294 17835 6296
rect 13445 6291 13511 6294
rect 17769 6291 17835 6294
rect 18781 6354 18847 6357
rect 19149 6354 19215 6357
rect 18781 6352 19215 6354
rect 18781 6296 18786 6352
rect 18842 6296 19154 6352
rect 19210 6296 19215 6352
rect 18781 6294 19215 6296
rect 18781 6291 18847 6294
rect 19149 6291 19215 6294
rect 0 6218 800 6248
rect 3877 6218 3943 6221
rect 0 6216 3943 6218
rect 0 6160 3882 6216
rect 3938 6160 3943 6216
rect 0 6158 3943 6160
rect 0 6128 800 6158
rect 3877 6155 3943 6158
rect 6821 6218 6887 6221
rect 17953 6218 18019 6221
rect 6821 6216 18019 6218
rect 6821 6160 6826 6216
rect 6882 6160 17958 6216
rect 18014 6160 18019 6216
rect 6821 6158 18019 6160
rect 6821 6155 6887 6158
rect 17953 6155 18019 6158
rect 9765 6082 9831 6085
rect 11145 6082 11211 6085
rect 9765 6080 11211 6082
rect 9765 6024 9770 6080
rect 9826 6024 11150 6080
rect 11206 6024 11211 6080
rect 9765 6022 11211 6024
rect 9765 6019 9831 6022
rect 11145 6019 11211 6022
rect 17677 6082 17743 6085
rect 21265 6082 21331 6085
rect 17677 6080 21331 6082
rect 17677 6024 17682 6080
rect 17738 6024 21270 6080
rect 21326 6024 21331 6080
rect 17677 6022 21331 6024
rect 17677 6019 17743 6022
rect 21265 6019 21331 6022
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 3601 5946 3667 5949
rect 6637 5946 6703 5949
rect 3601 5944 6703 5946
rect 3601 5888 3606 5944
rect 3662 5888 6642 5944
rect 6698 5888 6703 5944
rect 3601 5886 6703 5888
rect 3601 5883 3667 5886
rect 6637 5883 6703 5886
rect 9673 5946 9739 5949
rect 13721 5946 13787 5949
rect 9673 5944 13787 5946
rect 9673 5888 9678 5944
rect 9734 5888 13726 5944
rect 13782 5888 13787 5944
rect 9673 5886 13787 5888
rect 9673 5883 9739 5886
rect 13721 5883 13787 5886
rect 16941 5946 17007 5949
rect 18045 5946 18111 5949
rect 16941 5944 18111 5946
rect 16941 5888 16946 5944
rect 17002 5888 18050 5944
rect 18106 5888 18111 5944
rect 16941 5886 18111 5888
rect 16941 5883 17007 5886
rect 18045 5883 18111 5886
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 5625 5810 5691 5813
rect 7189 5810 7255 5813
rect 8293 5810 8359 5813
rect 5625 5808 8359 5810
rect 5625 5752 5630 5808
rect 5686 5752 7194 5808
rect 7250 5752 8298 5808
rect 8354 5752 8359 5808
rect 5625 5750 8359 5752
rect 5625 5747 5691 5750
rect 7189 5747 7255 5750
rect 8293 5747 8359 5750
rect 10777 5810 10843 5813
rect 12801 5810 12867 5813
rect 17769 5810 17835 5813
rect 10777 5808 12082 5810
rect 10777 5752 10782 5808
rect 10838 5752 12082 5808
rect 10777 5750 12082 5752
rect 10777 5747 10843 5750
rect 3969 5674 4035 5677
rect 6126 5674 6132 5676
rect 3969 5672 6132 5674
rect 3969 5616 3974 5672
rect 4030 5616 6132 5672
rect 3969 5614 6132 5616
rect 3969 5611 4035 5614
rect 6126 5612 6132 5614
rect 6196 5612 6202 5676
rect 6637 5674 6703 5677
rect 8569 5674 8635 5677
rect 6637 5672 8635 5674
rect 6637 5616 6642 5672
rect 6698 5616 8574 5672
rect 8630 5616 8635 5672
rect 6637 5614 8635 5616
rect 6637 5611 6703 5614
rect 8569 5611 8635 5614
rect 11102 5614 11714 5674
rect 6453 5538 6519 5541
rect 11102 5538 11162 5614
rect 6453 5536 11162 5538
rect 6453 5480 6458 5536
rect 6514 5480 11162 5536
rect 6453 5478 11162 5480
rect 6453 5475 6519 5478
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 11654 5402 11714 5614
rect 12022 5538 12082 5750
rect 12801 5808 17835 5810
rect 12801 5752 12806 5808
rect 12862 5752 17774 5808
rect 17830 5752 17835 5808
rect 12801 5750 17835 5752
rect 12801 5747 12867 5750
rect 17769 5747 17835 5750
rect 19425 5810 19491 5813
rect 22000 5810 22800 5840
rect 19425 5808 22800 5810
rect 19425 5752 19430 5808
rect 19486 5752 22800 5808
rect 19425 5750 22800 5752
rect 19425 5747 19491 5750
rect 22000 5720 22800 5750
rect 12157 5674 12223 5677
rect 12617 5674 12683 5677
rect 12157 5672 12683 5674
rect 12157 5616 12162 5672
rect 12218 5616 12622 5672
rect 12678 5616 12683 5672
rect 12157 5614 12683 5616
rect 12157 5611 12223 5614
rect 12617 5611 12683 5614
rect 13537 5674 13603 5677
rect 17125 5674 17191 5677
rect 13537 5672 17191 5674
rect 13537 5616 13542 5672
rect 13598 5616 17130 5672
rect 17186 5616 17191 5672
rect 13537 5614 17191 5616
rect 13537 5611 13603 5614
rect 17125 5611 17191 5614
rect 15009 5538 15075 5541
rect 12022 5536 15075 5538
rect 12022 5480 15014 5536
rect 15070 5480 15075 5536
rect 12022 5478 15075 5480
rect 15009 5475 15075 5478
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 17585 5402 17651 5405
rect 11654 5400 17651 5402
rect 11654 5344 17590 5400
rect 17646 5344 17651 5400
rect 11654 5342 17651 5344
rect 17585 5339 17651 5342
rect 0 5266 800 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 800 5206
rect 4061 5203 4127 5206
rect 6821 5266 6887 5269
rect 13813 5266 13879 5269
rect 20161 5266 20227 5269
rect 6821 5264 13738 5266
rect 6821 5208 6826 5264
rect 6882 5208 13738 5264
rect 6821 5206 13738 5208
rect 6821 5203 6887 5206
rect 3141 5130 3207 5133
rect 9949 5130 10015 5133
rect 12065 5130 12131 5133
rect 3141 5128 9874 5130
rect 3141 5072 3146 5128
rect 3202 5072 9874 5128
rect 3141 5070 9874 5072
rect 3141 5067 3207 5070
rect 9814 4994 9874 5070
rect 9949 5128 12131 5130
rect 9949 5072 9954 5128
rect 10010 5072 12070 5128
rect 12126 5072 12131 5128
rect 9949 5070 12131 5072
rect 13678 5130 13738 5206
rect 13813 5264 20227 5266
rect 13813 5208 13818 5264
rect 13874 5208 20166 5264
rect 20222 5208 20227 5264
rect 13813 5206 20227 5208
rect 13813 5203 13879 5206
rect 20161 5203 20227 5206
rect 19374 5130 19380 5132
rect 13678 5070 19380 5130
rect 9949 5067 10015 5070
rect 12065 5067 12131 5070
rect 19374 5068 19380 5070
rect 19444 5068 19450 5132
rect 14273 4994 14339 4997
rect 9814 4992 14339 4994
rect 9814 4936 14278 4992
rect 14334 4936 14339 4992
rect 9814 4934 14339 4936
rect 14273 4931 14339 4934
rect 15377 4994 15443 4997
rect 16021 4994 16087 4997
rect 16481 4994 16547 4997
rect 18689 4994 18755 4997
rect 15377 4992 18755 4994
rect 15377 4936 15382 4992
rect 15438 4936 16026 4992
rect 16082 4936 16486 4992
rect 16542 4936 18694 4992
rect 18750 4936 18755 4992
rect 15377 4934 18755 4936
rect 15377 4931 15443 4934
rect 16021 4931 16087 4934
rect 16481 4931 16547 4934
rect 18689 4931 18755 4934
rect 7808 4928 8128 4929
rect 0 4858 800 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 2221 4858 2287 4861
rect 12433 4858 12499 4861
rect 13537 4858 13603 4861
rect 0 4856 2287 4858
rect 0 4800 2226 4856
rect 2282 4800 2287 4856
rect 0 4798 2287 4800
rect 0 4768 800 4798
rect 2221 4795 2287 4798
rect 9446 4856 13603 4858
rect 9446 4800 12438 4856
rect 12494 4800 13542 4856
rect 13598 4800 13603 4856
rect 9446 4798 13603 4800
rect 6361 4722 6427 4725
rect 9446 4722 9506 4798
rect 12433 4795 12499 4798
rect 13537 4795 13603 4798
rect 15101 4858 15167 4861
rect 18597 4858 18663 4861
rect 15101 4856 18663 4858
rect 15101 4800 15106 4856
rect 15162 4800 18602 4856
rect 18658 4800 18663 4856
rect 15101 4798 18663 4800
rect 15101 4795 15167 4798
rect 18597 4795 18663 4798
rect 6361 4720 9506 4722
rect 6361 4664 6366 4720
rect 6422 4664 9506 4720
rect 6361 4662 9506 4664
rect 9581 4722 9647 4725
rect 21173 4722 21239 4725
rect 9581 4720 21239 4722
rect 9581 4664 9586 4720
rect 9642 4664 21178 4720
rect 21234 4664 21239 4720
rect 9581 4662 21239 4664
rect 6361 4659 6427 4662
rect 9581 4659 9647 4662
rect 21173 4659 21239 4662
rect 2773 4586 2839 4589
rect 3233 4586 3299 4589
rect 20805 4586 20871 4589
rect 2773 4584 20871 4586
rect 2773 4528 2778 4584
rect 2834 4528 3238 4584
rect 3294 4528 20810 4584
rect 20866 4528 20871 4584
rect 2773 4526 20871 4528
rect 2773 4523 2839 4526
rect 3233 4523 3299 4526
rect 20805 4523 20871 4526
rect 5349 4450 5415 4453
rect 7741 4450 7807 4453
rect 5349 4448 7807 4450
rect 5349 4392 5354 4448
rect 5410 4392 7746 4448
rect 7802 4392 7807 4448
rect 5349 4390 7807 4392
rect 5349 4387 5415 4390
rect 7741 4387 7807 4390
rect 8569 4450 8635 4453
rect 10961 4450 11027 4453
rect 8569 4448 11027 4450
rect 8569 4392 8574 4448
rect 8630 4392 10966 4448
rect 11022 4392 11027 4448
rect 8569 4390 11027 4392
rect 8569 4387 8635 4390
rect 10961 4387 11027 4390
rect 11973 4450 12039 4453
rect 13905 4450 13971 4453
rect 11973 4448 13971 4450
rect 11973 4392 11978 4448
rect 12034 4392 13910 4448
rect 13966 4392 13971 4448
rect 11973 4390 13971 4392
rect 11973 4387 12039 4390
rect 13905 4387 13971 4390
rect 4376 4384 4696 4385
rect 0 4314 800 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 9581 4314 9647 4317
rect 16757 4314 16823 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 800 4254
rect 4061 4251 4127 4254
rect 4846 4312 9647 4314
rect 4846 4256 9586 4312
rect 9642 4256 9647 4312
rect 4846 4254 9647 4256
rect 3509 4178 3575 4181
rect 4061 4178 4127 4181
rect 4846 4178 4906 4254
rect 9581 4251 9647 4254
rect 13126 4312 16823 4314
rect 13126 4256 16762 4312
rect 16818 4256 16823 4312
rect 13126 4254 16823 4256
rect 3509 4176 4906 4178
rect 3509 4120 3514 4176
rect 3570 4120 4066 4176
rect 4122 4120 4906 4176
rect 3509 4118 4906 4120
rect 5809 4178 5875 4181
rect 13126 4178 13186 4254
rect 16757 4251 16823 4254
rect 5809 4176 13186 4178
rect 5809 4120 5814 4176
rect 5870 4120 13186 4176
rect 5809 4118 13186 4120
rect 13537 4178 13603 4181
rect 20069 4178 20135 4181
rect 13537 4176 20135 4178
rect 13537 4120 13542 4176
rect 13598 4120 20074 4176
rect 20130 4120 20135 4176
rect 13537 4118 20135 4120
rect 3509 4115 3575 4118
rect 4061 4115 4127 4118
rect 5809 4115 5875 4118
rect 13537 4115 13603 4118
rect 20069 4115 20135 4118
rect 2773 4042 2839 4045
rect 16665 4042 16731 4045
rect 2773 4040 16731 4042
rect 2773 3984 2778 4040
rect 2834 3984 16670 4040
rect 16726 3984 16731 4040
rect 2773 3982 16731 3984
rect 2773 3979 2839 3982
rect 16665 3979 16731 3982
rect 0 3906 800 3936
rect 7598 3906 7604 3908
rect 0 3846 7604 3906
rect 0 3816 800 3846
rect 7598 3844 7604 3846
rect 7668 3844 7674 3908
rect 10593 3906 10659 3909
rect 11881 3906 11947 3909
rect 10593 3904 11947 3906
rect 10593 3848 10598 3904
rect 10654 3848 11886 3904
rect 11942 3848 11947 3904
rect 10593 3846 11947 3848
rect 10593 3843 10659 3846
rect 11881 3843 11947 3846
rect 15469 3906 15535 3909
rect 18321 3906 18387 3909
rect 15469 3904 18387 3906
rect 15469 3848 15474 3904
rect 15530 3848 18326 3904
rect 18382 3848 18387 3904
rect 15469 3846 18387 3848
rect 15469 3843 15535 3846
rect 18321 3843 18387 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 4889 3770 4955 3773
rect 7097 3770 7163 3773
rect 4889 3768 7163 3770
rect 4889 3712 4894 3768
rect 4950 3712 7102 3768
rect 7158 3712 7163 3768
rect 4889 3710 7163 3712
rect 4889 3707 4955 3710
rect 7097 3707 7163 3710
rect 15101 3770 15167 3773
rect 19517 3770 19583 3773
rect 15101 3768 19583 3770
rect 15101 3712 15106 3768
rect 15162 3712 19522 3768
rect 19578 3712 19583 3768
rect 15101 3710 19583 3712
rect 15101 3707 15167 3710
rect 19517 3707 19583 3710
rect 3877 3634 3943 3637
rect 4521 3634 4587 3637
rect 13537 3634 13603 3637
rect 3877 3632 13603 3634
rect 3877 3576 3882 3632
rect 3938 3576 4526 3632
rect 4582 3576 13542 3632
rect 13598 3576 13603 3632
rect 3877 3574 13603 3576
rect 3877 3571 3943 3574
rect 4521 3571 4587 3574
rect 13537 3571 13603 3574
rect 16665 3634 16731 3637
rect 19333 3634 19399 3637
rect 16665 3632 19399 3634
rect 16665 3576 16670 3632
rect 16726 3576 19338 3632
rect 19394 3576 19399 3632
rect 16665 3574 19399 3576
rect 16665 3571 16731 3574
rect 19333 3571 19399 3574
rect 0 3498 800 3528
rect 3049 3498 3115 3501
rect 0 3496 3115 3498
rect 0 3440 3054 3496
rect 3110 3440 3115 3496
rect 0 3438 3115 3440
rect 0 3408 800 3438
rect 3049 3435 3115 3438
rect 7598 3436 7604 3500
rect 7668 3498 7674 3500
rect 19977 3498 20043 3501
rect 7668 3496 20043 3498
rect 7668 3440 19982 3496
rect 20038 3440 20043 3496
rect 7668 3438 20043 3440
rect 7668 3436 7674 3438
rect 19977 3435 20043 3438
rect 5257 3362 5323 3365
rect 8385 3362 8451 3365
rect 5257 3360 8451 3362
rect 5257 3304 5262 3360
rect 5318 3304 8390 3360
rect 8446 3304 8451 3360
rect 5257 3302 8451 3304
rect 5257 3299 5323 3302
rect 8385 3299 8451 3302
rect 14457 3362 14523 3365
rect 17217 3362 17283 3365
rect 14457 3360 17283 3362
rect 14457 3304 14462 3360
rect 14518 3304 17222 3360
rect 17278 3304 17283 3360
rect 14457 3302 17283 3304
rect 14457 3299 14523 3302
rect 17217 3299 17283 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 8661 3226 8727 3229
rect 10409 3226 10475 3229
rect 11053 3226 11119 3229
rect 15653 3226 15719 3229
rect 8661 3224 11119 3226
rect 8661 3168 8666 3224
rect 8722 3168 10414 3224
rect 10470 3168 11058 3224
rect 11114 3168 11119 3224
rect 8661 3166 11119 3168
rect 8661 3163 8727 3166
rect 10409 3163 10475 3166
rect 11053 3163 11119 3166
rect 13310 3224 15719 3226
rect 13310 3168 15658 3224
rect 15714 3168 15719 3224
rect 13310 3166 15719 3168
rect 4705 3090 4771 3093
rect 13310 3090 13370 3166
rect 15653 3163 15719 3166
rect 15837 3226 15903 3229
rect 16113 3226 16179 3229
rect 18597 3228 18663 3229
rect 18597 3226 18644 3228
rect 15837 3224 16179 3226
rect 15837 3168 15842 3224
rect 15898 3168 16118 3224
rect 16174 3168 16179 3224
rect 15837 3166 16179 3168
rect 18552 3224 18644 3226
rect 18552 3168 18602 3224
rect 18552 3166 18644 3168
rect 15837 3163 15903 3166
rect 16113 3163 16179 3166
rect 18597 3164 18644 3166
rect 18708 3164 18714 3228
rect 18597 3163 18663 3164
rect 4705 3088 13370 3090
rect 4705 3032 4710 3088
rect 4766 3032 13370 3088
rect 4705 3030 13370 3032
rect 13537 3090 13603 3093
rect 19701 3090 19767 3093
rect 13537 3088 19767 3090
rect 13537 3032 13542 3088
rect 13598 3032 19706 3088
rect 19762 3032 19767 3088
rect 13537 3030 19767 3032
rect 4705 3027 4771 3030
rect 13537 3027 13603 3030
rect 19701 3027 19767 3030
rect 0 2954 800 2984
rect 2037 2954 2103 2957
rect 0 2952 2103 2954
rect 0 2896 2042 2952
rect 2098 2896 2103 2952
rect 0 2894 2103 2896
rect 0 2864 800 2894
rect 2037 2891 2103 2894
rect 4613 2954 4679 2957
rect 7281 2954 7347 2957
rect 14273 2954 14339 2957
rect 4613 2952 7347 2954
rect 4613 2896 4618 2952
rect 4674 2896 7286 2952
rect 7342 2896 7347 2952
rect 4613 2894 7347 2896
rect 4613 2891 4679 2894
rect 7281 2891 7347 2894
rect 7606 2952 14339 2954
rect 7606 2896 14278 2952
rect 14334 2896 14339 2952
rect 7606 2894 14339 2896
rect 2129 2818 2195 2821
rect 7606 2818 7666 2894
rect 14273 2891 14339 2894
rect 14825 2954 14891 2957
rect 16665 2954 16731 2957
rect 14825 2952 16731 2954
rect 14825 2896 14830 2952
rect 14886 2896 16670 2952
rect 16726 2896 16731 2952
rect 14825 2894 16731 2896
rect 14825 2891 14891 2894
rect 16665 2891 16731 2894
rect 2129 2816 7666 2818
rect 2129 2760 2134 2816
rect 2190 2760 7666 2816
rect 2129 2758 7666 2760
rect 8569 2818 8635 2821
rect 10869 2818 10935 2821
rect 8569 2816 10935 2818
rect 8569 2760 8574 2816
rect 8630 2760 10874 2816
rect 10930 2760 10935 2816
rect 8569 2758 10935 2760
rect 2129 2755 2195 2758
rect 8569 2755 8635 2758
rect 10869 2755 10935 2758
rect 15929 2818 15995 2821
rect 18873 2818 18939 2821
rect 15929 2816 18939 2818
rect 15929 2760 15934 2816
rect 15990 2760 18878 2816
rect 18934 2760 18939 2816
rect 15929 2758 18939 2760
rect 15929 2755 15995 2758
rect 18873 2755 18939 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 2773 2682 2839 2685
rect 6913 2682 6979 2685
rect 2773 2680 6979 2682
rect 2773 2624 2778 2680
rect 2834 2624 6918 2680
rect 6974 2624 6979 2680
rect 2773 2622 6979 2624
rect 2773 2619 2839 2622
rect 6913 2619 6979 2622
rect 0 2546 800 2576
rect 2405 2546 2471 2549
rect 0 2544 2471 2546
rect 0 2488 2410 2544
rect 2466 2488 2471 2544
rect 0 2486 2471 2488
rect 0 2456 800 2486
rect 2405 2483 2471 2486
rect 7373 2546 7439 2549
rect 16021 2546 16087 2549
rect 7373 2544 16087 2546
rect 7373 2488 7378 2544
rect 7434 2488 16026 2544
rect 16082 2488 16087 2544
rect 7373 2486 16087 2488
rect 7373 2483 7439 2486
rect 16021 2483 16087 2486
rect 10593 2410 10659 2413
rect 18137 2410 18203 2413
rect 10593 2408 18203 2410
rect 10593 2352 10598 2408
rect 10654 2352 18142 2408
rect 18198 2352 18203 2408
rect 10593 2350 18203 2352
rect 10593 2347 10659 2350
rect 18137 2347 18203 2350
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 0 1594 800 1624
rect 2589 1594 2655 1597
rect 0 1592 2655 1594
rect 0 1536 2594 1592
rect 2650 1536 2655 1592
rect 0 1534 2655 1536
rect 0 1504 800 1534
rect 2589 1531 2655 1534
rect 0 1050 800 1080
rect 1301 1050 1367 1053
rect 0 1048 1367 1050
rect 0 992 1306 1048
rect 1362 992 1367 1048
rect 0 990 1367 992
rect 0 960 800 990
rect 1301 987 1367 990
rect 0 642 800 672
rect 2221 642 2287 645
rect 0 640 2287 642
rect 0 584 2226 640
rect 2282 584 2287 640
rect 0 582 2287 584
rect 0 552 800 582
rect 2221 579 2287 582
rect 0 234 800 264
rect 1577 234 1643 237
rect 0 232 1643 234
rect 0 176 1582 232
rect 1638 176 1643 232
rect 0 174 1643 176
rect 0 144 800 174
rect 1577 171 1643 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7236 11460 7300 11524
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 7236 8876 7300 8940
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 6132 8664 6196 8668
rect 6132 8608 6182 8664
rect 6182 8608 6196 8664
rect 6132 8604 6196 8608
rect 17540 8604 17604 8668
rect 17540 8392 17604 8396
rect 17540 8336 17590 8392
rect 17590 8336 17604 8392
rect 17540 8332 17604 8336
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 8340 8060 8404 8124
rect 8340 7788 8404 7852
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 19564 6760 19628 6764
rect 19564 6704 19578 6760
rect 19578 6704 19628 6760
rect 19564 6700 19628 6704
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 18644 6428 18708 6492
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 6132 5612 6196 5676
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 19380 5068 19444 5132
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7604 3844 7668 3908
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 7604 3436 7668 3500
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 18644 3224 18708 3228
rect 18644 3168 18658 3224
rect 18658 3168 18708 3224
rect 18644 3164 18708 3168
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7235 11524 7301 11525
rect 7235 11460 7236 11524
rect 7300 11460 7301 11524
rect 7235 11459 7301 11460
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 7238 8941 7298 11459
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7235 8940 7301 8941
rect 7235 8876 7236 8940
rect 7300 8876 7301 8940
rect 7235 8875 7301 8876
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 6131 8668 6197 8669
rect 6131 8604 6132 8668
rect 6196 8604 6197 8668
rect 6131 8603 6197 8604
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 6134 5677 6194 8603
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 8339 8124 8405 8125
rect 8339 8060 8340 8124
rect 8404 8060 8405 8124
rect 8339 8059 8405 8060
rect 8342 7853 8402 8059
rect 8339 7852 8405 7853
rect 8339 7788 8340 7852
rect 8404 7788 8405 7852
rect 8339 7787 8405 7788
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 6131 5676 6197 5677
rect 6131 5612 6132 5676
rect 6196 5612 6197 5676
rect 6131 5611 6197 5612
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7603 3908 7669 3909
rect 7603 3844 7604 3908
rect 7668 3844 7669 3908
rect 7603 3843 7669 3844
rect 7606 3501 7666 3843
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7603 3500 7669 3501
rect 7603 3436 7604 3500
rect 7668 3436 7669 3500
rect 7603 3435 7669 3436
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 17539 8668 17605 8669
rect 17539 8604 17540 8668
rect 17604 8604 17605 8668
rect 17539 8603 17605 8604
rect 17542 8397 17602 8603
rect 17539 8396 17605 8397
rect 17539 8332 17540 8396
rect 17604 8332 17605 8396
rect 17539 8331 17605 8332
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 19563 6764 19629 6765
rect 19563 6700 19564 6764
rect 19628 6700 19629 6764
rect 19563 6699 19629 6700
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18643 6492 18709 6493
rect 18643 6428 18644 6492
rect 18708 6428 18709 6492
rect 18643 6427 18709 6428
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18646 3229 18706 6427
rect 19379 5132 19445 5133
rect 19379 5068 19380 5132
rect 19444 5130 19445 5132
rect 19566 5130 19626 6699
rect 19444 5070 19626 5130
rect 19444 5068 19445 5070
rect 19379 5067 19445 5068
rect 18643 3228 18709 3229
rect 18643 3164 18644 3228
rect 18708 3164 18709 3228
rect 18643 3163 18709 3164
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608763374
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608763374
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1608763374
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608763374
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1608763374
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608763374
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1608763374
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1608763374
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1608763374
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608763374
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1608763374
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1608763374
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1608763374
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608763374
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1608763374
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1608763374
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1608763374
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608763374
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1608763374
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1608763374
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1608763374
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1608763374
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608763374
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_52
timestamp 1608763374
transform 1 0 5888 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1608763374
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608763374
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1608763374
transform 1 0 3496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1608763374
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_24
timestamp 1608763374
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_28
timestamp 1608763374
transform 1 0 3680 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1608763374
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1608763374
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_40
timestamp 1608763374
transform 1 0 4784 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608763374
transform 1 0 2392 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608763374
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608763374
transform 1 0 2944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608763374
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1608763374
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1608763374
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1608763374
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_18
timestamp 1608763374
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608763374
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1608763374
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1608763374
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608763374
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1608763374
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1608763374
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1608763374
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1608763374
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1608763374
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608763374
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1608763374
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1608763374
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1608763374
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1608763374
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1608763374
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608763374
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1608763374
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1608763374
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_45
timestamp 1608763374
transform 1 0 5244 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1608763374
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1608763374
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1608763374
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1608763374
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1608763374
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1608763374
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_29
timestamp 1608763374
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp 1608763374
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1608763374
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1608763374
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608763374
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608763374
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2852 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608763374
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1608763374
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1608763374
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1608763374
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1608763374
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608763374
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608763374
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608763374
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608763374
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1608763374
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1608763374
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1608763374
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608763374
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1608763374
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1608763374
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1608763374
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1608763374
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1608763374
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1608763374
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608763374
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_84
timestamp 1608763374
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608763374
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1608763374
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1608763374
transform 1 0 7728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_60
timestamp 1608763374
transform 1 0 6624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_56
timestamp 1608763374
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1608763374
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 5336 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1608763374
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_44
timestamp 1608763374
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1608763374
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1608763374
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608763374
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_25
timestamp 1608763374
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1608763374
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1608763374
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1608763374
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1608763374
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608763374
transform 1 0 1564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2116 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2852 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608763374
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1608763374
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_9
timestamp 1608763374
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1608763374
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608763374
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1608763374
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1608763374
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608763374
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1608763374
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1608763374
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1608763374
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1608763374
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1608763374
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 10856 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608763374
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_105
timestamp 1608763374
transform 1 0 10764 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1608763374
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_116
timestamp 1608763374
transform 1 0 11776 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1608763374
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 9200 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1608763374
transform 1 0 9752 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_98
timestamp 1608763374
transform 1 0 10120 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1608763374
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 7728 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_66
timestamp 1608763374
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_70
timestamp 1608763374
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1608763374
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_82
timestamp 1608763374
transform 1 0 8648 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1608763374
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608763374
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1608763374
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1608763374
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1608763374
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_49
timestamp 1608763374
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_45
timestamp 1608763374
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1608763374
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1608763374
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1608763374
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_37
timestamp 1608763374
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1608763374
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_33
timestamp 1608763374
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1608763374
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_29
timestamp 1608763374
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_25
timestamp 1608763374
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1608763374
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_21
timestamp 1608763374
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608763374
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608763374
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608763374
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1608763374
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1608763374
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1608763374
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1608763374
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608763374
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608763374
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1608763374
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608763374
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1608763374
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1608763374
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1608763374
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608763374
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1608763374
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1608763374
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1608763374
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1608763374
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_132
timestamp 1608763374
transform 1 0 13248 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_144
timestamp 1608763374
transform 1 0 14352 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608763374
transform 1 0 10856 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1608763374
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_113
timestamp 1608763374
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_117
timestamp 1608763374
transform 1 0 11868 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_125
timestamp 1608763374
transform 1 0 12604 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1608763374
transform 1 0 9844 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608763374
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1608763374
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1608763374
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1608763374
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_104
timestamp 1608763374
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_79
timestamp 1608763374
transform 1 0 8372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_75
timestamp 1608763374
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1608763374
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1608763374
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1608763374
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1608763374
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1608763374
transform 1 0 6532 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1608763374
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1608763374
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1608763374
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_47
timestamp 1608763374
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_43
timestamp 1608763374
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_36
timestamp 1608763374
transform 1 0 4416 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_39
timestamp 1608763374
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608763374
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1608763374
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1608763374
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1608763374
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608763374
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2300 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608763374
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1608763374
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1608763374
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_19
timestamp 1608763374
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608763374
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608763374
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608763374
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1608763374
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608763374
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1608763374
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1608763374
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1608763374
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1608763374
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608763374
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1608763374
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1608763374
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608763374
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608763374
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1608763374
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1608763374
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1608763374
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1608763374
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_163
timestamp 1608763374
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1608763374
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1608763374
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_138
timestamp 1608763374
transform 1 0 13800 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1608763374
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 11316 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608763374
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1608763374
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_112
timestamp 1608763374
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1608763374
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608763374
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 9936 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608763374
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_87
timestamp 1608763374
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1608763374
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_88
timestamp 1608763374
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_92
timestamp 1608763374
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608763374
transform 1 0 8556 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1608763374
transform 1 0 8280 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 8096 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1608763374
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1608763374
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_74
timestamp 1608763374
transform 1 0 7912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_78
timestamp 1608763374
transform 1 0 8280 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608763374
transform 1 0 5980 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 5704 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608763374
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_48
timestamp 1608763374
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_50
timestamp 1608763374
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_56
timestamp 1608763374
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1608763374
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608763374
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608763374
transform 1 0 3036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 4232 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608763374
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_25
timestamp 1608763374
transform 1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_26
timestamp 1608763374
transform 1 0 3496 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_32
timestamp 1608763374
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2944 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1608763374
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1608763374
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608763374
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2300 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2208 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1608763374
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_10
timestamp 1608763374
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608763374
transform 1 0 1656 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608763374
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608763374
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1608763374
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1608763374
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608763374
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1608763374
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1608763374
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608763374
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_167
timestamp 1608763374
transform 1 0 16468 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1608763374
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608763374
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_155
timestamp 1608763374
transform 1 0 15364 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_126
timestamp 1608763374
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_130
timestamp 1608763374
transform 1 0 13064 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_135
timestamp 1608763374
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1608763374
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_143
timestamp 1608763374
transform 1 0 14260 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608763374
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1608763374
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608763374
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1608763374
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1608763374
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1608763374
transform 1 0 9752 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1608763374
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1608763374
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 8096 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1608763374
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_75
timestamp 1608763374
transform 1 0 8004 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1608763374
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1608763374
transform 1 0 5612 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608763374
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_45
timestamp 1608763374
transform 1 0 5244 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1608763374
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1608763374
transform 1 0 4416 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1608763374
transform 1 0 3404 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_21
timestamp 1608763374
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1608763374
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608763374
transform 1 0 1564 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2116 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608763374
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1608763374
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1608763374
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1608763374
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608763374
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608763374
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608763374
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608763374
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1608763374
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1608763374
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1608763374
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608763374
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1608763374
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1608763374
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1608763374
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1608763374
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_130
timestamp 1608763374
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1608763374
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1608763374
transform 1 0 11500 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_106
timestamp 1608763374
transform 1 0 10856 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_111
timestamp 1608763374
transform 1 0 11316 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_122
timestamp 1608763374
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608763374
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608763374
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1608763374
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1608763374
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1608763374
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1608763374
transform 1 0 8280 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_76
timestamp 1608763374
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608763374
transform 1 0 6164 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 6624 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_48
timestamp 1608763374
transform 1 0 5520 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_52
timestamp 1608763374
transform 1 0 5888 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1608763374
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608763374
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_24
timestamp 1608763374
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1608763374
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608763374
transform 1 0 1472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2760 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608763374
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608763374
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_8
timestamp 1608763374
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1608763374
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608763374
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1608763374
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1608763374
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608763374
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1608763374
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1608763374
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1608763374
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1608763374
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1608763374
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1608763374
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1608763374
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608763374
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1608763374
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_119
timestamp 1608763374
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1608763374
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_111
timestamp 1608763374
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_107
timestamp 1608763374
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 9108 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_84
timestamp 1608763374
transform 1 0 8832 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_103
timestamp 1608763374
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1608763374
transform 1 0 7176 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1608763374
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_79
timestamp 1608763374
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1608763374
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608763374
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_55
timestamp 1608763374
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_50
timestamp 1608763374
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1608763374
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_46
timestamp 1608763374
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_35
timestamp 1608763374
transform 1 0 4324 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_39
timestamp 1608763374
transform 1 0 4692 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608763374
transform 1 0 1472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 2852 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2024 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608763374
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1608763374
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_8
timestamp 1608763374
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_16
timestamp 1608763374
transform 1 0 2576 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608763374
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608763374
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1608763374
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1608763374
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1608763374
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1608763374
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1608763374
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608763374
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1608763374
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1608763374
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1608763374
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1608763374
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1608763374
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1608763374
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_140
timestamp 1608763374
transform 1 0 13984 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1608763374
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1608763374
transform 1 0 12144 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_124
timestamp 1608763374
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608763374
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 10304 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608763374
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1608763374
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1608763374
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_96
timestamp 1608763374
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 6992 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_63
timestamp 1608763374
transform 1 0 6900 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1608763374
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1608763374
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1608763374
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608763374
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 4692 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608763374
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 4508 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1608763374
transform 1 0 3312 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_28
timestamp 1608763374
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_35
timestamp 1608763374
transform 1 0 4324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608763374
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608763374
transform 1 0 2944 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2208 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608763374
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1608763374
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1608763374
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1608763374
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608763374
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1608763374
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1608763374
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608763374
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1608763374
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1608763374
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_147
timestamp 1608763374
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1608763374
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_163
timestamp 1608763374
transform 1 0 16100 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_143
timestamp 1608763374
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1608763374
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_135
timestamp 1608763374
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1608763374
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 12972 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 1608763374
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608763374
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1608763374
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1608763374
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1608763374
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1608763374
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1608763374
transform 1 0 9384 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608763374
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_85
timestamp 1608763374
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_89
timestamp 1608763374
transform 1 0 9292 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1608763374
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608763374
transform 1 0 7268 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 8280 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1608763374
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_76
timestamp 1608763374
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1608763374
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 5060 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608763374
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608763374
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1608763374
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608763374
transform 1 0 4600 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608763374
transform 1 0 3496 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_23
timestamp 1608763374
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_35
timestamp 1608763374
transform 1 0 4324 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_41
timestamp 1608763374
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608763374
transform 1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2300 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608763374
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608763374
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1608763374
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1608763374
transform 1 0 2852 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608763374
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608763374
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608763374
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608763374
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608763374
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1608763374
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1608763374
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_194
timestamp 1608763374
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1608763374
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608763374
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_167
timestamp 1608763374
transform 1 0 16468 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1608763374
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1608763374
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_170
timestamp 1608763374
transform 1 0 16744 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_182
timestamp 1608763374
transform 1 0 17848 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_158
timestamp 1608763374
transform 1 0 15640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1608763374
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1608763374
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1608763374
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1608763374
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608763374
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1608763374
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1608763374
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_147
timestamp 1608763374
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_146
timestamp 1608763374
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1608763374
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_142
timestamp 1608763374
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1608763374
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1608763374
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_135
timestamp 1608763374
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1608763374
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1608763374
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1608763374
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1608763374
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_126
timestamp 1608763374
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1608763374
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608763374
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1608763374
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_122
timestamp 1608763374
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1608763374
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_118
timestamp 1608763374
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1608763374
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_114
timestamp 1608763374
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_111
timestamp 1608763374
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1608763374
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 9844 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 9752 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608763374
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1608763374
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1608763374
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608763374
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608763374
transform 1 0 8832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608763374
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_87
timestamp 1608763374
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 7268 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608763374
transform 1 0 7820 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1608763374
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1608763374
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_64
timestamp 1608763374
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_83
timestamp 1608763374
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608763374
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608763374
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1608763374
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1608763374
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1608763374
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608763374
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 5244 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1608763374
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1608763374
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1608763374
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1608763374
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1608763374
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608763374
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608763374
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1608763374
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1608763374
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_26
timestamp 1608763374
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 2576 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608763374
transform 1 0 2392 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 2944 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1608763374
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_12
timestamp 1608763374
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1608763374
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 1656 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 1656 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608763374
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608763374
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1608763374
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1608763374
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608763374
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608763374
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1608763374
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1608763374
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1608763374
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1608763374
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1608763374
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_190
timestamp 1608763374
transform 1 0 18584 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_194
timestamp 1608763374
transform 1 0 18952 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1608763374
transform 1 0 19228 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1608763374
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1608763374
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1608763374
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_166
timestamp 1608763374
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 16192 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_162
timestamp 1608763374
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_158
timestamp 1608763374
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608763374
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1608763374
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1608763374
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1608763374
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1608763374
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1608763374
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1608763374
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1608763374
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_125
timestamp 1608763374
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1608763374
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 11960 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_114
timestamp 1608763374
transform 1 0 11592 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1608763374
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1608763374
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1608763374
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608763374
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_86
timestamp 1608763374
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1608763374
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 7176 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1608763374
transform 1 0 7084 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1608763374
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 5244 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_61
timestamp 1608763374
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608763374
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608763374
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1608763374
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1608763374
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608763374
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1608763374
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608763374
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608763374
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1608763374
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1608763374
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608763374
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_209
timestamp 1608763374
transform 1 0 20332 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1608763374
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608763374
transform 1 0 19044 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608763374
transform 1 0 19596 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1608763374
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_192
timestamp 1608763374
transform 1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1608763374
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_205
timestamp 1608763374
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608763374
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1608763374
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_184
timestamp 1608763374
transform 1 0 18032 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_167
timestamp 1608763374
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1608763374
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1608763374
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1608763374
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1608763374
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1608763374
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1608763374
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_147
timestamp 1608763374
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1608763374
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1608763374
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1608763374
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1608763374
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1608763374
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608763374
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1608763374
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1608763374
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608763374
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1608763374
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 10028 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1608763374
transform 1 0 9016 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_85
timestamp 1608763374
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1608763374
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1608763374
transform 1 0 7360 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1608763374
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1608763374
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 5060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608763374
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608763374
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1608763374
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 3312 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_40
timestamp 1608763374
transform 1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1608763374
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608763374
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1608763374
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1608763374
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1608763374
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608763374
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608763374
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1608763374
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1608763374
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608763374
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608763374
transform 1 0 18492 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_193
timestamp 1608763374
transform 1 0 18860 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1608763374
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_186
timestamp 1608763374
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_182
timestamp 1608763374
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_178
timestamp 1608763374
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1608763374
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1608763374
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1608763374
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1608763374
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_158
timestamp 1608763374
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1608763374
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608763374
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1608763374
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1608763374
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1608763374
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1608763374
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1608763374
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1608763374
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_126
timestamp 1608763374
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608763374
transform 1 0 11316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1608763374
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1608763374
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_114
timestamp 1608763374
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_118
timestamp 1608763374
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1608763374
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608763374
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1608763374
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608763374
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 7544 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1608763374
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608763374
transform 1 0 6164 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1608763374
transform 1 0 5152 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_42
timestamp 1608763374
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp 1608763374
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1608763374
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1608763374
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608763374
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_23
timestamp 1608763374
transform 1 0 3220 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1608763374
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1608763374
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_38
timestamp 1608763374
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 1748 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608763374
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1608763374
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608763374
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_217
timestamp 1608763374
transform 1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1608763374
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1608763374
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_189
timestamp 1608763374
transform 1 0 18492 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1608763374
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1608763374
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_201
timestamp 1608763374
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1608763374
transform 1 0 19964 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608763374
transform 1 0 18124 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608763374
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1608763374
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1608763374
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608763374
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp 1608763374
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1608763374
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_165
timestamp 1608763374
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1608763374
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1608763374
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1608763374
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1608763374
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1608763374
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1608763374
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1608763374
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_137
timestamp 1608763374
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_133
timestamp 1608763374
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1608763374
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608763374
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 11224 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_108
timestamp 1608763374
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1608763374
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_117
timestamp 1608763374
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1608763374
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1608763374
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1608763374
transform 1 0 10212 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_97
timestamp 1608763374
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608763374
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 8556 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1608763374
transform 1 0 7544 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_68
timestamp 1608763374
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_79
timestamp 1608763374
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608763374
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_55
timestamp 1608763374
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608763374
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1608763374
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608763374
transform 1 0 4232 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 4692 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1608763374
transform 1 0 3128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_31
timestamp 1608763374
transform 1 0 3956 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_37
timestamp 1608763374
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 1472 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608763374
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608763374
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_20
timestamp 1608763374
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608763374
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608763374
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608763374
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608763374
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1608763374
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608763374
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1608763374
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1608763374
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1608763374
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1608763374
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1608763374
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_202
timestamp 1608763374
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1608763374
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_198
timestamp 1608763374
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1608763374
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1608763374
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1608763374
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1608763374
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1608763374
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1608763374
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_186
timestamp 1608763374
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608763374
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1608763374
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1608763374
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_178
timestamp 1608763374
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1608763374
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_174
timestamp 1608763374
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1608763374
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1608763374
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1608763374
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1608763374
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1608763374
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 1608763374
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1608763374
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_159
timestamp 1608763374
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_158
timestamp 1608763374
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1608763374
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608763374
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1608763374
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1608763374
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1608763374
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 13892 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1608763374
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_136
timestamp 1608763374
transform 1 0 13616 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1608763374
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1608763374
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1608763374
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 12144 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1608763374
transform 1 0 11224 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1608763374
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608763374
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1608763374
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 10304 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1608763374
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1608763374
transform 1 0 10672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_97
timestamp 1608763374
transform 1 0 10028 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608763374
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608763374
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_89
timestamp 1608763374
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1608763374
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1608763374
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_83
timestamp 1608763374
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608763374
transform 1 0 8004 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608763374
transform 1 0 8464 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 8464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1608763374
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_79
timestamp 1608763374
transform 1 0 8372 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1608763374
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608763374
transform 1 0 7176 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1608763374
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1608763374
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 6716 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1608763374
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1608763374
transform 1 0 5612 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608763374
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1608763374
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1608763374
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1608763374
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1608763374
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1608763374
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1608763374
transform 1 0 4600 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1608763374
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608763374
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1608763374
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1608763374
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1608763374
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_25
timestamp 1608763374
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608763374
transform 1 0 3128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_22
timestamp 1608763374
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_20
timestamp 1608763374
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1608763374
transform 1 0 2300 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1608763374
transform 1 0 2116 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608763374
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608763374
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1608763374
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1608763374
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1608763374
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1608763374
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608763374
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608763374
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 20516 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1608763374
transform 1 0 20332 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1608763374
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1608763374
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608763374
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_205
timestamp 1608763374
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1608763374
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1608763374
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1608763374
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1608763374
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_185
timestamp 1608763374
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_181
timestamp 1608763374
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 1608763374
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1608763374
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_169
timestamp 1608763374
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1608763374
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608763374
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1608763374
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1608763374
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_161
timestamp 1608763374
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1608763374
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1608763374
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 11868 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1608763374
transform 1 0 11132 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_113
timestamp 1608763374
transform 1 0 11500 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1608763374
transform 1 0 11776 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608763374
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1608763374
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1608763374
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1608763374
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608763374
transform 1 0 8280 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_75
timestamp 1608763374
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608763374
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 6532 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1608763374
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_50
timestamp 1608763374
transform 1 0 5704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1608763374
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608763374
transform 1 0 4416 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608763374
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1608763374
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1608763374
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1608763374
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 1748 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608763374
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1608763374
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608763374
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608763374
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608763374
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1608763374
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1608763374
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_208
timestamp 1608763374
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1608763374
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1608763374
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1608763374
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1608763374
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1608763374
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 17112 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608763374
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1608763374
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1608763374
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1608763374
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1608763374
transform 1 0 14536 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 16376 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1608763374
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_159
timestamp 1608763374
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_163
timestamp 1608763374
transform 1 0 16100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1608763374
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_126
timestamp 1608763374
transform 1 0 12696 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1608763374
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1608763374
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1608763374
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608763374
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608763374
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 12052 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp 1608763374
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 11592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1608763374
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1608763374
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608763374
transform 1 0 9660 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1608763374
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1608763374
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_102
timestamp 1608763374
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608763374
transform 1 0 8464 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1608763374
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608763374
transform 1 0 5520 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608763374
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1608763374
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1608763374
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 3864 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1608763374
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1608763374
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608763374
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1608763374
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1608763374
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1608763374
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608763374
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608763374
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608763374
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1608763374
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1608763374
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1608763374
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608763374
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_205
timestamp 1608763374
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_201
timestamp 1608763374
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1608763374
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1608763374
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_193
timestamp 1608763374
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1608763374
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1608763374
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1608763374
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_185
timestamp 1608763374
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 15916 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608763374
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_147
timestamp 1608763374
transform 1 0 14628 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608763374
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1608763374
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1608763374
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1608763374
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1608763374
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1608763374
transform 1 0 13524 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1608763374
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608763374
transform 1 0 12512 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 10856 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1608763374
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_103
timestamp 1608763374
transform 1 0 10580 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_99
timestamp 1608763374
transform 1 0 10212 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608763374
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608763374
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1608763374
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_86
timestamp 1608763374
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_63
timestamp 1608763374
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1608763374
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1608763374
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_76
timestamp 1608763374
transform 1 0 8096 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1608763374
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 5428 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1608763374
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608763374
transform 1 0 4416 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608763374
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_22
timestamp 1608763374
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1608763374
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1608763374
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 1656 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608763374
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1608763374
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608763374
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1608763374
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_mem_bottom_track_1.prog_clk_A
timestamp 1608763374
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1608763374
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1608763374
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1608763374
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1608763374
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1608763374
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1608763374
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1608763374
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_192
timestamp 1608763374
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1608763374
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1608763374
transform 1 0 17296 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608763374
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1608763374
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1608763374
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1608763374
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608763374
transform 1 0 16284 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_158
timestamp 1608763374
transform 1 0 15640 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_162
timestamp 1608763374
transform 1 0 16008 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 14168 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1608763374
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1608763374
transform 1 0 13616 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1608763374
transform 1 0 10948 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1608763374
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608763374
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1608763374
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1608763374
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608763374
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 9292 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1608763374
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 7636 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_68
timestamp 1608763374
transform 1 0 7360 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608763374
transform 1 0 5060 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608763374
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_52
timestamp 1608763374
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_56
timestamp 1608763374
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1608763374
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1608763374
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608763374
transform 1 0 4048 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608763374
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_30
timestamp 1608763374
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_41
timestamp 1608763374
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608763374
transform 1 0 2024 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608763374
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1608763374
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1608763374
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1608763374
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608763374
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608763374
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1608763374
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1608763374
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608763374
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1608763374
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1608763374
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_202
timestamp 1608763374
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1608763374
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1608763374
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1608763374
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1608763374
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1608763374
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1608763374
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 16008 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608763374
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1608763374
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_160
timestamp 1608763374
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 13432 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1608763374
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_132
timestamp 1608763374
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 11316 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_105
timestamp 1608763374
transform 1 0 10764 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608763374
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608763374
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608763374
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_96
timestamp 1608763374
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_100
timestamp 1608763374
transform 1 0 10304 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1608763374
transform 1 0 7176 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1608763374
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp 1608763374
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1608763374
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 5980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1608763374
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp 1608763374
transform 1 0 5704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1608763374
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp 1608763374
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608763374
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608763374
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1608763374
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1608763374
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1608763374
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1608763374
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 1380 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608763374
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1608763374
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608763374
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608763374
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1608763374
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608763374
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608763374
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1608763374
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1608763374
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_216
timestamp 1608763374
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1608763374
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_212
timestamp 1608763374
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1608763374
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1608763374
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_205
timestamp 1608763374
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1608763374
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1608763374
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_200
timestamp 1608763374
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1608763374
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_196
timestamp 1608763374
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1608763374
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1608763374
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1608763374
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1608763374
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 16652 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608763374
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_185
timestamp 1608763374
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1608763374
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1608763374
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1608763374
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_173
timestamp 1608763374
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_177
timestamp 1608763374
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608763374
transform 1 0 16192 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608763374
transform 1 0 15456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_159
timestamp 1608763374
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1608763374
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1608763374
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608763374
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608763374
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 1608763374
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1608763374
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_150
timestamp 1608763374
transform 1 0 14904 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1608763374
transform 1 0 14076 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1608763374
transform 1 0 14076 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 13340 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_127
timestamp 1608763374
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_131
timestamp 1608763374
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_139
timestamp 1608763374
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1608763374
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608763374
transform 1 0 11960 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608763374
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1608763374
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_117
timestamp 1608763374
transform 1 0 11868 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_116
timestamp 1608763374
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1608763374
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 10304 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608763374
transform 1 0 10672 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1608763374
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_94
timestamp 1608763374
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1608763374
transform 1 0 10212 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608763374
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608763374
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1608763374
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 1608763374
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608763374
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 7176 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 8280 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1608763374
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_82
timestamp 1608763374
transform 1 0 8648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1608763374
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp 1608763374
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 5520 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608763374
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1608763374
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608763374
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_53
timestamp 1608763374
transform 1 0 5980 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608763374
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_45
timestamp 1608763374
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_49
timestamp 1608763374
transform 1 0 5612 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 4140 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608763374
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1608763374
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608763374
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1608763374
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1608763374
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_28
timestamp 1608763374
transform 1 0 3680 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 2208 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608763374
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_10
timestamp 1608763374
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_10
timestamp 1608763374
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608763374
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1608763374
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608763374
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608763374
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1608763374
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1608763374
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608763374
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1608763374
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_212
timestamp 1608763374
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1608763374
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp 1608763374
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1608763374
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_204
timestamp 1608763374
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1608763374
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1608763374
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1608763374
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_192
timestamp 1608763374
transform 1 0 18768 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1608763374
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608763374
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 17664 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1608763374
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1608763374
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1608763374
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608763374
transform 1 0 14720 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 16008 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1608763374
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 1608763374
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1608763374
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_159
timestamp 1608763374
transform 1 0 15732 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 13984 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_126
timestamp 1608763374
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_130
timestamp 1608763374
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_134
timestamp 1608763374
transform 1 0 13432 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608763374
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608763374
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608763374
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1608763374
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1608763374
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 9476 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_84
timestamp 1608763374
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_88
timestamp 1608763374
transform 1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1608763374
transform 1 0 6992 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1608763374
transform 1 0 8004 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1608763374
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1608763374
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608763374
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608763374
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_42
timestamp 1608763374
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1608763374
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608763374
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1608763374
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608763374
transform 1 0 3772 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1608763374
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp 1608763374
transform 1 0 3312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp 1608763374
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608763374
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1608763374
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1608763374
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_9
timestamp 1608763374
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1608763374
transform 1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_17
timestamp 1608763374
transform 1 0 2668 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_20
timestamp 1608763374
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608763374
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608763374
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1608763374
transform 1 0 21068 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1608763374
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1608763374
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608763374
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1608763374
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1608763374
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608763374
transform 1 0 17940 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1608763374
transform 1 0 16928 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_170
timestamp 1608763374
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_181
timestamp 1608763374
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1608763374
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 15272 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608763374
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_147
timestamp 1608763374
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608763374
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608763374
transform 1 0 13984 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1608763374
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1608763374
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 12328 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1608763374
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608763374
transform 1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 10672 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608763374
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1608763374
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1608763374
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1608763374
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1608763374
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1608763374
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1608763374
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1608763374
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1608763374
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1608763374
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1608763374
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608763374
transform 1 0 5336 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608763374
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1608763374
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_42
timestamp 1608763374
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_55
timestamp 1608763374
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608763374
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1608763374
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1608763374
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1608763374
transform 1 0 4416 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608763374
transform 1 0 1748 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608763374
transform 1 0 2760 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608763374
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1608763374
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_16
timestamp 1608763374
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608763374
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1608763374
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1608763374
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1608763374
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1608763374
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1608763374
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1608763374
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1608763374
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_205
timestamp 1608763374
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp 1608763374
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_196
timestamp 1608763374
transform 1 0 19136 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1608763374
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1608763374
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608763374
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_174
timestamp 1608763374
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1608763374
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1608763374
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1608763374
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 14628 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1608763374
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1608763374
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 12972 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1608763374
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1608763374
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1608763374
transform 1 0 11224 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608763374
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1608763374
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_107
timestamp 1608763374
transform 1 0 10948 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1608763374
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1608763374
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608763374
transform 1 0 9752 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1608763374
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1608763374
transform 1 0 10580 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608763374
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1608763374
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_82
timestamp 1608763374
transform 1 0 8648 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608763374
transform 1 0 5244 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608763374
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1608763374
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1608763374
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1608763374
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1608763374
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 3588 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1608763374
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1608763374
transform 1 0 1472 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 1932 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608763374
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608763374
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1608763374
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608763374
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608763374
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608763374
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1608763374
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1608763374
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1608763374
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1608763374
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1608763374
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_207
timestamp 1608763374
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1608763374
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1608763374
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1608763374
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_195
timestamp 1608763374
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_191
timestamp 1608763374
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 16652 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 17756 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 18124 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_175
timestamp 1608763374
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_179
timestamp 1608763374
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp 1608763374
transform 1 0 17940 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1608763374
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608763374
transform 1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608763374
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1608763374
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1608763374
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_165
timestamp 1608763374
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1608763374
transform 1 0 12972 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1608763374
transform 1 0 13984 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_126
timestamp 1608763374
transform 1 0 12696 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1608763374
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 12144 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1608763374
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1608763374
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_113
timestamp 1608763374
transform 1 0 11500 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1608763374
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608763374
transform 1 0 9936 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608763374
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608763374
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1608763374
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 7912 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1608763374
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1608763374
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_67
timestamp 1608763374
transform 1 0 7268 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1608763374
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763374
transform 1 0 5428 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608763374
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 3220 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608763374
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1608763374
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1608763374
transform 1 0 4876 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 1472 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608763374
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1608763374
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_20
timestamp 1608763374
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608763374
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608763374
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1608763374
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608763374
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1608763374
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1608763374
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608763374
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_215
timestamp 1608763374
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608763374
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1608763374
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608763374
transform 1 0 19780 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608763374
transform 1 0 19964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608763374
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1608763374
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_198
timestamp 1608763374
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_202
timestamp 1608763374
transform 1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608763374
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608763374
transform 1 0 18584 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1608763374
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1608763374
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1608763374
transform 1 0 19228 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1608763374
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_194
timestamp 1608763374
transform 1 0 18952 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608763374
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608763374
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608763374
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608763374
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608763374
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608763374
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608763374
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 17112 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1608763374
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_180
timestamp 1608763374
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608763374
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1608763374
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1608763374
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 16376 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1608763374
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608763374
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608763374
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1608763374
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_164
timestamp 1608763374
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608763374
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 14536 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1608763374
transform 1 0 15364 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608763374
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1608763374
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608763374
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp 1608763374
transform 1 0 15088 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608763374
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1608763374
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1608763374
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_141
timestamp 1608763374
transform 1 0 14076 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608763374
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1608763374
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_137
timestamp 1608763374
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608763374
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 13156 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1608763374
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1608763374
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608763374
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608763374
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608763374
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1608763374
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1608763374
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608763374
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763374
transform 1 0 11500 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115
timestamp 1608763374
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1608763374
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_111
timestamp 1608763374
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_111
timestamp 1608763374
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608763374
transform 1 0 10488 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608763374
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608763374
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608763374
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1608763374
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_99
timestamp 1608763374
transform 1 0 10212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 8740 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608763374
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1608763374
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1608763374
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1608763374
transform 1 0 8280 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1608763374
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1608763374
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1608763374
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608763374
transform 1 0 6992 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608763374
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1608763374
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608763374
transform 1 0 6164 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608763374
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608763374
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608763374
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48
timestamp 1608763374
transform 1 0 5520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1608763374
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1608763374
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1608763374
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1608763374
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763374
transform 1 0 4048 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763374
transform 1 0 4508 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608763374
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1608763374
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608763374
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28
timestamp 1608763374
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_28
timestamp 1608763374
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_32
timestamp 1608763374
transform 1 0 4048 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608763374
transform 1 0 2852 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608763374
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1608763374
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1608763374
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1608763374
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1608763374
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1608763374
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1608763374
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1608763374
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1608763374
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1608763374
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1608763374
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608763374
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1608763374
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1608763374
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7
timestamp 1608763374
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608763374
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608763374
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1608763374
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1608763374
transform 1 0 1380 0 1 2720
box -38 -48 222 592
<< labels >>
rlabel metal2 s 21638 0 21694 800 4 SC_IN_BOT
port 1 nsew
rlabel metal2 s 22098 0 22154 800 4 SC_OUT_BOT
port 2 nsew
rlabel metal2 s 202 0 258 800 4 bottom_left_grid_pin_42_
port 3 nsew
rlabel metal2 s 570 0 626 800 4 bottom_left_grid_pin_43_
port 4 nsew
rlabel metal2 s 1030 0 1086 800 4 bottom_left_grid_pin_44_
port 5 nsew
rlabel metal2 s 1490 0 1546 800 4 bottom_left_grid_pin_45_
port 6 nsew
rlabel metal2 s 1950 0 2006 800 4 bottom_left_grid_pin_46_
port 7 nsew
rlabel metal2 s 2318 0 2374 800 4 bottom_left_grid_pin_47_
port 8 nsew
rlabel metal2 s 2778 0 2834 800 4 bottom_left_grid_pin_48_
port 9 nsew
rlabel metal2 s 3238 0 3294 800 4 bottom_left_grid_pin_49_
port 10 nsew
rlabel metal2 s 21178 0 21234 800 4 bottom_right_grid_pin_1_
port 11 nsew
rlabel metal3 s 22000 5720 22800 5840 4 ccff_head
port 12 nsew
rlabel metal3 s 22000 17144 22800 17264 4 ccff_tail
port 13 nsew
rlabel metal3 s 0 3816 800 3936 4 chanx_left_in[0]
port 14 nsew
rlabel metal3 s 0 8440 800 8560 4 chanx_left_in[10]
port 15 nsew
rlabel metal3 s 0 8984 800 9104 4 chanx_left_in[11]
port 16 nsew
rlabel metal3 s 0 9392 800 9512 4 chanx_left_in[12]
port 17 nsew
rlabel metal3 s 0 9936 800 10056 4 chanx_left_in[13]
port 18 nsew
rlabel metal3 s 0 10344 800 10464 4 chanx_left_in[14]
port 19 nsew
rlabel metal3 s 0 10752 800 10872 4 chanx_left_in[15]
port 20 nsew
rlabel metal3 s 0 11296 800 11416 4 chanx_left_in[16]
port 21 nsew
rlabel metal3 s 0 11704 800 11824 4 chanx_left_in[17]
port 22 nsew
rlabel metal3 s 0 12248 800 12368 4 chanx_left_in[18]
port 23 nsew
rlabel metal3 s 0 12656 800 12776 4 chanx_left_in[19]
port 24 nsew
rlabel metal3 s 0 4224 800 4344 4 chanx_left_in[1]
port 25 nsew
rlabel metal3 s 0 4768 800 4888 4 chanx_left_in[2]
port 26 nsew
rlabel metal3 s 0 5176 800 5296 4 chanx_left_in[3]
port 27 nsew
rlabel metal3 s 0 5720 800 5840 4 chanx_left_in[4]
port 28 nsew
rlabel metal3 s 0 6128 800 6248 4 chanx_left_in[5]
port 29 nsew
rlabel metal3 s 0 6672 800 6792 4 chanx_left_in[6]
port 30 nsew
rlabel metal3 s 0 7080 800 7200 4 chanx_left_in[7]
port 31 nsew
rlabel metal3 s 0 7488 800 7608 4 chanx_left_in[8]
port 32 nsew
rlabel metal3 s 0 8032 800 8152 4 chanx_left_in[9]
port 33 nsew
rlabel metal3 s 0 13200 800 13320 4 chanx_left_out[0]
port 34 nsew
rlabel metal3 s 0 17824 800 17944 4 chanx_left_out[10]
port 35 nsew
rlabel metal3 s 0 18232 800 18352 4 chanx_left_out[11]
port 36 nsew
rlabel metal3 s 0 18776 800 18896 4 chanx_left_out[12]
port 37 nsew
rlabel metal3 s 0 19184 800 19304 4 chanx_left_out[13]
port 38 nsew
rlabel metal3 s 0 19728 800 19848 4 chanx_left_out[14]
port 39 nsew
rlabel metal3 s 0 20136 800 20256 4 chanx_left_out[15]
port 40 nsew
rlabel metal3 s 0 20544 800 20664 4 chanx_left_out[16]
port 41 nsew
rlabel metal3 s 0 21088 800 21208 4 chanx_left_out[17]
port 42 nsew
rlabel metal3 s 0 21496 800 21616 4 chanx_left_out[18]
port 43 nsew
rlabel metal3 s 0 22040 800 22160 4 chanx_left_out[19]
port 44 nsew
rlabel metal3 s 0 13608 800 13728 4 chanx_left_out[1]
port 45 nsew
rlabel metal3 s 0 14016 800 14136 4 chanx_left_out[2]
port 46 nsew
rlabel metal3 s 0 14560 800 14680 4 chanx_left_out[3]
port 47 nsew
rlabel metal3 s 0 14968 800 15088 4 chanx_left_out[4]
port 48 nsew
rlabel metal3 s 0 15512 800 15632 4 chanx_left_out[5]
port 49 nsew
rlabel metal3 s 0 15920 800 16040 4 chanx_left_out[6]
port 50 nsew
rlabel metal3 s 0 16464 800 16584 4 chanx_left_out[7]
port 51 nsew
rlabel metal3 s 0 16872 800 16992 4 chanx_left_out[8]
port 52 nsew
rlabel metal3 s 0 17280 800 17400 4 chanx_left_out[9]
port 53 nsew
rlabel metal2 s 3698 0 3754 800 4 chany_bottom_in[0]
port 54 nsew
rlabel metal2 s 8022 0 8078 800 4 chany_bottom_in[10]
port 55 nsew
rlabel metal2 s 8482 0 8538 800 4 chany_bottom_in[11]
port 56 nsew
rlabel metal2 s 8942 0 8998 800 4 chany_bottom_in[12]
port 57 nsew
rlabel metal2 s 9402 0 9458 800 4 chany_bottom_in[13]
port 58 nsew
rlabel metal2 s 9770 0 9826 800 4 chany_bottom_in[14]
port 59 nsew
rlabel metal2 s 10230 0 10286 800 4 chany_bottom_in[15]
port 60 nsew
rlabel metal2 s 10690 0 10746 800 4 chany_bottom_in[16]
port 61 nsew
rlabel metal2 s 11150 0 11206 800 4 chany_bottom_in[17]
port 62 nsew
rlabel metal2 s 11610 0 11666 800 4 chany_bottom_in[18]
port 63 nsew
rlabel metal2 s 11978 0 12034 800 4 chany_bottom_in[19]
port 64 nsew
rlabel metal2 s 4066 0 4122 800 4 chany_bottom_in[1]
port 65 nsew
rlabel metal2 s 4526 0 4582 800 4 chany_bottom_in[2]
port 66 nsew
rlabel metal2 s 4986 0 5042 800 4 chany_bottom_in[3]
port 67 nsew
rlabel metal2 s 5446 0 5502 800 4 chany_bottom_in[4]
port 68 nsew
rlabel metal2 s 5906 0 5962 800 4 chany_bottom_in[5]
port 69 nsew
rlabel metal2 s 6274 0 6330 800 4 chany_bottom_in[6]
port 70 nsew
rlabel metal2 s 6734 0 6790 800 4 chany_bottom_in[7]
port 71 nsew
rlabel metal2 s 7194 0 7250 800 4 chany_bottom_in[8]
port 72 nsew
rlabel metal2 s 7654 0 7710 800 4 chany_bottom_in[9]
port 73 nsew
rlabel metal2 s 12438 0 12494 800 4 chany_bottom_out[0]
port 74 nsew
rlabel metal2 s 16854 0 16910 800 4 chany_bottom_out[10]
port 75 nsew
rlabel metal2 s 17314 0 17370 800 4 chany_bottom_out[11]
port 76 nsew
rlabel metal2 s 17682 0 17738 800 4 chany_bottom_out[12]
port 77 nsew
rlabel metal2 s 18142 0 18198 800 4 chany_bottom_out[13]
port 78 nsew
rlabel metal2 s 18602 0 18658 800 4 chany_bottom_out[14]
port 79 nsew
rlabel metal2 s 19062 0 19118 800 4 chany_bottom_out[15]
port 80 nsew
rlabel metal2 s 19430 0 19486 800 4 chany_bottom_out[16]
port 81 nsew
rlabel metal2 s 19890 0 19946 800 4 chany_bottom_out[17]
port 82 nsew
rlabel metal2 s 20350 0 20406 800 4 chany_bottom_out[18]
port 83 nsew
rlabel metal2 s 20810 0 20866 800 4 chany_bottom_out[19]
port 84 nsew
rlabel metal2 s 12898 0 12954 800 4 chany_bottom_out[1]
port 85 nsew
rlabel metal2 s 13358 0 13414 800 4 chany_bottom_out[2]
port 86 nsew
rlabel metal2 s 13726 0 13782 800 4 chany_bottom_out[3]
port 87 nsew
rlabel metal2 s 14186 0 14242 800 4 chany_bottom_out[4]
port 88 nsew
rlabel metal2 s 14646 0 14702 800 4 chany_bottom_out[5]
port 89 nsew
rlabel metal2 s 15106 0 15162 800 4 chany_bottom_out[6]
port 90 nsew
rlabel metal2 s 15474 0 15530 800 4 chany_bottom_out[7]
port 91 nsew
rlabel metal2 s 15934 0 15990 800 4 chany_bottom_out[8]
port 92 nsew
rlabel metal2 s 16394 0 16450 800 4 chany_bottom_out[9]
port 93 nsew
rlabel metal3 s 0 144 800 264 4 left_bottom_grid_pin_34_
port 94 nsew
rlabel metal3 s 0 552 800 672 4 left_bottom_grid_pin_35_
port 95 nsew
rlabel metal3 s 0 960 800 1080 4 left_bottom_grid_pin_36_
port 96 nsew
rlabel metal3 s 0 1504 800 1624 4 left_bottom_grid_pin_37_
port 97 nsew
rlabel metal3 s 0 1912 800 2032 4 left_bottom_grid_pin_38_
port 98 nsew
rlabel metal3 s 0 2456 800 2576 4 left_bottom_grid_pin_39_
port 99 nsew
rlabel metal3 s 0 2864 800 2984 4 left_bottom_grid_pin_40_
port 100 nsew
rlabel metal3 s 0 3408 800 3528 4 left_bottom_grid_pin_41_
port 101 nsew
rlabel metal3 s 0 22448 800 22568 4 left_top_grid_pin_1_
port 102 nsew
rlabel metal2 s 22558 0 22614 800 4 prog_clk_0_S_in
port 103 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 104 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 105 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22568
string GDS_FILE /ef/openfpga/openlane/runs/sb_2__2_/results/magic/sb_2__2_.gds
string GDS_END 1445034
string GDS_START 81916
<< end >>
