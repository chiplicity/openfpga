magic
tech sky130A
magscale 1 2
timestamp 1605112181
<< locali >>
rect 9321 18819 9355 18921
rect 11805 17731 11839 17833
rect 20821 11679 20855 11781
rect 18797 10999 18831 11305
rect 11989 8415 12023 8517
rect 12541 5015 12575 5117
<< viali >>
rect 16405 25449 16439 25483
rect 20177 25449 20211 25483
rect 23029 25449 23063 25483
rect 16221 25313 16255 25347
rect 18889 25313 18923 25347
rect 19993 25313 20027 25347
rect 21741 25313 21775 25347
rect 22845 25313 22879 25347
rect 24593 25313 24627 25347
rect 19073 25177 19107 25211
rect 21925 25177 21959 25211
rect 24777 25109 24811 25143
rect 16957 24769 16991 24803
rect 12541 24701 12575 24735
rect 13645 24701 13679 24735
rect 14197 24701 14231 24735
rect 14749 24701 14783 24735
rect 15301 24701 15335 24735
rect 15853 24701 15887 24735
rect 18061 24701 18095 24735
rect 19349 24701 19383 24735
rect 19533 24701 19567 24735
rect 20821 24701 20855 24735
rect 20913 24701 20947 24735
rect 22017 24701 22051 24735
rect 24593 24701 24627 24735
rect 25145 24701 25179 24735
rect 21833 24633 21867 24667
rect 12725 24565 12759 24599
rect 13093 24565 13127 24599
rect 13829 24565 13863 24599
rect 14933 24565 14967 24599
rect 16037 24565 16071 24599
rect 16405 24565 16439 24599
rect 16773 24565 16807 24599
rect 17785 24565 17819 24599
rect 18245 24565 18279 24599
rect 18889 24565 18923 24599
rect 19717 24565 19751 24599
rect 20177 24565 20211 24599
rect 21097 24565 21131 24599
rect 22201 24565 22235 24599
rect 22845 24565 22879 24599
rect 24409 24565 24443 24599
rect 24777 24565 24811 24599
rect 15853 24361 15887 24395
rect 17141 24361 17175 24395
rect 18245 24361 18279 24395
rect 19441 24361 19475 24395
rect 21189 24361 21223 24395
rect 22569 24361 22603 24395
rect 23673 24361 23707 24395
rect 13185 24225 13219 24259
rect 15761 24225 15795 24259
rect 16957 24225 16991 24259
rect 18061 24225 18095 24259
rect 19257 24225 19291 24259
rect 21005 24225 21039 24259
rect 22385 24225 22419 24259
rect 23489 24225 23523 24259
rect 24593 24225 24627 24259
rect 13277 24157 13311 24191
rect 13369 24157 13403 24191
rect 16037 24157 16071 24191
rect 10885 24021 10919 24055
rect 12449 24021 12483 24055
rect 12817 24021 12851 24055
rect 14933 24021 14967 24055
rect 15393 24021 15427 24055
rect 22109 24021 22143 24055
rect 24777 24021 24811 24055
rect 10793 23817 10827 23851
rect 14749 23817 14783 23851
rect 16313 23817 16347 23851
rect 21557 23817 21591 23851
rect 22661 23817 22695 23851
rect 23489 23817 23523 23851
rect 11345 23681 11379 23715
rect 14933 23681 14967 23715
rect 22385 23681 22419 23715
rect 23949 23681 23983 23715
rect 11161 23613 11195 23647
rect 12449 23613 12483 23647
rect 12716 23613 12750 23647
rect 17509 23613 17543 23647
rect 18061 23613 18095 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 22477 23613 22511 23647
rect 23765 23613 23799 23647
rect 25053 23613 25087 23647
rect 25605 23613 25639 23647
rect 11897 23545 11931 23579
rect 15200 23545 15234 23579
rect 18306 23545 18340 23579
rect 21097 23545 21131 23579
rect 10701 23477 10735 23511
rect 11253 23477 11287 23511
rect 12265 23477 12299 23511
rect 13829 23477 13863 23511
rect 16957 23477 16991 23511
rect 17785 23477 17819 23511
rect 19441 23477 19475 23511
rect 20085 23477 20119 23511
rect 23121 23477 23155 23511
rect 24685 23477 24719 23511
rect 25237 23477 25271 23511
rect 10885 23273 10919 23307
rect 12541 23273 12575 23307
rect 13461 23273 13495 23307
rect 15577 23273 15611 23307
rect 15945 23273 15979 23307
rect 18981 23273 19015 23307
rect 21097 23273 21131 23307
rect 11406 23205 11440 23239
rect 14105 23205 14139 23239
rect 16374 23205 16408 23239
rect 23121 23205 23155 23239
rect 24409 23205 24443 23239
rect 14013 23137 14047 23171
rect 16129 23137 16163 23171
rect 20913 23137 20947 23171
rect 22845 23137 22879 23171
rect 24133 23137 24167 23171
rect 11161 23069 11195 23103
rect 14197 23069 14231 23103
rect 14933 23069 14967 23103
rect 19073 23069 19107 23103
rect 19165 23069 19199 23103
rect 25421 23069 25455 23103
rect 13185 22933 13219 22967
rect 13645 22933 13679 22967
rect 17509 22933 17543 22967
rect 18061 22933 18095 22967
rect 18613 22933 18647 22967
rect 19717 22933 19751 22967
rect 23765 22933 23799 22967
rect 12817 22729 12851 22763
rect 13277 22729 13311 22763
rect 14749 22729 14783 22763
rect 15945 22729 15979 22763
rect 18245 22729 18279 22763
rect 21557 22729 21591 22763
rect 23397 22729 23431 22763
rect 17417 22661 17451 22695
rect 25237 22661 25271 22695
rect 11621 22593 11655 22627
rect 13369 22593 13403 22627
rect 16865 22593 16899 22627
rect 17049 22593 17083 22627
rect 17785 22593 17819 22627
rect 18797 22593 18831 22627
rect 24041 22593 24075 22627
rect 16313 22525 16347 22559
rect 16773 22525 16807 22559
rect 21373 22525 21407 22559
rect 21925 22525 21959 22559
rect 22477 22525 22511 22559
rect 23765 22525 23799 22559
rect 24501 22525 24535 22559
rect 25053 22525 25087 22559
rect 25605 22525 25639 22559
rect 13614 22457 13648 22491
rect 15301 22457 15335 22491
rect 19064 22457 19098 22491
rect 11161 22389 11195 22423
rect 16405 22389 16439 22423
rect 18613 22389 18647 22423
rect 20177 22389 20211 22423
rect 21005 22389 21039 22423
rect 22661 22389 22695 22423
rect 23121 22389 23155 22423
rect 24869 22389 24903 22423
rect 12449 22185 12483 22219
rect 13001 22185 13035 22219
rect 15117 22185 15151 22219
rect 16497 22185 16531 22219
rect 17969 22185 18003 22219
rect 18889 22185 18923 22219
rect 22753 22185 22787 22219
rect 13921 22117 13955 22151
rect 16589 22117 16623 22151
rect 20545 22117 20579 22151
rect 11069 22049 11103 22083
rect 11336 22049 11370 22083
rect 15301 22049 15335 22083
rect 17509 22049 17543 22083
rect 19165 22049 19199 22083
rect 19441 22049 19475 22083
rect 21281 22049 21315 22083
rect 24593 22049 24627 22083
rect 14013 21981 14047 22015
rect 14105 21981 14139 22015
rect 15577 21981 15611 22015
rect 18061 21981 18095 22015
rect 18153 21981 18187 22015
rect 22845 21981 22879 22015
rect 23029 21981 23063 22015
rect 13553 21913 13587 21947
rect 17601 21913 17635 21947
rect 21465 21913 21499 21947
rect 9321 21845 9355 21879
rect 10885 21845 10919 21879
rect 13461 21845 13495 21879
rect 14657 21845 14691 21879
rect 16037 21845 16071 21879
rect 17141 21845 17175 21879
rect 22017 21845 22051 21879
rect 22385 21845 22419 21879
rect 24777 21845 24811 21879
rect 9045 21641 9079 21675
rect 11805 21641 11839 21675
rect 12173 21641 12207 21675
rect 13369 21641 13403 21675
rect 14289 21641 14323 21675
rect 14473 21641 14507 21675
rect 15485 21641 15519 21675
rect 17049 21641 17083 21675
rect 18061 21641 18095 21675
rect 19441 21641 19475 21675
rect 22845 21641 22879 21675
rect 23213 21641 23247 21675
rect 25053 21641 25087 21675
rect 9873 21505 9907 21539
rect 10701 21505 10735 21539
rect 11345 21505 11379 21539
rect 13461 21505 13495 21539
rect 14933 21505 14967 21539
rect 15025 21505 15059 21539
rect 16497 21505 16531 21539
rect 16589 21505 16623 21539
rect 18613 21505 18647 21539
rect 19073 21505 19107 21539
rect 9597 21437 9631 21471
rect 16405 21437 16439 21471
rect 20545 21437 20579 21471
rect 24317 21437 24351 21471
rect 10333 21369 10367 21403
rect 11161 21369 11195 21403
rect 15945 21369 15979 21403
rect 17785 21369 17819 21403
rect 18521 21369 18555 21403
rect 20790 21369 20824 21403
rect 24593 21369 24627 21403
rect 9229 21301 9263 21335
rect 9689 21301 9723 21335
rect 10793 21301 10827 21335
rect 11253 21301 11287 21335
rect 12449 21301 12483 21335
rect 14013 21301 14047 21335
rect 14841 21301 14875 21335
rect 16037 21301 16071 21335
rect 17417 21301 17451 21335
rect 18429 21301 18463 21335
rect 19809 21301 19843 21335
rect 20453 21301 20487 21335
rect 21925 21301 21959 21335
rect 22477 21301 22511 21335
rect 24133 21301 24167 21335
rect 25605 21301 25639 21335
rect 12541 21097 12575 21131
rect 13553 21097 13587 21131
rect 17233 21097 17267 21131
rect 17693 21097 17727 21131
rect 19901 21097 19935 21131
rect 21833 21097 21867 21131
rect 13921 21029 13955 21063
rect 15546 21029 15580 21063
rect 22284 21029 22318 21063
rect 24777 21029 24811 21063
rect 10313 20961 10347 20995
rect 12449 20961 12483 20995
rect 12909 20961 12943 20995
rect 15301 20961 15335 20995
rect 18153 20961 18187 20995
rect 19533 20961 19567 20995
rect 19717 20961 19751 20995
rect 20361 20961 20395 20995
rect 20913 20961 20947 20995
rect 21465 20961 21499 20995
rect 22017 20961 22051 20995
rect 24501 20961 24535 20995
rect 10057 20893 10091 20927
rect 13001 20893 13035 20927
rect 13093 20893 13127 20927
rect 18245 20893 18279 20927
rect 18337 20893 18371 20927
rect 11437 20825 11471 20859
rect 23949 20825 23983 20859
rect 7665 20757 7699 20791
rect 9321 20757 9355 20791
rect 14565 20757 14599 20791
rect 16681 20757 16715 20791
rect 17785 20757 17819 20791
rect 18797 20757 18831 20791
rect 19165 20757 19199 20791
rect 19349 20757 19383 20791
rect 21097 20757 21131 20791
rect 23397 20757 23431 20791
rect 9597 20553 9631 20587
rect 10793 20553 10827 20587
rect 11805 20553 11839 20587
rect 12173 20553 12207 20587
rect 15301 20553 15335 20587
rect 15853 20553 15887 20587
rect 17509 20553 17543 20587
rect 23029 20553 23063 20587
rect 16405 20485 16439 20519
rect 11437 20417 11471 20451
rect 12725 20417 12759 20451
rect 13921 20417 13955 20451
rect 16865 20417 16899 20451
rect 16957 20417 16991 20451
rect 21557 20417 21591 20451
rect 22661 20417 22695 20451
rect 23673 20417 23707 20451
rect 7573 20349 7607 20383
rect 12449 20349 12483 20383
rect 18061 20349 18095 20383
rect 19533 20349 19567 20383
rect 7481 20281 7515 20315
rect 7840 20281 7874 20315
rect 10333 20281 10367 20315
rect 11161 20281 11195 20315
rect 13829 20281 13863 20315
rect 14177 20281 14211 20315
rect 16221 20281 16255 20315
rect 16773 20281 16807 20315
rect 18337 20281 18371 20315
rect 19441 20281 19475 20315
rect 19800 20281 19834 20315
rect 21833 20281 21867 20315
rect 22477 20281 22511 20315
rect 23397 20281 23431 20315
rect 23918 20281 23952 20315
rect 8953 20213 8987 20247
rect 9965 20213 9999 20247
rect 10701 20213 10735 20247
rect 11253 20213 11287 20247
rect 13277 20213 13311 20247
rect 17785 20213 17819 20247
rect 18797 20213 18831 20247
rect 20913 20213 20947 20247
rect 22017 20213 22051 20247
rect 22385 20213 22419 20247
rect 25053 20213 25087 20247
rect 7849 20009 7883 20043
rect 11069 20009 11103 20043
rect 12725 20009 12759 20043
rect 13921 20009 13955 20043
rect 15025 20009 15059 20043
rect 15761 20009 15795 20043
rect 17233 20009 17267 20043
rect 18337 20009 18371 20043
rect 20637 20009 20671 20043
rect 22845 20009 22879 20043
rect 23949 20009 23983 20043
rect 24317 20009 24351 20043
rect 18797 19941 18831 19975
rect 21189 19941 21223 19975
rect 22109 19941 22143 19975
rect 7757 19873 7791 19907
rect 9689 19873 9723 19907
rect 9956 19873 9990 19907
rect 12173 19873 12207 19907
rect 14105 19873 14139 19907
rect 16109 19873 16143 19907
rect 18521 19873 18555 19907
rect 19625 19873 19659 19907
rect 20269 19873 20303 19907
rect 20913 19873 20947 19907
rect 22753 19873 22787 19907
rect 24409 19873 24443 19907
rect 8033 19805 8067 19839
rect 12817 19805 12851 19839
rect 12909 19805 12943 19839
rect 14749 19805 14783 19839
rect 15853 19805 15887 19839
rect 19717 19805 19751 19839
rect 19901 19805 19935 19839
rect 22937 19805 22971 19839
rect 24593 19805 24627 19839
rect 19257 19737 19291 19771
rect 21649 19737 21683 19771
rect 22385 19737 22419 19771
rect 24961 19737 24995 19771
rect 7389 19669 7423 19703
rect 12357 19669 12391 19703
rect 13369 19669 13403 19703
rect 13829 19669 13863 19703
rect 18153 19669 18187 19703
rect 23673 19669 23707 19703
rect 7481 19465 7515 19499
rect 9965 19465 9999 19499
rect 11897 19465 11931 19499
rect 16405 19465 16439 19499
rect 19717 19465 19751 19499
rect 22477 19465 22511 19499
rect 24685 19465 24719 19499
rect 7113 19329 7147 19363
rect 11437 19329 11471 19363
rect 16957 19329 16991 19363
rect 17417 19329 17451 19363
rect 18613 19329 18647 19363
rect 20269 19329 20303 19363
rect 21833 19329 21867 19363
rect 24317 19329 24351 19363
rect 8033 19261 8067 19295
rect 8289 19261 8323 19295
rect 12265 19261 12299 19295
rect 12817 19261 12851 19295
rect 13084 19261 13118 19295
rect 15945 19261 15979 19295
rect 16773 19261 16807 19295
rect 17877 19261 17911 19295
rect 18429 19261 18463 19295
rect 21189 19261 21223 19295
rect 21741 19261 21775 19295
rect 23121 19261 23155 19295
rect 25053 19261 25087 19295
rect 25237 19261 25271 19295
rect 25973 19261 26007 19295
rect 7849 19193 7883 19227
rect 10609 19193 10643 19227
rect 11253 19193 11287 19227
rect 15393 19193 15427 19227
rect 19165 19193 19199 19227
rect 20085 19193 20119 19227
rect 20821 19193 20855 19227
rect 21649 19193 21683 19227
rect 23489 19193 23523 19227
rect 25513 19193 25547 19227
rect 9413 19125 9447 19159
rect 10793 19125 10827 19159
rect 11161 19125 11195 19159
rect 12725 19125 12759 19159
rect 14197 19125 14231 19159
rect 14749 19125 14783 19159
rect 15301 19125 15335 19159
rect 16313 19125 16347 19159
rect 16865 19125 16899 19159
rect 18061 19125 18095 19159
rect 18521 19125 18555 19159
rect 19533 19125 19567 19159
rect 20177 19125 20211 19159
rect 21281 19125 21315 19159
rect 23673 19125 23707 19159
rect 24041 19125 24075 19159
rect 24133 19125 24167 19159
rect 8033 18921 8067 18955
rect 8401 18921 8435 18955
rect 9321 18921 9355 18955
rect 11621 18921 11655 18955
rect 13185 18921 13219 18955
rect 15945 18921 15979 18955
rect 19717 18921 19751 18955
rect 22109 18921 22143 18955
rect 24225 18921 24259 18955
rect 10793 18853 10827 18887
rect 11253 18853 11287 18887
rect 12050 18853 12084 18887
rect 18521 18853 18555 18887
rect 19349 18853 19383 18887
rect 20269 18853 20303 18887
rect 21649 18853 21683 18887
rect 22468 18853 22502 18887
rect 24501 18853 24535 18887
rect 8769 18785 8803 18819
rect 9321 18785 9355 18819
rect 9413 18785 9447 18819
rect 10057 18785 10091 18819
rect 11805 18785 11839 18819
rect 14197 18785 14231 18819
rect 14473 18785 14507 18819
rect 16865 18785 16899 18819
rect 17601 18785 17635 18819
rect 18429 18785 18463 18819
rect 21097 18785 21131 18819
rect 25053 18785 25087 18819
rect 25145 18785 25179 18819
rect 10149 18717 10183 18751
rect 10241 18717 10275 18751
rect 15301 18717 15335 18751
rect 16957 18717 16991 18751
rect 17141 18717 17175 18751
rect 18613 18717 18647 18751
rect 19809 18717 19843 18751
rect 20729 18717 20763 18751
rect 22201 18717 22235 18751
rect 25237 18717 25271 18751
rect 17969 18649 18003 18683
rect 9689 18581 9723 18615
rect 13737 18581 13771 18615
rect 14289 18581 14323 18615
rect 15025 18581 15059 18615
rect 16221 18581 16255 18615
rect 16497 18581 16531 18615
rect 18061 18581 18095 18615
rect 21281 18581 21315 18615
rect 23581 18581 23615 18615
rect 24685 18581 24719 18615
rect 10149 18377 10183 18411
rect 10701 18377 10735 18411
rect 11437 18377 11471 18411
rect 11897 18377 11931 18411
rect 12265 18377 12299 18411
rect 14749 18377 14783 18411
rect 21097 18377 21131 18411
rect 22017 18377 22051 18411
rect 23121 18377 23155 18411
rect 25053 18377 25087 18411
rect 14933 18309 14967 18343
rect 20821 18309 20855 18343
rect 8769 18241 8803 18275
rect 11069 18241 11103 18275
rect 13185 18241 13219 18275
rect 13829 18241 13863 18275
rect 15485 18241 15519 18275
rect 18337 18241 18371 18275
rect 20361 18241 20395 18275
rect 21925 18241 21959 18275
rect 22569 18241 22603 18275
rect 23397 18241 23431 18275
rect 9036 18173 9070 18207
rect 13645 18173 13679 18207
rect 16497 18173 16531 18207
rect 20913 18173 20947 18207
rect 21557 18173 21591 18207
rect 22477 18173 22511 18207
rect 23673 18173 23707 18207
rect 23929 18173 23963 18207
rect 8677 18105 8711 18139
rect 12817 18105 12851 18139
rect 15393 18105 15427 18139
rect 16773 18105 16807 18139
rect 17877 18105 17911 18139
rect 18604 18105 18638 18139
rect 22385 18105 22419 18139
rect 13277 18037 13311 18071
rect 13737 18037 13771 18071
rect 14289 18037 14323 18071
rect 15301 18037 15335 18071
rect 15945 18037 15979 18071
rect 16313 18037 16347 18071
rect 17325 18037 17359 18071
rect 19717 18037 19751 18071
rect 25605 18037 25639 18071
rect 9137 17833 9171 17867
rect 10701 17833 10735 17867
rect 11805 17833 11839 17867
rect 11897 17833 11931 17867
rect 12081 17833 12115 17867
rect 13645 17833 13679 17867
rect 14013 17833 14047 17867
rect 17233 17833 17267 17867
rect 17693 17833 17727 17867
rect 19165 17833 19199 17867
rect 22937 17833 22971 17867
rect 23949 17833 23983 17867
rect 24409 17833 24443 17867
rect 25329 17833 25363 17867
rect 11621 17765 11655 17799
rect 12449 17765 12483 17799
rect 8585 17697 8619 17731
rect 10057 17697 10091 17731
rect 11805 17697 11839 17731
rect 12541 17697 12575 17731
rect 13553 17697 13587 17731
rect 14105 17697 14139 17731
rect 15301 17697 15335 17731
rect 15568 17697 15602 17731
rect 18052 17697 18086 17731
rect 20453 17697 20487 17731
rect 21180 17697 21214 17731
rect 24317 17697 24351 17731
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 12725 17629 12759 17663
rect 14197 17629 14231 17663
rect 14933 17629 14967 17663
rect 17785 17629 17819 17663
rect 20913 17629 20947 17663
rect 24501 17629 24535 17663
rect 9689 17561 9723 17595
rect 16681 17561 16715 17595
rect 25053 17561 25087 17595
rect 13185 17493 13219 17527
rect 19809 17493 19843 17527
rect 20269 17493 20303 17527
rect 22293 17493 22327 17527
rect 23305 17493 23339 17527
rect 23765 17493 23799 17527
rect 9137 17289 9171 17323
rect 10517 17289 10551 17323
rect 11621 17289 11655 17323
rect 14105 17289 14139 17323
rect 15209 17289 15243 17323
rect 16129 17289 16163 17323
rect 19625 17289 19659 17323
rect 23121 17289 23155 17323
rect 25605 17289 25639 17323
rect 12081 17221 12115 17255
rect 16037 17221 16071 17255
rect 9597 17153 9631 17187
rect 9689 17153 9723 17187
rect 10977 17153 11011 17187
rect 13185 17153 13219 17187
rect 14013 17153 14047 17187
rect 14565 17153 14599 17187
rect 14749 17153 14783 17187
rect 16589 17153 16623 17187
rect 16681 17153 16715 17187
rect 17509 17153 17543 17187
rect 18705 17153 18739 17187
rect 10701 17085 10735 17119
rect 12265 17085 12299 17119
rect 12909 17085 12943 17119
rect 14473 17085 14507 17119
rect 16497 17085 16531 17119
rect 18429 17085 18463 17119
rect 20177 17085 20211 17119
rect 22201 17085 22235 17119
rect 22569 17085 22603 17119
rect 23673 17085 23707 17119
rect 9045 17017 9079 17051
rect 9505 17017 9539 17051
rect 11989 17017 12023 17051
rect 17877 17017 17911 17051
rect 20422 17017 20456 17051
rect 23940 17017 23974 17051
rect 10149 16949 10183 16983
rect 12541 16949 12575 16983
rect 13001 16949 13035 16983
rect 13645 16949 13679 16983
rect 15577 16949 15611 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 19073 16949 19107 16983
rect 20085 16949 20119 16983
rect 21557 16949 21591 16983
rect 23489 16949 23523 16983
rect 25053 16949 25087 16983
rect 9229 16745 9263 16779
rect 9873 16745 9907 16779
rect 12817 16745 12851 16779
rect 13645 16745 13679 16779
rect 14749 16745 14783 16779
rect 16313 16745 16347 16779
rect 16681 16745 16715 16779
rect 16865 16745 16899 16779
rect 18429 16745 18463 16779
rect 20269 16745 20303 16779
rect 21925 16745 21959 16779
rect 22477 16745 22511 16779
rect 24041 16745 24075 16779
rect 24501 16745 24535 16779
rect 14197 16677 14231 16711
rect 15117 16677 15151 16711
rect 17325 16677 17359 16711
rect 18889 16677 18923 16711
rect 23765 16677 23799 16711
rect 11345 16609 11379 16643
rect 11437 16609 11471 16643
rect 11704 16609 11738 16643
rect 13921 16609 13955 16643
rect 15669 16609 15703 16643
rect 15761 16609 15795 16643
rect 17233 16609 17267 16643
rect 18797 16609 18831 16643
rect 19809 16609 19843 16643
rect 21281 16609 21315 16643
rect 21373 16609 21407 16643
rect 22293 16609 22327 16643
rect 22845 16609 22879 16643
rect 24409 16609 24443 16643
rect 25053 16609 25087 16643
rect 25513 16609 25547 16643
rect 15853 16541 15887 16575
rect 17509 16541 17543 16575
rect 18061 16541 18095 16575
rect 19073 16541 19107 16575
rect 21465 16541 21499 16575
rect 22937 16541 22971 16575
rect 23029 16541 23063 16575
rect 24593 16541 24627 16575
rect 10885 16473 10919 16507
rect 15301 16405 15335 16439
rect 19441 16405 19475 16439
rect 20545 16405 20579 16439
rect 20913 16405 20947 16439
rect 11805 16201 11839 16235
rect 15393 16201 15427 16235
rect 17509 16201 17543 16235
rect 18061 16201 18095 16235
rect 19073 16201 19107 16235
rect 23489 16201 23523 16235
rect 24685 16201 24719 16235
rect 25145 16201 25179 16235
rect 12449 16133 12483 16167
rect 21649 16133 21683 16167
rect 23673 16133 23707 16167
rect 10333 16065 10367 16099
rect 11437 16065 11471 16099
rect 13001 16065 13035 16099
rect 14013 16065 14047 16099
rect 16221 16065 16255 16099
rect 18613 16065 18647 16099
rect 19993 16065 20027 16099
rect 20637 16065 20671 16099
rect 22201 16065 22235 16099
rect 24317 16065 24351 16099
rect 10701 15997 10735 16031
rect 11253 15997 11287 16031
rect 13921 15997 13955 16031
rect 14280 15997 14314 16031
rect 16681 15997 16715 16031
rect 20453 15997 20487 16031
rect 24041 15997 24075 16031
rect 25237 15997 25271 16031
rect 25973 15997 26007 16031
rect 16957 15929 16991 15963
rect 19625 15929 19659 15963
rect 21189 15929 21223 15963
rect 22109 15929 22143 15963
rect 25513 15929 25547 15963
rect 9965 15861 9999 15895
rect 10793 15861 10827 15895
rect 11161 15861 11195 15895
rect 12173 15861 12207 15895
rect 12817 15861 12851 15895
rect 12909 15861 12943 15895
rect 13461 15861 13495 15895
rect 16589 15861 16623 15895
rect 17785 15861 17819 15895
rect 18429 15861 18463 15895
rect 18521 15861 18555 15895
rect 20085 15861 20119 15895
rect 20545 15861 20579 15895
rect 21465 15861 21499 15895
rect 22017 15861 22051 15895
rect 22753 15861 22787 15895
rect 23121 15861 23155 15895
rect 24133 15861 24167 15895
rect 12725 15657 12759 15691
rect 14657 15657 14691 15691
rect 15117 15657 15151 15691
rect 16313 15657 16347 15691
rect 16773 15657 16807 15691
rect 17233 15657 17267 15691
rect 17969 15657 18003 15691
rect 18337 15657 18371 15691
rect 18981 15657 19015 15691
rect 19257 15657 19291 15691
rect 20913 15657 20947 15691
rect 22477 15657 22511 15691
rect 24501 15657 24535 15691
rect 24869 15657 24903 15691
rect 11253 15589 11287 15623
rect 11590 15589 11624 15623
rect 14197 15589 14231 15623
rect 15761 15589 15795 15623
rect 20729 15589 20763 15623
rect 25329 15589 25363 15623
rect 11345 15521 11379 15555
rect 13921 15521 13955 15555
rect 15485 15521 15519 15555
rect 17141 15521 17175 15555
rect 19625 15521 19659 15555
rect 20361 15521 20395 15555
rect 21281 15521 21315 15555
rect 22569 15521 22603 15555
rect 22836 15521 22870 15555
rect 25053 15521 25087 15555
rect 10333 15453 10367 15487
rect 17325 15453 17359 15487
rect 19717 15453 19751 15487
rect 19901 15453 19935 15487
rect 21373 15453 21407 15487
rect 21557 15453 21591 15487
rect 10793 15385 10827 15419
rect 13829 15385 13863 15419
rect 13277 15317 13311 15351
rect 16589 15317 16623 15351
rect 18705 15317 18739 15351
rect 21925 15317 21959 15351
rect 23949 15317 23983 15351
rect 10793 15113 10827 15147
rect 11805 15113 11839 15147
rect 12449 15113 12483 15147
rect 14749 15113 14783 15147
rect 17325 15113 17359 15147
rect 21189 15113 21223 15147
rect 21833 15113 21867 15147
rect 22385 15113 22419 15147
rect 23029 15113 23063 15147
rect 23397 15113 23431 15147
rect 25421 15113 25455 15147
rect 26249 15113 26283 15147
rect 10333 15045 10367 15079
rect 23673 15045 23707 15079
rect 25053 15045 25087 15079
rect 9965 14977 9999 15011
rect 11253 14977 11287 15011
rect 11345 14977 11379 15011
rect 13001 14977 13035 15011
rect 14289 14977 14323 15011
rect 15393 14977 15427 15011
rect 18797 14977 18831 15011
rect 24225 14977 24259 15011
rect 12817 14909 12851 14943
rect 14013 14909 14047 14943
rect 18613 14909 18647 14943
rect 19809 14909 19843 14943
rect 20065 14909 20099 14943
rect 22477 14909 22511 14943
rect 25237 14909 25271 14943
rect 25789 14909 25823 14943
rect 12265 14841 12299 14875
rect 12909 14841 12943 14875
rect 15660 14841 15694 14875
rect 17877 14841 17911 14875
rect 18705 14841 18739 14875
rect 19349 14841 19383 14875
rect 19717 14841 19751 14875
rect 10701 14773 10735 14807
rect 11161 14773 11195 14807
rect 13737 14773 13771 14807
rect 15301 14773 15335 14807
rect 16773 14773 16807 14807
rect 18245 14773 18279 14807
rect 22661 14773 22695 14807
rect 24041 14773 24075 14807
rect 24133 14773 24167 14807
rect 24685 14773 24719 14807
rect 10609 14569 10643 14603
rect 12725 14569 12759 14603
rect 13185 14569 13219 14603
rect 13645 14569 13679 14603
rect 14657 14569 14691 14603
rect 16037 14569 16071 14603
rect 18521 14569 18555 14603
rect 19901 14569 19935 14603
rect 20729 14569 20763 14603
rect 20913 14569 20947 14603
rect 23949 14569 23983 14603
rect 25237 14569 25271 14603
rect 19349 14501 19383 14535
rect 20269 14501 20303 14535
rect 10957 14433 10991 14467
rect 14013 14433 14047 14467
rect 15945 14433 15979 14467
rect 17397 14433 17431 14467
rect 19717 14433 19751 14467
rect 21281 14433 21315 14467
rect 22109 14433 22143 14467
rect 22836 14433 22870 14467
rect 25053 14433 25087 14467
rect 10241 14365 10275 14399
rect 10701 14365 10735 14399
rect 13553 14365 13587 14399
rect 14105 14365 14139 14399
rect 14289 14365 14323 14399
rect 16129 14365 16163 14399
rect 17141 14365 17175 14399
rect 21373 14365 21407 14399
rect 21465 14365 21499 14399
rect 22569 14365 22603 14399
rect 15577 14297 15611 14331
rect 12081 14229 12115 14263
rect 15025 14229 15059 14263
rect 16865 14229 16899 14263
rect 22477 14229 22511 14263
rect 24501 14229 24535 14263
rect 24961 14229 24995 14263
rect 10333 14025 10367 14059
rect 12173 14025 12207 14059
rect 12817 14025 12851 14059
rect 16129 14025 16163 14059
rect 18613 14025 18647 14059
rect 20177 14025 20211 14059
rect 21281 14025 21315 14059
rect 22017 14025 22051 14059
rect 25513 14025 25547 14059
rect 26065 14025 26099 14059
rect 9965 13889 9999 13923
rect 11345 13889 11379 13923
rect 13369 13889 13403 13923
rect 14381 13889 14415 13923
rect 16589 13889 16623 13923
rect 16773 13889 16807 13923
rect 17785 13889 17819 13923
rect 21833 13889 21867 13923
rect 22661 13889 22695 13923
rect 24041 13889 24075 13923
rect 11253 13821 11287 13855
rect 11805 13821 11839 13855
rect 12725 13821 12759 13855
rect 13277 13821 13311 13855
rect 17417 13821 17451 13855
rect 18797 13821 18831 13855
rect 19053 13821 19087 13855
rect 20913 13821 20947 13855
rect 23121 13821 23155 13855
rect 23489 13821 23523 13855
rect 24133 13821 24167 13855
rect 24389 13821 24423 13855
rect 10609 13753 10643 13787
rect 11161 13753 11195 13787
rect 13921 13753 13955 13787
rect 14289 13753 14323 13787
rect 14648 13753 14682 13787
rect 16957 13753 16991 13787
rect 22477 13753 22511 13787
rect 10793 13685 10827 13719
rect 13185 13685 13219 13719
rect 15761 13685 15795 13719
rect 16497 13685 16531 13719
rect 18337 13685 18371 13719
rect 22385 13685 22419 13719
rect 9781 13481 9815 13515
rect 10333 13481 10367 13515
rect 10701 13481 10735 13515
rect 12173 13481 12207 13515
rect 13645 13481 13679 13515
rect 14749 13481 14783 13515
rect 15117 13481 15151 13515
rect 17877 13481 17911 13515
rect 20269 13481 20303 13515
rect 20913 13481 20947 13515
rect 22845 13481 22879 13515
rect 23489 13481 23523 13515
rect 24041 13481 24075 13515
rect 25053 13481 25087 13515
rect 11060 13413 11094 13447
rect 16037 13413 16071 13447
rect 18245 13413 18279 13447
rect 20729 13413 20763 13447
rect 22937 13413 22971 13447
rect 10793 13345 10827 13379
rect 12909 13345 12943 13379
rect 14013 13345 14047 13379
rect 18337 13345 18371 13379
rect 19625 13345 19659 13379
rect 21281 13345 21315 13379
rect 24409 13345 24443 13379
rect 24501 13345 24535 13379
rect 25421 13345 25455 13379
rect 13553 13277 13587 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 18521 13277 18555 13311
rect 19717 13277 19751 13311
rect 19901 13277 19935 13311
rect 21373 13277 21407 13311
rect 21557 13277 21591 13311
rect 23121 13277 23155 13311
rect 23949 13277 23983 13311
rect 24593 13277 24627 13311
rect 15577 13209 15611 13243
rect 17325 13209 17359 13243
rect 22109 13209 22143 13243
rect 18889 13141 18923 13175
rect 19257 13141 19291 13175
rect 22477 13141 22511 13175
rect 9965 12937 9999 12971
rect 10793 12937 10827 12971
rect 12265 12937 12299 12971
rect 16221 12937 16255 12971
rect 18245 12937 18279 12971
rect 19717 12937 19751 12971
rect 21741 12937 21775 12971
rect 25513 12937 25547 12971
rect 15117 12869 15151 12903
rect 15761 12869 15795 12903
rect 24041 12869 24075 12903
rect 10333 12801 10367 12835
rect 11345 12801 11379 12835
rect 13645 12801 13679 12835
rect 16773 12801 16807 12835
rect 17509 12801 17543 12835
rect 18889 12801 18923 12835
rect 22569 12801 22603 12835
rect 24133 12801 24167 12835
rect 11253 12733 11287 12767
rect 12449 12733 12483 12767
rect 13185 12733 13219 12767
rect 13737 12733 13771 12767
rect 14004 12733 14038 12767
rect 17877 12733 17911 12767
rect 18705 12733 18739 12767
rect 19809 12733 19843 12767
rect 22293 12733 22327 12767
rect 10701 12665 10735 12699
rect 11161 12665 11195 12699
rect 12725 12665 12759 12699
rect 16681 12665 16715 12699
rect 19349 12665 19383 12699
rect 20054 12665 20088 12699
rect 23121 12665 23155 12699
rect 23489 12665 23523 12699
rect 24400 12665 24434 12699
rect 11897 12597 11931 12631
rect 16129 12597 16163 12631
rect 16589 12597 16623 12631
rect 18613 12597 18647 12631
rect 21189 12597 21223 12631
rect 22201 12597 22235 12631
rect 11253 12393 11287 12427
rect 13829 12393 13863 12427
rect 14197 12393 14231 12427
rect 15301 12393 15335 12427
rect 16313 12393 16347 12427
rect 16773 12393 16807 12427
rect 20177 12393 20211 12427
rect 20637 12393 20671 12427
rect 22845 12393 22879 12427
rect 23305 12393 23339 12427
rect 24961 12393 24995 12427
rect 10885 12325 10919 12359
rect 11796 12325 11830 12359
rect 15669 12325 15703 12359
rect 17601 12325 17635 12359
rect 18337 12325 18371 12359
rect 21158 12325 21192 12359
rect 23848 12325 23882 12359
rect 25513 12325 25547 12359
rect 15761 12257 15795 12291
rect 19165 12257 19199 12291
rect 20913 12257 20947 12291
rect 23581 12257 23615 12291
rect 11529 12189 11563 12223
rect 15117 12189 15151 12223
rect 15945 12189 15979 12223
rect 17693 12189 17727 12223
rect 17785 12189 17819 12223
rect 19257 12189 19291 12223
rect 19349 12189 19383 12223
rect 17233 12121 17267 12155
rect 12909 12053 12943 12087
rect 14657 12053 14691 12087
rect 17141 12053 17175 12087
rect 18705 12053 18739 12087
rect 18797 12053 18831 12087
rect 19901 12053 19935 12087
rect 22293 12053 22327 12087
rect 11621 11849 11655 11883
rect 15209 11849 15243 11883
rect 16221 11849 16255 11883
rect 17509 11849 17543 11883
rect 20637 11849 20671 11883
rect 23121 11849 23155 11883
rect 25329 11849 25363 11883
rect 20821 11781 20855 11815
rect 20913 11781 20947 11815
rect 22477 11781 22511 11815
rect 12725 11713 12759 11747
rect 16957 11713 16991 11747
rect 21097 11713 21131 11747
rect 24225 11713 24259 11747
rect 24961 11713 24995 11747
rect 12449 11645 12483 11679
rect 13185 11645 13219 11679
rect 13829 11645 13863 11679
rect 16773 11645 16807 11679
rect 18061 11645 18095 11679
rect 20821 11645 20855 11679
rect 21353 11645 21387 11679
rect 13737 11577 13771 11611
rect 14074 11577 14108 11611
rect 18328 11577 18362 11611
rect 19993 11577 20027 11611
rect 23489 11577 23523 11611
rect 24685 11577 24719 11611
rect 11897 11509 11931 11543
rect 15853 11509 15887 11543
rect 16405 11509 16439 11543
rect 16865 11509 16899 11543
rect 17785 11509 17819 11543
rect 19441 11509 19475 11543
rect 24317 11509 24351 11543
rect 24777 11509 24811 11543
rect 13829 11305 13863 11339
rect 14473 11305 14507 11339
rect 15117 11305 15151 11339
rect 16589 11305 16623 11339
rect 18429 11305 18463 11339
rect 18797 11305 18831 11339
rect 19349 11305 19383 11339
rect 20269 11305 20303 11339
rect 20913 11305 20947 11339
rect 21281 11305 21315 11339
rect 22293 11305 22327 11339
rect 22753 11305 22787 11339
rect 24225 11305 24259 11339
rect 24869 11305 24903 11339
rect 25513 11305 25547 11339
rect 12449 11169 12483 11203
rect 12716 11169 12750 11203
rect 15853 11169 15887 11203
rect 17316 11169 17350 11203
rect 15945 11101 15979 11135
rect 16037 11101 16071 11135
rect 17049 11101 17083 11135
rect 10885 11033 10919 11067
rect 15485 11033 15519 11067
rect 16865 11033 16899 11067
rect 19809 11237 19843 11271
rect 23090 11237 23124 11271
rect 19533 11169 19567 11203
rect 22845 11169 22879 11203
rect 25329 11169 25363 11203
rect 21373 11101 21407 11135
rect 21465 11101 21499 11135
rect 19073 11033 19107 11067
rect 21925 11033 21959 11067
rect 11897 10965 11931 10999
rect 12357 10965 12391 10999
rect 18797 10965 18831 10999
rect 20729 10965 20763 10999
rect 10793 10761 10827 10795
rect 14197 10761 14231 10795
rect 17049 10761 17083 10795
rect 17785 10761 17819 10795
rect 19533 10761 19567 10795
rect 19717 10761 19751 10795
rect 23397 10761 23431 10795
rect 25789 10761 25823 10795
rect 12449 10693 12483 10727
rect 18061 10693 18095 10727
rect 10701 10625 10735 10659
rect 11437 10625 11471 10659
rect 13001 10625 13035 10659
rect 13737 10625 13771 10659
rect 14657 10625 14691 10659
rect 14841 10625 14875 10659
rect 15301 10625 15335 10659
rect 16221 10625 16255 10659
rect 16405 10625 16439 10659
rect 18705 10625 18739 10659
rect 19993 10625 20027 10659
rect 21649 10625 21683 10659
rect 22569 10625 22603 10659
rect 24317 10625 24351 10659
rect 25329 10625 25363 10659
rect 11161 10557 11195 10591
rect 12909 10557 12943 10591
rect 18429 10557 18463 10591
rect 19901 10557 19935 10591
rect 21465 10557 21499 10591
rect 24133 10557 24167 10591
rect 24777 10557 24811 10591
rect 12817 10489 12851 10523
rect 15669 10489 15703 10523
rect 17417 10489 17451 10523
rect 18521 10489 18555 10523
rect 20545 10489 20579 10523
rect 20913 10489 20947 10523
rect 11253 10421 11287 10455
rect 11805 10421 11839 10455
rect 12173 10421 12207 10455
rect 14105 10421 14139 10455
rect 14565 10421 14599 10455
rect 15761 10421 15795 10455
rect 16129 10421 16163 10455
rect 19165 10421 19199 10455
rect 21005 10421 21039 10455
rect 21373 10421 21407 10455
rect 22109 10421 22143 10455
rect 22477 10421 22511 10455
rect 23029 10421 23063 10455
rect 23765 10421 23799 10455
rect 24225 10421 24259 10455
rect 12725 10217 12759 10251
rect 13277 10217 13311 10251
rect 14749 10217 14783 10251
rect 15577 10217 15611 10251
rect 16129 10217 16163 10251
rect 16681 10217 16715 10251
rect 17693 10217 17727 10251
rect 18245 10217 18279 10251
rect 19257 10217 19291 10251
rect 19625 10217 19659 10251
rect 21373 10217 21407 10251
rect 22385 10217 22419 10251
rect 22753 10217 22787 10251
rect 22937 10217 22971 10251
rect 23857 10217 23891 10251
rect 25329 10217 25363 10251
rect 14197 10149 14231 10183
rect 17601 10149 17635 10183
rect 23397 10149 23431 10183
rect 11612 10081 11646 10115
rect 14105 10081 14139 10115
rect 16037 10081 16071 10115
rect 18797 10081 18831 10115
rect 19717 10081 19751 10115
rect 21281 10081 21315 10115
rect 23949 10081 23983 10115
rect 24216 10081 24250 10115
rect 11345 10013 11379 10047
rect 16313 10013 16347 10047
rect 17877 10013 17911 10047
rect 19901 10013 19935 10047
rect 21557 10013 21591 10047
rect 15117 9945 15151 9979
rect 17233 9945 17267 9979
rect 19165 9945 19199 9979
rect 10885 9877 10919 9911
rect 13921 9877 13955 9911
rect 15669 9877 15703 9911
rect 17141 9877 17175 9911
rect 20637 9877 20671 9911
rect 20913 9877 20947 9911
rect 21925 9877 21959 9911
rect 17785 9673 17819 9707
rect 20085 9673 20119 9707
rect 21925 9673 21959 9707
rect 22661 9673 22695 9707
rect 23857 9673 23891 9707
rect 24961 9673 24995 9707
rect 25237 9673 25271 9707
rect 15117 9605 15151 9639
rect 19441 9605 19475 9639
rect 20453 9605 20487 9639
rect 11345 9537 11379 9571
rect 13001 9537 13035 9571
rect 14749 9537 14783 9571
rect 15853 9537 15887 9571
rect 16957 9537 16991 9571
rect 21005 9537 21039 9571
rect 21097 9537 21131 9571
rect 21557 9537 21591 9571
rect 24501 9537 24535 9571
rect 25421 9537 25455 9571
rect 14381 9469 14415 9503
rect 15669 9469 15703 9503
rect 16681 9469 16715 9503
rect 18061 9469 18095 9503
rect 20913 9469 20947 9503
rect 22109 9469 22143 9503
rect 12817 9401 12851 9435
rect 13829 9401 13863 9435
rect 15577 9401 15611 9435
rect 18306 9401 18340 9435
rect 23029 9401 23063 9435
rect 24317 9401 24351 9435
rect 11253 9333 11287 9367
rect 11897 9333 11931 9367
rect 12265 9333 12299 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 13461 9333 13495 9367
rect 15209 9333 15243 9367
rect 16221 9333 16255 9367
rect 17509 9333 17543 9367
rect 20545 9333 20579 9367
rect 23489 9333 23523 9367
rect 24225 9333 24259 9367
rect 12909 9129 12943 9163
rect 14013 9129 14047 9163
rect 14841 9129 14875 9163
rect 17601 9129 17635 9163
rect 19441 9129 19475 9163
rect 20085 9129 20119 9163
rect 20545 9129 20579 9163
rect 22845 9129 22879 9163
rect 24317 9129 24351 9163
rect 15844 9061 15878 9095
rect 11785 8993 11819 9027
rect 15117 8993 15151 9027
rect 18328 8993 18362 9027
rect 20729 8993 20763 9027
rect 20913 8993 20947 9027
rect 21169 8993 21203 9027
rect 24225 8993 24259 9027
rect 11529 8925 11563 8959
rect 14381 8925 14415 8959
rect 15577 8925 15611 8959
rect 18061 8925 18095 8959
rect 24409 8925 24443 8959
rect 14933 8857 14967 8891
rect 23765 8857 23799 8891
rect 10885 8789 10919 8823
rect 11437 8789 11471 8823
rect 16957 8789 16991 8823
rect 17969 8789 18003 8823
rect 20361 8789 20395 8823
rect 22293 8789 22327 8823
rect 23397 8789 23431 8823
rect 23857 8789 23891 8823
rect 10333 8585 10367 8619
rect 10793 8585 10827 8619
rect 12541 8585 12575 8619
rect 16129 8585 16163 8619
rect 16497 8585 16531 8619
rect 17877 8585 17911 8619
rect 18337 8585 18371 8619
rect 20361 8585 20395 8619
rect 23121 8585 23155 8619
rect 23489 8585 23523 8619
rect 25237 8585 25271 8619
rect 11989 8517 12023 8551
rect 15485 8517 15519 8551
rect 11437 8449 11471 8483
rect 13185 8449 13219 8483
rect 13553 8449 13587 8483
rect 14013 8449 14047 8483
rect 22017 8449 22051 8483
rect 11805 8381 11839 8415
rect 11989 8381 12023 8415
rect 12265 8381 12299 8415
rect 13001 8381 13035 8415
rect 14105 8381 14139 8415
rect 14372 8381 14406 8415
rect 18981 8381 19015 8415
rect 21281 8381 21315 8415
rect 21833 8381 21867 8415
rect 23857 8381 23891 8415
rect 10701 8313 10735 8347
rect 11253 8313 11287 8347
rect 12909 8313 12943 8347
rect 16589 8313 16623 8347
rect 18889 8313 18923 8347
rect 19226 8313 19260 8347
rect 21925 8313 21959 8347
rect 22477 8313 22511 8347
rect 24124 8313 24158 8347
rect 11161 8245 11195 8279
rect 17417 8245 17451 8279
rect 21005 8245 21039 8279
rect 21465 8245 21499 8279
rect 12541 8041 12575 8075
rect 14013 8041 14047 8075
rect 15301 8041 15335 8075
rect 15669 8041 15703 8075
rect 17785 8041 17819 8075
rect 18061 8041 18095 8075
rect 18705 8041 18739 8075
rect 21281 8041 21315 8075
rect 23949 8041 23983 8075
rect 25053 8041 25087 8075
rect 10149 7973 10183 8007
rect 14105 7973 14139 8007
rect 15761 7973 15795 8007
rect 17233 7973 17267 8007
rect 19257 7973 19291 8007
rect 19717 7973 19751 8007
rect 21373 7973 21407 8007
rect 9873 7905 9907 7939
rect 11417 7905 11451 7939
rect 16313 7905 16347 7939
rect 18613 7905 18647 7939
rect 22825 7905 22859 7939
rect 11161 7837 11195 7871
rect 14289 7837 14323 7871
rect 15945 7837 15979 7871
rect 18797 7837 18831 7871
rect 19809 7837 19843 7871
rect 21465 7837 21499 7871
rect 22569 7837 22603 7871
rect 22109 7769 22143 7803
rect 10885 7701 10919 7735
rect 13093 7701 13127 7735
rect 13645 7701 13679 7735
rect 15117 7701 15151 7735
rect 18245 7701 18279 7735
rect 20545 7701 20579 7735
rect 20913 7701 20947 7735
rect 22477 7701 22511 7735
rect 24501 7701 24535 7735
rect 9413 7497 9447 7531
rect 11253 7497 11287 7531
rect 11805 7497 11839 7531
rect 12173 7497 12207 7531
rect 12449 7497 12483 7531
rect 14105 7497 14139 7531
rect 16129 7497 16163 7531
rect 16405 7497 16439 7531
rect 17877 7497 17911 7531
rect 20453 7497 20487 7531
rect 21465 7497 21499 7531
rect 21833 7497 21867 7531
rect 13737 7429 13771 7463
rect 16773 7429 16807 7463
rect 20361 7429 20395 7463
rect 13001 7361 13035 7395
rect 15485 7361 15519 7395
rect 15669 7361 15703 7395
rect 19441 7361 19475 7395
rect 21097 7361 21131 7395
rect 22661 7361 22695 7395
rect 23489 7361 23523 7395
rect 9045 7293 9079 7327
rect 9873 7293 9907 7327
rect 12909 7293 12943 7327
rect 14565 7293 14599 7327
rect 18705 7293 18739 7327
rect 19257 7293 19291 7327
rect 19901 7293 19935 7327
rect 20821 7293 20855 7327
rect 23673 7293 23707 7327
rect 23940 7293 23974 7327
rect 9781 7225 9815 7259
rect 10118 7225 10152 7259
rect 14841 7225 14875 7259
rect 15393 7225 15427 7259
rect 20913 7225 20947 7259
rect 12817 7157 12851 7191
rect 14381 7157 14415 7191
rect 15025 7157 15059 7191
rect 16957 7157 16991 7191
rect 17509 7157 17543 7191
rect 18337 7157 18371 7191
rect 18889 7157 18923 7191
rect 19349 7157 19383 7191
rect 22017 7157 22051 7191
rect 22385 7157 22419 7191
rect 22477 7157 22511 7191
rect 23121 7157 23155 7191
rect 25053 7157 25087 7191
rect 11069 6953 11103 6987
rect 12081 6953 12115 6987
rect 12173 6953 12207 6987
rect 12541 6953 12575 6987
rect 13737 6953 13771 6987
rect 14289 6953 14323 6987
rect 14565 6953 14599 6987
rect 15117 6953 15151 6987
rect 16681 6953 16715 6987
rect 17417 6953 17451 6987
rect 17969 6953 18003 6987
rect 22385 6953 22419 6987
rect 12633 6885 12667 6919
rect 9956 6817 9990 6851
rect 15301 6817 15335 6851
rect 15568 6817 15602 6851
rect 17877 6817 17911 6851
rect 18153 6817 18187 6851
rect 18501 6817 18535 6851
rect 20545 6817 20579 6851
rect 21261 6817 21295 6851
rect 23397 6817 23431 6851
rect 23857 6817 23891 6851
rect 9689 6749 9723 6783
rect 12725 6749 12759 6783
rect 13461 6749 13495 6783
rect 18245 6749 18279 6783
rect 21005 6749 21039 6783
rect 23949 6749 23983 6783
rect 24041 6749 24075 6783
rect 25053 6749 25087 6783
rect 23029 6681 23063 6715
rect 11713 6613 11747 6647
rect 19625 6613 19659 6647
rect 23489 6613 23523 6647
rect 24501 6613 24535 6647
rect 7849 6409 7883 6443
rect 10793 6409 10827 6443
rect 11897 6409 11931 6443
rect 12265 6409 12299 6443
rect 15945 6409 15979 6443
rect 17509 6409 17543 6443
rect 21097 6409 21131 6443
rect 21649 6409 21683 6443
rect 22109 6409 22143 6443
rect 24409 6409 24443 6443
rect 9413 6341 9447 6375
rect 12725 6341 12759 6375
rect 23489 6341 23523 6375
rect 10333 6273 10367 6307
rect 11437 6273 11471 6307
rect 13829 6273 13863 6307
rect 14013 6273 14047 6307
rect 15393 6273 15427 6307
rect 15577 6273 15611 6307
rect 17877 6273 17911 6307
rect 18705 6273 18739 6307
rect 24961 6273 24995 6307
rect 8033 6205 8067 6239
rect 8289 6205 8323 6239
rect 10701 6205 10735 6239
rect 11161 6205 11195 6239
rect 13277 6205 13311 6239
rect 13737 6205 13771 6239
rect 16865 6205 16899 6239
rect 18521 6205 18555 6239
rect 19717 6205 19751 6239
rect 22201 6205 22235 6239
rect 22753 6205 22787 6239
rect 24317 6205 24351 6239
rect 24869 6205 24903 6239
rect 11253 6137 11287 6171
rect 15301 6137 15335 6171
rect 16773 6137 16807 6171
rect 19962 6137 19996 6171
rect 13369 6069 13403 6103
rect 14381 6069 14415 6103
rect 14749 6069 14783 6103
rect 14933 6069 14967 6103
rect 16313 6069 16347 6103
rect 17049 6069 17083 6103
rect 18153 6069 18187 6103
rect 18613 6069 18647 6103
rect 19165 6069 19199 6103
rect 19533 6069 19567 6103
rect 22385 6069 22419 6103
rect 23949 6069 23983 6103
rect 24777 6069 24811 6103
rect 8125 5865 8159 5899
rect 9965 5865 9999 5899
rect 11713 5865 11747 5899
rect 12817 5865 12851 5899
rect 13461 5865 13495 5899
rect 14013 5865 14047 5899
rect 15485 5865 15519 5899
rect 17141 5865 17175 5899
rect 17785 5865 17819 5899
rect 18153 5865 18187 5899
rect 19625 5865 19659 5899
rect 20269 5865 20303 5899
rect 20637 5865 20671 5899
rect 22385 5865 22419 5899
rect 23029 5865 23063 5899
rect 23857 5865 23891 5899
rect 24593 5865 24627 5899
rect 18490 5797 18524 5831
rect 21250 5797 21284 5831
rect 23305 5797 23339 5831
rect 10333 5729 10367 5763
rect 12081 5729 12115 5763
rect 16017 5729 16051 5763
rect 18245 5729 18279 5763
rect 21005 5729 21039 5763
rect 25053 5729 25087 5763
rect 10793 5661 10827 5695
rect 12173 5661 12207 5695
rect 12357 5661 12391 5695
rect 14105 5661 14139 5695
rect 14197 5661 14231 5695
rect 15761 5661 15795 5695
rect 23949 5661 23983 5695
rect 24041 5661 24075 5695
rect 14933 5593 14967 5627
rect 13645 5525 13679 5559
rect 23489 5525 23523 5559
rect 24869 5525 24903 5559
rect 25237 5525 25271 5559
rect 11253 5321 11287 5355
rect 13737 5321 13771 5355
rect 14013 5321 14047 5355
rect 15577 5321 15611 5355
rect 16129 5321 16163 5355
rect 23121 5321 23155 5355
rect 25789 5321 25823 5355
rect 12633 5253 12667 5287
rect 23489 5253 23523 5287
rect 11345 5185 11379 5219
rect 13093 5185 13127 5219
rect 13277 5185 13311 5219
rect 18797 5185 18831 5219
rect 19625 5185 19659 5219
rect 20361 5185 20395 5219
rect 21097 5185 21131 5219
rect 12265 5117 12299 5151
rect 12541 5117 12575 5151
rect 14197 5117 14231 5151
rect 14453 5117 14487 5151
rect 16865 5117 16899 5151
rect 17417 5117 17451 5151
rect 20177 5117 20211 5151
rect 21373 5117 21407 5151
rect 21925 5117 21959 5151
rect 22477 5117 22511 5151
rect 23857 5117 23891 5151
rect 11897 5049 11931 5083
rect 17877 5049 17911 5083
rect 18613 5049 18647 5083
rect 22385 5049 22419 5083
rect 24124 5049 24158 5083
rect 12541 4981 12575 5015
rect 13001 4981 13035 5015
rect 16589 4981 16623 5015
rect 17049 4981 17083 5015
rect 18245 4981 18279 5015
rect 18705 4981 18739 5015
rect 19257 4981 19291 5015
rect 19809 4981 19843 5015
rect 20269 4981 20303 5015
rect 21557 4981 21591 5015
rect 22661 4981 22695 5015
rect 25237 4981 25271 5015
rect 12081 4777 12115 4811
rect 12449 4777 12483 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 14841 4777 14875 4811
rect 15669 4777 15703 4811
rect 16313 4777 16347 4811
rect 18337 4777 18371 4811
rect 19901 4777 19935 4811
rect 23029 4777 23063 4811
rect 23397 4777 23431 4811
rect 24593 4777 24627 4811
rect 25053 4777 25087 4811
rect 11805 4709 11839 4743
rect 12817 4709 12851 4743
rect 18245 4709 18279 4743
rect 18705 4709 18739 4743
rect 19441 4709 19475 4743
rect 20545 4709 20579 4743
rect 21373 4709 21407 4743
rect 24409 4709 24443 4743
rect 24961 4709 24995 4743
rect 14105 4641 14139 4675
rect 15761 4641 15795 4675
rect 16865 4641 16899 4675
rect 21925 4641 21959 4675
rect 12909 4573 12943 4607
rect 13093 4573 13127 4607
rect 15945 4573 15979 4607
rect 17049 4573 17083 4607
rect 18797 4573 18831 4607
rect 18981 4573 19015 4607
rect 20913 4573 20947 4607
rect 23489 4573 23523 4607
rect 23673 4573 23707 4607
rect 25145 4573 25179 4607
rect 14289 4505 14323 4539
rect 15301 4505 15335 4539
rect 17601 4505 17635 4539
rect 16773 4437 16807 4471
rect 20177 4437 20211 4471
rect 22109 4437 22143 4471
rect 22569 4437 22603 4471
rect 22845 4437 22879 4471
rect 24133 4437 24167 4471
rect 13001 4233 13035 4267
rect 13369 4233 13403 4267
rect 14841 4233 14875 4267
rect 15945 4233 15979 4267
rect 17877 4233 17911 4267
rect 18981 4233 19015 4267
rect 21465 4233 21499 4267
rect 21925 4233 21959 4267
rect 23121 4233 23155 4267
rect 25605 4233 25639 4267
rect 11897 4165 11931 4199
rect 14381 4165 14415 4199
rect 15301 4097 15335 4131
rect 15393 4097 15427 4131
rect 16313 4097 16347 4131
rect 18337 4097 18371 4131
rect 22569 4097 22603 4131
rect 23489 4097 23523 4131
rect 11253 4029 11287 4063
rect 12173 4029 12207 4063
rect 12449 4029 12483 4063
rect 13553 4029 13587 4063
rect 16405 4029 16439 4063
rect 17509 4029 17543 4063
rect 18153 4029 18187 4063
rect 19441 4029 19475 4063
rect 22385 4029 22419 4063
rect 22477 4029 22511 4063
rect 23673 4029 23707 4063
rect 13829 3961 13863 3995
rect 16681 3961 16715 3995
rect 19686 3961 19720 3995
rect 23918 3961 23952 3995
rect 11161 3893 11195 3927
rect 11437 3893 11471 3927
rect 12633 3893 12667 3927
rect 14749 3893 14783 3927
rect 15209 3893 15243 3927
rect 19349 3893 19383 3927
rect 20821 3893 20855 3927
rect 22017 3893 22051 3927
rect 25053 3893 25087 3927
rect 11345 3689 11379 3723
rect 13001 3689 13035 3723
rect 13369 3689 13403 3723
rect 14473 3689 14507 3723
rect 16129 3689 16163 3723
rect 18705 3689 18739 3723
rect 19257 3689 19291 3723
rect 19625 3689 19659 3723
rect 19717 3689 19751 3723
rect 20269 3689 20303 3723
rect 22937 3689 22971 3723
rect 23673 3689 23707 3723
rect 24409 3689 24443 3723
rect 25053 3689 25087 3723
rect 25421 3689 25455 3723
rect 10149 3621 10183 3655
rect 15577 3621 15611 3655
rect 20637 3621 20671 3655
rect 21373 3621 21407 3655
rect 24501 3621 24535 3655
rect 11161 3553 11195 3587
rect 12265 3553 12299 3587
rect 13737 3553 13771 3587
rect 14841 3553 14875 3587
rect 15301 3553 15335 3587
rect 17040 3553 17074 3587
rect 21557 3553 21591 3587
rect 21824 3553 21858 3587
rect 13829 3485 13863 3519
rect 14013 3485 14047 3519
rect 16773 3485 16807 3519
rect 19901 3485 19935 3519
rect 24593 3485 24627 3519
rect 12173 3349 12207 3383
rect 12449 3349 12483 3383
rect 16589 3349 16623 3383
rect 18153 3349 18187 3383
rect 19073 3349 19107 3383
rect 24041 3349 24075 3383
rect 10793 3145 10827 3179
rect 11161 3145 11195 3179
rect 11805 3145 11839 3179
rect 12265 3145 12299 3179
rect 12633 3145 12667 3179
rect 14289 3145 14323 3179
rect 14841 3145 14875 3179
rect 15209 3145 15243 3179
rect 17785 3145 17819 3179
rect 18061 3145 18095 3179
rect 19349 3145 19383 3179
rect 21833 3145 21867 3179
rect 22385 3145 22419 3179
rect 23121 3145 23155 3179
rect 23489 3145 23523 3179
rect 24409 3145 24443 3179
rect 24777 3145 24811 3179
rect 25513 3145 25547 3179
rect 10333 3077 10367 3111
rect 11437 3077 11471 3111
rect 25145 3077 25179 3111
rect 18613 3009 18647 3043
rect 19717 3009 19751 3043
rect 20361 3009 20395 3043
rect 10149 2941 10183 2975
rect 11253 2941 11287 2975
rect 12909 2941 12943 2975
rect 13165 2941 13199 2975
rect 15393 2941 15427 2975
rect 15649 2941 15683 2975
rect 18429 2941 18463 2975
rect 20453 2941 20487 2975
rect 20720 2941 20754 2975
rect 23673 2941 23707 2975
rect 24961 2941 24995 2975
rect 23949 2873 23983 2907
rect 16773 2805 16807 2839
rect 17325 2805 17359 2839
rect 18521 2805 18555 2839
rect 10885 2601 10919 2635
rect 12633 2601 12667 2635
rect 14013 2601 14047 2635
rect 15301 2601 15335 2635
rect 16313 2601 16347 2635
rect 17325 2601 17359 2635
rect 17785 2601 17819 2635
rect 18153 2601 18187 2635
rect 19717 2601 19751 2635
rect 21189 2601 21223 2635
rect 22201 2601 22235 2635
rect 22569 2601 22603 2635
rect 23673 2601 23707 2635
rect 11345 2533 11379 2567
rect 24317 2533 24351 2567
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 12449 2465 12483 2499
rect 13001 2465 13035 2499
rect 14289 2465 14323 2499
rect 16681 2465 16715 2499
rect 18337 2465 18371 2499
rect 18593 2465 18627 2499
rect 20913 2465 20947 2499
rect 21557 2465 21591 2499
rect 22753 2465 22787 2499
rect 23305 2465 23339 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25329 2465 25363 2499
rect 25881 2465 25915 2499
rect 13093 2397 13127 2431
rect 13277 2397 13311 2431
rect 15853 2397 15887 2431
rect 16773 2397 16807 2431
rect 16957 2397 16991 2431
rect 20637 2397 20671 2431
rect 21649 2397 21683 2431
rect 21833 2397 21867 2431
rect 13737 2329 13771 2363
rect 22937 2329 22971 2363
rect 25513 2329 25547 2363
rect 10517 2261 10551 2295
rect 11621 2261 11655 2295
rect 14473 2261 14507 2295
rect 14841 2261 14875 2295
rect 16129 2261 16163 2295
<< metal1 >>
rect 21634 26664 21640 26716
rect 21692 26704 21698 26716
rect 24762 26704 24768 26716
rect 21692 26676 24768 26704
rect 21692 26664 21698 26676
rect 24762 26664 24768 26676
rect 24820 26664 24826 26716
rect 16114 26392 16120 26444
rect 16172 26432 16178 26444
rect 24578 26432 24584 26444
rect 16172 26404 24584 26432
rect 16172 26392 16178 26404
rect 24578 26392 24584 26404
rect 24636 26392 24642 26444
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 16393 25483 16451 25489
rect 16393 25449 16405 25483
rect 16439 25480 16451 25483
rect 18690 25480 18696 25492
rect 16439 25452 18696 25480
rect 16439 25449 16451 25452
rect 16393 25443 16451 25449
rect 18690 25440 18696 25452
rect 18748 25440 18754 25492
rect 20165 25483 20223 25489
rect 20165 25449 20177 25483
rect 20211 25449 20223 25483
rect 20165 25443 20223 25449
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25480 23075 25483
rect 24670 25480 24676 25492
rect 23063 25452 24676 25480
rect 23063 25449 23075 25452
rect 23017 25443 23075 25449
rect 20180 25412 20208 25443
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 26878 25412 26884 25424
rect 20180 25384 26884 25412
rect 26878 25372 26884 25384
rect 26936 25372 26942 25424
rect 16209 25347 16267 25353
rect 16209 25313 16221 25347
rect 16255 25344 16267 25347
rect 16390 25344 16396 25356
rect 16255 25316 16396 25344
rect 16255 25313 16267 25316
rect 16209 25307 16267 25313
rect 16390 25304 16396 25316
rect 16448 25304 16454 25356
rect 18874 25344 18880 25356
rect 18835 25316 18880 25344
rect 18874 25304 18880 25316
rect 18932 25304 18938 25356
rect 19981 25347 20039 25353
rect 19981 25313 19993 25347
rect 20027 25344 20039 25347
rect 20254 25344 20260 25356
rect 20027 25316 20260 25344
rect 20027 25313 20039 25316
rect 19981 25307 20039 25313
rect 20254 25304 20260 25316
rect 20312 25304 20318 25356
rect 21729 25347 21787 25353
rect 21729 25313 21741 25347
rect 21775 25344 21787 25347
rect 21818 25344 21824 25356
rect 21775 25316 21824 25344
rect 21775 25313 21787 25316
rect 21729 25307 21787 25313
rect 21818 25304 21824 25316
rect 21876 25304 21882 25356
rect 22830 25344 22836 25356
rect 22791 25316 22836 25344
rect 22830 25304 22836 25316
rect 22888 25304 22894 25356
rect 24026 25304 24032 25356
rect 24084 25344 24090 25356
rect 24581 25347 24639 25353
rect 24581 25344 24593 25347
rect 24084 25316 24593 25344
rect 24084 25304 24090 25316
rect 24581 25313 24593 25316
rect 24627 25313 24639 25347
rect 24581 25307 24639 25313
rect 26142 25276 26148 25288
rect 19076 25248 26148 25276
rect 19076 25217 19104 25248
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 19061 25211 19119 25217
rect 19061 25177 19073 25211
rect 19107 25177 19119 25211
rect 19061 25171 19119 25177
rect 21913 25211 21971 25217
rect 21913 25177 21925 25211
rect 21959 25208 21971 25211
rect 24118 25208 24124 25220
rect 21959 25180 24124 25208
rect 21959 25177 21971 25180
rect 21913 25171 21971 25177
rect 24118 25168 24124 25180
rect 24176 25168 24182 25220
rect 24762 25140 24768 25152
rect 24723 25112 24768 25140
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 16945 24803 17003 24809
rect 16945 24769 16957 24803
rect 16991 24800 17003 24803
rect 17862 24800 17868 24812
rect 16991 24772 17868 24800
rect 16991 24769 17003 24772
rect 16945 24763 17003 24769
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 12529 24735 12587 24741
rect 12529 24701 12541 24735
rect 12575 24732 12587 24735
rect 12575 24704 12940 24732
rect 12575 24701 12587 24704
rect 12529 24695 12587 24701
rect 12912 24608 12940 24704
rect 13170 24692 13176 24744
rect 13228 24732 13234 24744
rect 13633 24735 13691 24741
rect 13633 24732 13645 24735
rect 13228 24704 13645 24732
rect 13228 24692 13234 24704
rect 13633 24701 13645 24704
rect 13679 24732 13691 24735
rect 14185 24735 14243 24741
rect 14185 24732 14197 24735
rect 13679 24704 14197 24732
rect 13679 24701 13691 24704
rect 13633 24695 13691 24701
rect 14185 24701 14197 24704
rect 14231 24701 14243 24735
rect 14185 24695 14243 24701
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 14737 24735 14795 24741
rect 14737 24732 14749 24735
rect 14424 24704 14749 24732
rect 14424 24692 14430 24704
rect 14737 24701 14749 24704
rect 14783 24732 14795 24735
rect 15289 24735 15347 24741
rect 15289 24732 15301 24735
rect 14783 24704 15301 24732
rect 14783 24701 14795 24704
rect 14737 24695 14795 24701
rect 15289 24701 15301 24704
rect 15335 24701 15347 24735
rect 15289 24695 15347 24701
rect 15841 24735 15899 24741
rect 15841 24701 15853 24735
rect 15887 24732 15899 24735
rect 16298 24732 16304 24744
rect 15887 24704 16304 24732
rect 15887 24701 15899 24704
rect 15841 24695 15899 24701
rect 16298 24692 16304 24704
rect 16356 24692 16362 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 17788 24704 18061 24732
rect 15102 24664 15108 24676
rect 13832 24636 15108 24664
rect 12710 24596 12716 24608
rect 12671 24568 12716 24596
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 12894 24556 12900 24608
rect 12952 24596 12958 24608
rect 13832 24605 13860 24636
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 16482 24664 16488 24676
rect 16040 24636 16488 24664
rect 13081 24599 13139 24605
rect 13081 24596 13093 24599
rect 12952 24568 13093 24596
rect 12952 24556 12958 24568
rect 13081 24565 13093 24568
rect 13127 24565 13139 24599
rect 13081 24559 13139 24565
rect 13817 24599 13875 24605
rect 13817 24565 13829 24599
rect 13863 24565 13875 24599
rect 14918 24596 14924 24608
rect 14879 24568 14924 24596
rect 13817 24559 13875 24565
rect 14918 24556 14924 24568
rect 14976 24556 14982 24608
rect 16040 24605 16068 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 16025 24599 16083 24605
rect 16025 24565 16037 24599
rect 16071 24565 16083 24599
rect 16025 24559 16083 24565
rect 16298 24556 16304 24608
rect 16356 24596 16362 24608
rect 16393 24599 16451 24605
rect 16393 24596 16405 24599
rect 16356 24568 16405 24596
rect 16356 24556 16362 24568
rect 16393 24565 16405 24568
rect 16439 24565 16451 24599
rect 16393 24559 16451 24565
rect 16574 24556 16580 24608
rect 16632 24596 16638 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16632 24568 16773 24596
rect 16632 24556 16638 24568
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 16761 24559 16819 24565
rect 17218 24556 17224 24608
rect 17276 24596 17282 24608
rect 17788 24605 17816 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 18690 24692 18696 24744
rect 18748 24732 18754 24744
rect 19337 24735 19395 24741
rect 19337 24732 19349 24735
rect 18748 24704 19349 24732
rect 18748 24692 18754 24704
rect 19337 24701 19349 24704
rect 19383 24732 19395 24735
rect 19521 24735 19579 24741
rect 19521 24732 19533 24735
rect 19383 24704 19533 24732
rect 19383 24701 19395 24704
rect 19337 24695 19395 24701
rect 19521 24701 19533 24704
rect 19567 24701 19579 24735
rect 19521 24695 19579 24701
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24732 20867 24735
rect 20901 24735 20959 24741
rect 20901 24732 20913 24735
rect 20855 24704 20913 24732
rect 20855 24701 20867 24704
rect 20809 24695 20867 24701
rect 20901 24701 20913 24704
rect 20947 24732 20959 24735
rect 21726 24732 21732 24744
rect 20947 24704 21732 24732
rect 20947 24701 20959 24704
rect 20901 24695 20959 24701
rect 21726 24692 21732 24704
rect 21784 24692 21790 24744
rect 22005 24735 22063 24741
rect 22005 24701 22017 24735
rect 22051 24732 22063 24735
rect 22186 24732 22192 24744
rect 22051 24704 22192 24732
rect 22051 24701 22063 24704
rect 22005 24695 22063 24701
rect 22186 24692 22192 24704
rect 22244 24692 22250 24744
rect 24578 24732 24584 24744
rect 24539 24704 24584 24732
rect 24578 24692 24584 24704
rect 24636 24732 24642 24744
rect 25133 24735 25191 24741
rect 25133 24732 25145 24735
rect 24636 24704 25145 24732
rect 24636 24692 24642 24704
rect 25133 24701 25145 24704
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 19242 24664 19248 24676
rect 18248 24636 19248 24664
rect 18248 24605 18276 24636
rect 19242 24624 19248 24636
rect 19300 24624 19306 24676
rect 20622 24664 20628 24676
rect 19720 24636 20628 24664
rect 17773 24599 17831 24605
rect 17773 24596 17785 24599
rect 17276 24568 17785 24596
rect 17276 24556 17282 24568
rect 17773 24565 17785 24568
rect 17819 24565 17831 24599
rect 17773 24559 17831 24565
rect 18233 24599 18291 24605
rect 18233 24565 18245 24599
rect 18279 24565 18291 24599
rect 18233 24559 18291 24565
rect 18414 24556 18420 24608
rect 18472 24596 18478 24608
rect 18874 24596 18880 24608
rect 18472 24568 18880 24596
rect 18472 24556 18478 24568
rect 18874 24556 18880 24568
rect 18932 24556 18938 24608
rect 19720 24605 19748 24636
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 21818 24664 21824 24676
rect 20732 24636 21824 24664
rect 20732 24608 20760 24636
rect 21818 24624 21824 24636
rect 21876 24624 21882 24676
rect 22738 24664 22744 24676
rect 22204 24636 22744 24664
rect 19705 24599 19763 24605
rect 19705 24565 19717 24599
rect 19751 24565 19763 24599
rect 19705 24559 19763 24565
rect 20165 24599 20223 24605
rect 20165 24565 20177 24599
rect 20211 24596 20223 24599
rect 20254 24596 20260 24608
rect 20211 24568 20260 24596
rect 20211 24565 20223 24568
rect 20165 24559 20223 24565
rect 20254 24556 20260 24568
rect 20312 24556 20318 24608
rect 20714 24556 20720 24608
rect 20772 24556 20778 24608
rect 21082 24596 21088 24608
rect 21043 24568 21088 24596
rect 21082 24556 21088 24568
rect 21140 24556 21146 24608
rect 22204 24605 22232 24636
rect 22738 24624 22744 24636
rect 22796 24624 22802 24676
rect 22189 24599 22247 24605
rect 22189 24565 22201 24599
rect 22235 24565 22247 24599
rect 22830 24596 22836 24608
rect 22791 24568 22836 24596
rect 22189 24559 22247 24565
rect 22830 24556 22836 24568
rect 22888 24556 22894 24608
rect 24026 24556 24032 24608
rect 24084 24596 24090 24608
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 24084 24568 24409 24596
rect 24084 24556 24090 24568
rect 24397 24565 24409 24568
rect 24443 24565 24455 24599
rect 24397 24559 24455 24565
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 24765 24599 24823 24605
rect 24765 24596 24777 24599
rect 24728 24568 24777 24596
rect 24728 24556 24734 24568
rect 24765 24565 24777 24568
rect 24811 24565 24823 24599
rect 24765 24559 24823 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 15838 24392 15844 24404
rect 15799 24364 15844 24392
rect 15838 24352 15844 24364
rect 15896 24352 15902 24404
rect 17129 24395 17187 24401
rect 17129 24361 17141 24395
rect 17175 24392 17187 24395
rect 17310 24392 17316 24404
rect 17175 24364 17316 24392
rect 17175 24361 17187 24364
rect 17129 24355 17187 24361
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 17954 24352 17960 24404
rect 18012 24392 18018 24404
rect 18233 24395 18291 24401
rect 18233 24392 18245 24395
rect 18012 24364 18245 24392
rect 18012 24352 18018 24364
rect 18233 24361 18245 24364
rect 18279 24361 18291 24395
rect 18233 24355 18291 24361
rect 19429 24395 19487 24401
rect 19429 24361 19441 24395
rect 19475 24392 19487 24395
rect 20070 24392 20076 24404
rect 19475 24364 20076 24392
rect 19475 24361 19487 24364
rect 19429 24355 19487 24361
rect 20070 24352 20076 24364
rect 20128 24352 20134 24404
rect 21177 24395 21235 24401
rect 21177 24361 21189 24395
rect 21223 24392 21235 24395
rect 22002 24392 22008 24404
rect 21223 24364 22008 24392
rect 21223 24361 21235 24364
rect 21177 24355 21235 24361
rect 22002 24352 22008 24364
rect 22060 24352 22066 24404
rect 22557 24395 22615 24401
rect 22557 24361 22569 24395
rect 22603 24392 22615 24395
rect 23382 24392 23388 24404
rect 22603 24364 23388 24392
rect 22603 24361 22615 24364
rect 22557 24355 22615 24361
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 23658 24392 23664 24404
rect 23619 24364 23664 24392
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 12710 24216 12716 24268
rect 12768 24256 12774 24268
rect 13173 24259 13231 24265
rect 13173 24256 13185 24259
rect 12768 24228 13185 24256
rect 12768 24216 12774 24228
rect 13173 24225 13185 24228
rect 13219 24225 13231 24259
rect 13173 24219 13231 24225
rect 14734 24216 14740 24268
rect 14792 24256 14798 24268
rect 15749 24259 15807 24265
rect 15749 24256 15761 24259
rect 14792 24228 15761 24256
rect 14792 24216 14798 24228
rect 15749 24225 15761 24228
rect 15795 24225 15807 24259
rect 16942 24256 16948 24268
rect 16903 24228 16948 24256
rect 15749 24219 15807 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17586 24216 17592 24268
rect 17644 24256 17650 24268
rect 18049 24259 18107 24265
rect 18049 24256 18061 24259
rect 17644 24228 18061 24256
rect 17644 24216 17650 24228
rect 18049 24225 18061 24228
rect 18095 24225 18107 24259
rect 18049 24219 18107 24225
rect 19245 24259 19303 24265
rect 19245 24225 19257 24259
rect 19291 24256 19303 24259
rect 20162 24256 20168 24268
rect 19291 24228 20168 24256
rect 19291 24225 19303 24228
rect 19245 24219 19303 24225
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 20990 24256 20996 24268
rect 20951 24228 20996 24256
rect 20990 24216 20996 24228
rect 21048 24216 21054 24268
rect 22370 24256 22376 24268
rect 22331 24228 22376 24256
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 23474 24256 23480 24268
rect 23435 24228 23480 24256
rect 23474 24216 23480 24228
rect 23532 24216 23538 24268
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 24762 24256 24768 24268
rect 24627 24228 24768 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 24762 24216 24768 24228
rect 24820 24216 24826 24268
rect 13262 24188 13268 24200
rect 13223 24160 13268 24188
rect 13262 24148 13268 24160
rect 13320 24148 13326 24200
rect 13354 24148 13360 24200
rect 13412 24188 13418 24200
rect 16022 24188 16028 24200
rect 13412 24160 13457 24188
rect 15983 24160 16028 24188
rect 13412 24148 13418 24160
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 10873 24055 10931 24061
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11330 24052 11336 24064
rect 10919 24024 11336 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11330 24012 11336 24024
rect 11388 24052 11394 24064
rect 12437 24055 12495 24061
rect 12437 24052 12449 24055
rect 11388 24024 12449 24052
rect 11388 24012 11394 24024
rect 12437 24021 12449 24024
rect 12483 24052 12495 24055
rect 12526 24052 12532 24064
rect 12483 24024 12532 24052
rect 12483 24021 12495 24024
rect 12437 24015 12495 24021
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 12802 24052 12808 24064
rect 12763 24024 12808 24052
rect 12802 24012 12808 24024
rect 12860 24012 12866 24064
rect 14826 24012 14832 24064
rect 14884 24052 14890 24064
rect 14921 24055 14979 24061
rect 14921 24052 14933 24055
rect 14884 24024 14933 24052
rect 14884 24012 14890 24024
rect 14921 24021 14933 24024
rect 14967 24021 14979 24055
rect 14921 24015 14979 24021
rect 15381 24055 15439 24061
rect 15381 24021 15393 24055
rect 15427 24052 15439 24055
rect 16482 24052 16488 24064
rect 15427 24024 16488 24052
rect 15427 24021 15439 24024
rect 15381 24015 15439 24021
rect 16482 24012 16488 24024
rect 16540 24012 16546 24064
rect 22097 24055 22155 24061
rect 22097 24021 22109 24055
rect 22143 24052 22155 24055
rect 22186 24052 22192 24064
rect 22143 24024 22192 24052
rect 22143 24021 22155 24024
rect 22097 24015 22155 24021
rect 22186 24012 22192 24024
rect 22244 24012 22250 24064
rect 24118 24012 24124 24064
rect 24176 24052 24182 24064
rect 24765 24055 24823 24061
rect 24765 24052 24777 24055
rect 24176 24024 24777 24052
rect 24176 24012 24182 24024
rect 24765 24021 24777 24024
rect 24811 24021 24823 24055
rect 24765 24015 24823 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 10778 23848 10784 23860
rect 10739 23820 10784 23848
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 13906 23808 13912 23860
rect 13964 23848 13970 23860
rect 14734 23848 14740 23860
rect 13964 23820 14740 23848
rect 13964 23808 13970 23820
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 16022 23808 16028 23860
rect 16080 23848 16086 23860
rect 16301 23851 16359 23857
rect 16301 23848 16313 23851
rect 16080 23820 16313 23848
rect 16080 23808 16086 23820
rect 16301 23817 16313 23820
rect 16347 23817 16359 23851
rect 16301 23811 16359 23817
rect 21545 23851 21603 23857
rect 21545 23817 21557 23851
rect 21591 23848 21603 23851
rect 21634 23848 21640 23860
rect 21591 23820 21640 23848
rect 21591 23817 21603 23820
rect 21545 23811 21603 23817
rect 21634 23808 21640 23820
rect 21692 23808 21698 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23290 23848 23296 23860
rect 22695 23820 23296 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 23474 23848 23480 23860
rect 23435 23820 23480 23848
rect 23474 23808 23480 23820
rect 23532 23808 23538 23860
rect 11330 23712 11336 23724
rect 11291 23684 11336 23712
rect 11330 23672 11336 23684
rect 11388 23672 11394 23724
rect 14826 23672 14832 23724
rect 14884 23712 14890 23724
rect 14921 23715 14979 23721
rect 14921 23712 14933 23715
rect 14884 23684 14933 23712
rect 14884 23672 14890 23684
rect 14921 23681 14933 23684
rect 14967 23681 14979 23715
rect 22370 23712 22376 23724
rect 22283 23684 22376 23712
rect 14921 23675 14979 23681
rect 22370 23672 22376 23684
rect 22428 23712 22434 23724
rect 23382 23712 23388 23724
rect 22428 23684 23388 23712
rect 22428 23672 22434 23684
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 23492 23712 23520 23808
rect 23937 23715 23995 23721
rect 23937 23712 23949 23715
rect 23492 23684 23949 23712
rect 23937 23681 23949 23684
rect 23983 23681 23995 23715
rect 23937 23675 23995 23681
rect 11146 23644 11152 23656
rect 11107 23616 11152 23644
rect 11146 23604 11152 23616
rect 11204 23604 11210 23656
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 12704 23647 12762 23653
rect 12483 23616 12572 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 12544 23576 12572 23616
rect 12704 23613 12716 23647
rect 12750 23644 12762 23647
rect 13078 23644 13084 23656
rect 12750 23616 13084 23644
rect 12750 23613 12762 23616
rect 12704 23607 12762 23613
rect 13078 23604 13084 23616
rect 13136 23604 13142 23656
rect 14844 23576 14872 23672
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 17497 23647 17555 23653
rect 17497 23644 17509 23647
rect 16724 23616 17509 23644
rect 16724 23604 16730 23616
rect 17497 23613 17509 23616
rect 17543 23644 17555 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17543 23616 18061 23644
rect 17543 23613 17555 23616
rect 17497 23607 17555 23613
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 18782 23644 18788 23656
rect 18095 23616 18788 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18782 23604 18788 23616
rect 18840 23604 18846 23656
rect 21361 23647 21419 23653
rect 21361 23613 21373 23647
rect 21407 23644 21419 23647
rect 21450 23644 21456 23656
rect 21407 23616 21456 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 21450 23604 21456 23616
rect 21508 23644 21514 23656
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21508 23616 21925 23644
rect 21508 23604 21514 23616
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 21913 23607 21971 23613
rect 22465 23647 22523 23653
rect 22465 23613 22477 23647
rect 22511 23644 22523 23647
rect 22511 23616 23152 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 15194 23585 15200 23588
rect 15188 23576 15200 23585
rect 11931 23548 14872 23576
rect 15155 23548 15200 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 12728 23520 12756 23548
rect 15188 23539 15200 23548
rect 15194 23536 15200 23539
rect 15252 23536 15258 23588
rect 18230 23536 18236 23588
rect 18288 23585 18294 23588
rect 18288 23579 18352 23585
rect 18288 23545 18306 23579
rect 18340 23545 18352 23579
rect 18288 23539 18352 23545
rect 18288 23536 18294 23539
rect 20990 23536 20996 23588
rect 21048 23576 21054 23588
rect 21085 23579 21143 23585
rect 21085 23576 21097 23579
rect 21048 23548 21097 23576
rect 21048 23536 21054 23548
rect 21085 23545 21097 23548
rect 21131 23576 21143 23579
rect 21634 23576 21640 23588
rect 21131 23548 21640 23576
rect 21131 23545 21143 23548
rect 21085 23539 21143 23545
rect 21634 23536 21640 23548
rect 21692 23536 21698 23588
rect 23124 23520 23152 23616
rect 23566 23604 23572 23656
rect 23624 23644 23630 23656
rect 23753 23647 23811 23653
rect 23753 23644 23765 23647
rect 23624 23616 23765 23644
rect 23624 23604 23630 23616
rect 23753 23613 23765 23616
rect 23799 23613 23811 23647
rect 25038 23644 25044 23656
rect 24999 23616 25044 23644
rect 23753 23607 23811 23613
rect 25038 23604 25044 23616
rect 25096 23644 25102 23656
rect 25593 23647 25651 23653
rect 25593 23644 25605 23647
rect 25096 23616 25605 23644
rect 25096 23604 25102 23616
rect 25593 23613 25605 23616
rect 25639 23613 25651 23647
rect 25593 23607 25651 23613
rect 10686 23508 10692 23520
rect 10599 23480 10692 23508
rect 10686 23468 10692 23480
rect 10744 23508 10750 23520
rect 11238 23508 11244 23520
rect 10744 23480 11244 23508
rect 10744 23468 10750 23480
rect 11238 23468 11244 23480
rect 11296 23468 11302 23520
rect 12253 23511 12311 23517
rect 12253 23477 12265 23511
rect 12299 23508 12311 23511
rect 12618 23508 12624 23520
rect 12299 23480 12624 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 12618 23468 12624 23480
rect 12676 23468 12682 23520
rect 12710 23468 12716 23520
rect 12768 23468 12774 23520
rect 13354 23468 13360 23520
rect 13412 23508 13418 23520
rect 13817 23511 13875 23517
rect 13817 23508 13829 23511
rect 13412 23480 13829 23508
rect 13412 23468 13418 23480
rect 13817 23477 13829 23480
rect 13863 23477 13875 23511
rect 16942 23508 16948 23520
rect 16903 23480 16948 23508
rect 13817 23471 13875 23477
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 17586 23468 17592 23520
rect 17644 23508 17650 23520
rect 17773 23511 17831 23517
rect 17773 23508 17785 23511
rect 17644 23480 17785 23508
rect 17644 23468 17650 23480
rect 17773 23477 17785 23480
rect 17819 23477 17831 23511
rect 17773 23471 17831 23477
rect 19242 23468 19248 23520
rect 19300 23508 19306 23520
rect 19429 23511 19487 23517
rect 19429 23508 19441 23511
rect 19300 23480 19441 23508
rect 19300 23468 19306 23480
rect 19429 23477 19441 23480
rect 19475 23477 19487 23511
rect 19429 23471 19487 23477
rect 20073 23511 20131 23517
rect 20073 23477 20085 23511
rect 20119 23508 20131 23511
rect 20162 23508 20168 23520
rect 20119 23480 20168 23508
rect 20119 23477 20131 23480
rect 20073 23471 20131 23477
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 23106 23508 23112 23520
rect 23067 23480 23112 23508
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 24673 23511 24731 23517
rect 24673 23477 24685 23511
rect 24719 23508 24731 23511
rect 24762 23508 24768 23520
rect 24719 23480 24768 23508
rect 24719 23477 24731 23480
rect 24673 23471 24731 23477
rect 24762 23468 24768 23480
rect 24820 23468 24826 23520
rect 25222 23508 25228 23520
rect 25183 23480 25228 23508
rect 25222 23468 25228 23480
rect 25280 23468 25286 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 10873 23307 10931 23313
rect 10873 23273 10885 23307
rect 10919 23304 10931 23307
rect 10962 23304 10968 23316
rect 10919 23276 10968 23304
rect 10919 23273 10931 23276
rect 10873 23267 10931 23273
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 12526 23304 12532 23316
rect 12487 23276 12532 23304
rect 12526 23264 12532 23276
rect 12584 23304 12590 23316
rect 13078 23304 13084 23316
rect 12584 23276 13084 23304
rect 12584 23264 12590 23276
rect 13078 23264 13084 23276
rect 13136 23264 13142 23316
rect 13262 23264 13268 23316
rect 13320 23304 13326 23316
rect 13449 23307 13507 23313
rect 13449 23304 13461 23307
rect 13320 23276 13461 23304
rect 13320 23264 13326 23276
rect 13449 23273 13461 23276
rect 13495 23273 13507 23307
rect 13449 23267 13507 23273
rect 15565 23307 15623 23313
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 15838 23304 15844 23316
rect 15611 23276 15844 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 15838 23264 15844 23276
rect 15896 23264 15902 23316
rect 15933 23307 15991 23313
rect 15933 23273 15945 23307
rect 15979 23304 15991 23307
rect 16022 23304 16028 23316
rect 15979 23276 16028 23304
rect 15979 23273 15991 23276
rect 15933 23267 15991 23273
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 18969 23307 19027 23313
rect 18969 23304 18981 23307
rect 18012 23276 18981 23304
rect 18012 23264 18018 23276
rect 18969 23273 18981 23276
rect 19015 23273 19027 23307
rect 18969 23267 19027 23273
rect 21085 23307 21143 23313
rect 21085 23273 21097 23307
rect 21131 23304 21143 23307
rect 21358 23304 21364 23316
rect 21131 23276 21364 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 21358 23264 21364 23276
rect 21416 23264 21422 23316
rect 11146 23196 11152 23248
rect 11204 23236 11210 23248
rect 11394 23239 11452 23245
rect 11394 23236 11406 23239
rect 11204 23208 11406 23236
rect 11204 23196 11210 23208
rect 11394 23205 11406 23208
rect 11440 23205 11452 23239
rect 11394 23199 11452 23205
rect 12802 23196 12808 23248
rect 12860 23236 12866 23248
rect 14093 23239 14151 23245
rect 14093 23236 14105 23239
rect 12860 23208 14105 23236
rect 12860 23196 12866 23208
rect 14093 23205 14105 23208
rect 14139 23205 14151 23239
rect 16040 23236 16068 23264
rect 16362 23239 16420 23245
rect 16362 23236 16374 23239
rect 16040 23208 16374 23236
rect 14093 23199 14151 23205
rect 16362 23205 16374 23208
rect 16408 23205 16420 23239
rect 23106 23236 23112 23248
rect 23067 23208 23112 23236
rect 16362 23199 16420 23205
rect 23106 23196 23112 23208
rect 23164 23196 23170 23248
rect 23474 23196 23480 23248
rect 23532 23236 23538 23248
rect 24397 23239 24455 23245
rect 24397 23236 24409 23239
rect 23532 23208 24409 23236
rect 23532 23196 23538 23208
rect 24397 23205 24409 23208
rect 24443 23205 24455 23239
rect 24397 23199 24455 23205
rect 13814 23128 13820 23180
rect 13872 23168 13878 23180
rect 14001 23171 14059 23177
rect 14001 23168 14013 23171
rect 13872 23140 14013 23168
rect 13872 23128 13878 23140
rect 14001 23137 14013 23140
rect 14047 23137 14059 23171
rect 14001 23131 14059 23137
rect 15378 23128 15384 23180
rect 15436 23168 15442 23180
rect 16117 23171 16175 23177
rect 16117 23168 16129 23171
rect 15436 23140 16129 23168
rect 15436 23128 15442 23140
rect 16117 23137 16129 23140
rect 16163 23168 16175 23171
rect 16666 23168 16672 23180
rect 16163 23140 16672 23168
rect 16163 23137 16175 23140
rect 16117 23131 16175 23137
rect 16666 23128 16672 23140
rect 16724 23128 16730 23180
rect 20901 23171 20959 23177
rect 20901 23137 20913 23171
rect 20947 23168 20959 23171
rect 20990 23168 20996 23180
rect 20947 23140 20996 23168
rect 20947 23137 20959 23140
rect 20901 23131 20959 23137
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 22833 23171 22891 23177
rect 22833 23137 22845 23171
rect 22879 23168 22891 23171
rect 23290 23168 23296 23180
rect 22879 23140 23296 23168
rect 22879 23137 22891 23140
rect 22833 23131 22891 23137
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 23934 23128 23940 23180
rect 23992 23168 23998 23180
rect 24121 23171 24179 23177
rect 24121 23168 24133 23171
rect 23992 23140 24133 23168
rect 23992 23128 23998 23140
rect 24121 23137 24133 23140
rect 24167 23137 24179 23171
rect 24121 23131 24179 23137
rect 11054 23060 11060 23112
rect 11112 23100 11118 23112
rect 11149 23103 11207 23109
rect 11149 23100 11161 23103
rect 11112 23072 11161 23100
rect 11112 23060 11118 23072
rect 11149 23069 11161 23072
rect 11195 23069 11207 23103
rect 11149 23063 11207 23069
rect 13262 23060 13268 23112
rect 13320 23100 13326 23112
rect 14185 23103 14243 23109
rect 14185 23100 14197 23103
rect 13320 23072 14197 23100
rect 13320 23060 13326 23072
rect 14185 23069 14197 23072
rect 14231 23100 14243 23103
rect 14734 23100 14740 23112
rect 14231 23072 14740 23100
rect 14231 23069 14243 23072
rect 14185 23063 14243 23069
rect 14734 23060 14740 23072
rect 14792 23100 14798 23112
rect 14921 23103 14979 23109
rect 14921 23100 14933 23103
rect 14792 23072 14933 23100
rect 14792 23060 14798 23072
rect 14921 23069 14933 23072
rect 14967 23100 14979 23103
rect 15194 23100 15200 23112
rect 14967 23072 15200 23100
rect 14967 23069 14979 23072
rect 14921 23063 14979 23069
rect 15194 23060 15200 23072
rect 15252 23060 15258 23112
rect 18506 23060 18512 23112
rect 18564 23100 18570 23112
rect 19061 23103 19119 23109
rect 19061 23100 19073 23103
rect 18564 23072 19073 23100
rect 18564 23060 18570 23072
rect 19061 23069 19073 23072
rect 19107 23069 19119 23103
rect 19061 23063 19119 23069
rect 19153 23103 19211 23109
rect 19153 23069 19165 23103
rect 19199 23069 19211 23103
rect 25406 23100 25412 23112
rect 25367 23072 25412 23100
rect 19153 23063 19211 23069
rect 19168 23032 19196 23063
rect 25406 23060 25412 23072
rect 25464 23060 25470 23112
rect 18248 23004 19196 23032
rect 18248 22976 18276 23004
rect 13173 22967 13231 22973
rect 13173 22933 13185 22967
rect 13219 22964 13231 22967
rect 13354 22964 13360 22976
rect 13219 22936 13360 22964
rect 13219 22933 13231 22936
rect 13173 22927 13231 22933
rect 13354 22924 13360 22936
rect 13412 22924 13418 22976
rect 13630 22964 13636 22976
rect 13591 22936 13636 22964
rect 13630 22924 13636 22936
rect 13688 22924 13694 22976
rect 17494 22964 17500 22976
rect 17455 22936 17500 22964
rect 17494 22924 17500 22936
rect 17552 22964 17558 22976
rect 18049 22967 18107 22973
rect 18049 22964 18061 22967
rect 17552 22936 18061 22964
rect 17552 22924 17558 22936
rect 18049 22933 18061 22936
rect 18095 22964 18107 22967
rect 18230 22964 18236 22976
rect 18095 22936 18236 22964
rect 18095 22933 18107 22936
rect 18049 22927 18107 22933
rect 18230 22924 18236 22936
rect 18288 22924 18294 22976
rect 18598 22964 18604 22976
rect 18559 22936 18604 22964
rect 18598 22924 18604 22936
rect 18656 22924 18662 22976
rect 18782 22924 18788 22976
rect 18840 22964 18846 22976
rect 19705 22967 19763 22973
rect 19705 22964 19717 22967
rect 18840 22936 19717 22964
rect 18840 22924 18846 22936
rect 19705 22933 19717 22936
rect 19751 22964 19763 22967
rect 20530 22964 20536 22976
rect 19751 22936 20536 22964
rect 19751 22933 19763 22936
rect 19705 22927 19763 22933
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 23753 22967 23811 22973
rect 23753 22964 23765 22967
rect 23624 22936 23765 22964
rect 23624 22924 23630 22936
rect 23753 22933 23765 22936
rect 23799 22933 23811 22967
rect 23753 22927 23811 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 12802 22760 12808 22772
rect 12763 22732 12808 22760
rect 12802 22720 12808 22732
rect 12860 22720 12866 22772
rect 13262 22760 13268 22772
rect 13223 22732 13268 22760
rect 13262 22720 13268 22732
rect 13320 22720 13326 22772
rect 14734 22760 14740 22772
rect 14695 22732 14740 22760
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 15933 22763 15991 22769
rect 15933 22729 15945 22763
rect 15979 22760 15991 22763
rect 16022 22760 16028 22772
rect 15979 22732 16028 22760
rect 15979 22729 15991 22732
rect 15933 22723 15991 22729
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18233 22763 18291 22769
rect 18233 22760 18245 22763
rect 18012 22732 18245 22760
rect 18012 22720 18018 22732
rect 18233 22729 18245 22732
rect 18279 22729 18291 22763
rect 21542 22760 21548 22772
rect 21503 22732 21548 22760
rect 18233 22723 18291 22729
rect 21542 22720 21548 22732
rect 21600 22720 21606 22772
rect 23290 22720 23296 22772
rect 23348 22760 23354 22772
rect 23385 22763 23443 22769
rect 23385 22760 23397 22763
rect 23348 22732 23397 22760
rect 23348 22720 23354 22732
rect 23385 22729 23397 22732
rect 23431 22729 23443 22763
rect 23385 22723 23443 22729
rect 17405 22695 17463 22701
rect 17405 22692 17417 22695
rect 16868 22664 17417 22692
rect 11054 22584 11060 22636
rect 11112 22624 11118 22636
rect 11609 22627 11667 22633
rect 11609 22624 11621 22627
rect 11112 22596 11621 22624
rect 11112 22584 11118 22596
rect 11609 22593 11621 22596
rect 11655 22624 11667 22627
rect 12158 22624 12164 22636
rect 11655 22596 12164 22624
rect 11655 22593 11667 22596
rect 11609 22587 11667 22593
rect 12158 22584 12164 22596
rect 12216 22624 12222 22636
rect 12710 22624 12716 22636
rect 12216 22596 12716 22624
rect 12216 22584 12222 22596
rect 12710 22584 12716 22596
rect 12768 22624 12774 22636
rect 13357 22627 13415 22633
rect 13357 22624 13369 22627
rect 12768 22596 13369 22624
rect 12768 22584 12774 22596
rect 13357 22593 13369 22596
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16868 22633 16896 22664
rect 17405 22661 17417 22664
rect 17451 22661 17463 22695
rect 17405 22655 17463 22661
rect 24210 22652 24216 22704
rect 24268 22692 24274 22704
rect 25225 22695 25283 22701
rect 25225 22692 25237 22695
rect 24268 22664 25237 22692
rect 24268 22652 24274 22664
rect 25225 22661 25237 22664
rect 25271 22661 25283 22695
rect 25225 22655 25283 22661
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16632 22596 16865 22624
rect 16632 22584 16638 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 17034 22624 17040 22636
rect 16995 22596 17040 22624
rect 16853 22587 16911 22593
rect 17034 22584 17040 22596
rect 17092 22624 17098 22636
rect 17494 22624 17500 22636
rect 17092 22596 17500 22624
rect 17092 22584 17098 22596
rect 17494 22584 17500 22596
rect 17552 22624 17558 22636
rect 17773 22627 17831 22633
rect 17773 22624 17785 22627
rect 17552 22596 17785 22624
rect 17552 22584 17558 22596
rect 17773 22593 17785 22596
rect 17819 22593 17831 22627
rect 18782 22624 18788 22636
rect 18743 22596 18788 22624
rect 17773 22587 17831 22593
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 24026 22624 24032 22636
rect 23987 22596 24032 22624
rect 24026 22584 24032 22596
rect 24084 22584 24090 22636
rect 16301 22559 16359 22565
rect 16301 22525 16313 22559
rect 16347 22556 16359 22559
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16347 22528 16773 22556
rect 16347 22525 16359 22528
rect 16301 22519 16359 22525
rect 16761 22525 16773 22528
rect 16807 22556 16819 22559
rect 17402 22556 17408 22568
rect 16807 22528 17408 22556
rect 16807 22525 16819 22528
rect 16761 22519 16819 22525
rect 17402 22516 17408 22528
rect 17460 22516 17466 22568
rect 21266 22516 21272 22568
rect 21324 22556 21330 22568
rect 21361 22559 21419 22565
rect 21361 22556 21373 22559
rect 21324 22528 21373 22556
rect 21324 22516 21330 22528
rect 21361 22525 21373 22528
rect 21407 22556 21419 22559
rect 21913 22559 21971 22565
rect 21913 22556 21925 22559
rect 21407 22528 21925 22556
rect 21407 22525 21419 22528
rect 21361 22519 21419 22525
rect 21913 22525 21925 22528
rect 21959 22525 21971 22559
rect 21913 22519 21971 22525
rect 22465 22559 22523 22565
rect 22465 22525 22477 22559
rect 22511 22556 22523 22559
rect 23750 22556 23756 22568
rect 22511 22528 23152 22556
rect 23663 22528 23756 22556
rect 22511 22525 22523 22528
rect 22465 22519 22523 22525
rect 13602 22491 13660 22497
rect 13602 22488 13614 22491
rect 13464 22460 13614 22488
rect 13464 22432 13492 22460
rect 13602 22457 13614 22460
rect 13648 22457 13660 22491
rect 13602 22451 13660 22457
rect 13722 22448 13728 22500
rect 13780 22488 13786 22500
rect 15289 22491 15347 22497
rect 15289 22488 15301 22491
rect 13780 22460 15301 22488
rect 13780 22448 13786 22460
rect 15289 22457 15301 22460
rect 15335 22457 15347 22491
rect 15289 22451 15347 22457
rect 19052 22491 19110 22497
rect 19052 22457 19064 22491
rect 19098 22488 19110 22491
rect 19242 22488 19248 22500
rect 19098 22460 19248 22488
rect 19098 22457 19110 22460
rect 19052 22451 19110 22457
rect 19242 22448 19248 22460
rect 19300 22448 19306 22500
rect 11146 22420 11152 22432
rect 11107 22392 11152 22420
rect 11146 22380 11152 22392
rect 11204 22380 11210 22432
rect 13446 22380 13452 22432
rect 13504 22380 13510 22432
rect 16393 22423 16451 22429
rect 16393 22389 16405 22423
rect 16439 22420 16451 22423
rect 16666 22420 16672 22432
rect 16439 22392 16672 22420
rect 16439 22389 16451 22392
rect 16393 22383 16451 22389
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 18506 22380 18512 22432
rect 18564 22420 18570 22432
rect 18601 22423 18659 22429
rect 18601 22420 18613 22423
rect 18564 22392 18613 22420
rect 18564 22380 18570 22392
rect 18601 22389 18613 22392
rect 18647 22389 18659 22423
rect 18601 22383 18659 22389
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 20165 22423 20223 22429
rect 20165 22420 20177 22423
rect 20128 22392 20177 22420
rect 20128 22380 20134 22392
rect 20165 22389 20177 22392
rect 20211 22389 20223 22423
rect 20990 22420 20996 22432
rect 20951 22392 20996 22420
rect 20165 22383 20223 22389
rect 20990 22380 20996 22392
rect 21048 22380 21054 22432
rect 22646 22420 22652 22432
rect 22607 22392 22652 22420
rect 22646 22380 22652 22392
rect 22704 22380 22710 22432
rect 23124 22429 23152 22528
rect 23750 22516 23756 22528
rect 23808 22556 23814 22568
rect 24489 22559 24547 22565
rect 24489 22556 24501 22559
rect 23808 22528 24501 22556
rect 23808 22516 23814 22528
rect 24489 22525 24501 22528
rect 24535 22525 24547 22559
rect 25038 22556 25044 22568
rect 24999 22528 25044 22556
rect 24489 22519 24547 22525
rect 25038 22516 25044 22528
rect 25096 22556 25102 22568
rect 25593 22559 25651 22565
rect 25593 22556 25605 22559
rect 25096 22528 25605 22556
rect 25096 22516 25102 22528
rect 25593 22525 25605 22528
rect 25639 22525 25651 22559
rect 25593 22519 25651 22525
rect 23109 22423 23167 22429
rect 23109 22389 23121 22423
rect 23155 22420 23167 22423
rect 23198 22420 23204 22432
rect 23155 22392 23204 22420
rect 23155 22389 23167 22392
rect 23109 22383 23167 22389
rect 23198 22380 23204 22392
rect 23256 22380 23262 22432
rect 24026 22380 24032 22432
rect 24084 22420 24090 22432
rect 24857 22423 24915 22429
rect 24857 22420 24869 22423
rect 24084 22392 24869 22420
rect 24084 22380 24090 22392
rect 24857 22389 24869 22392
rect 24903 22389 24915 22423
rect 24857 22383 24915 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 11146 22176 11152 22228
rect 11204 22216 11210 22228
rect 12437 22219 12495 22225
rect 12437 22216 12449 22219
rect 11204 22188 12449 22216
rect 11204 22176 11210 22188
rect 12437 22185 12449 22188
rect 12483 22185 12495 22219
rect 12437 22179 12495 22185
rect 12710 22176 12716 22228
rect 12768 22216 12774 22228
rect 12989 22219 13047 22225
rect 12989 22216 13001 22219
rect 12768 22188 13001 22216
rect 12768 22176 12774 22188
rect 12989 22185 13001 22188
rect 13035 22216 13047 22219
rect 13170 22216 13176 22228
rect 13035 22188 13176 22216
rect 13035 22185 13047 22188
rect 12989 22179 13047 22185
rect 13170 22176 13176 22188
rect 13228 22176 13234 22228
rect 15105 22219 15163 22225
rect 15105 22185 15117 22219
rect 15151 22216 15163 22219
rect 15378 22216 15384 22228
rect 15151 22188 15384 22216
rect 15151 22185 15163 22188
rect 15105 22179 15163 22185
rect 15378 22176 15384 22188
rect 15436 22176 15442 22228
rect 16485 22219 16543 22225
rect 16485 22185 16497 22219
rect 16531 22216 16543 22219
rect 17034 22216 17040 22228
rect 16531 22188 17040 22216
rect 16531 22185 16543 22188
rect 16485 22179 16543 22185
rect 17034 22176 17040 22188
rect 17092 22176 17098 22228
rect 17957 22219 18015 22225
rect 17957 22185 17969 22219
rect 18003 22216 18015 22219
rect 18598 22216 18604 22228
rect 18003 22188 18604 22216
rect 18003 22185 18015 22188
rect 17957 22179 18015 22185
rect 13909 22151 13967 22157
rect 13909 22148 13921 22151
rect 13832 22120 13921 22148
rect 1394 22040 1400 22092
rect 1452 22080 1458 22092
rect 2314 22080 2320 22092
rect 1452 22052 2320 22080
rect 1452 22040 1458 22052
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 11054 22080 11060 22092
rect 10100 22052 11060 22080
rect 10100 22040 10106 22052
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11324 22083 11382 22089
rect 11324 22049 11336 22083
rect 11370 22080 11382 22083
rect 11790 22080 11796 22092
rect 11370 22052 11796 22080
rect 11370 22049 11382 22052
rect 11324 22043 11382 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 13354 22040 13360 22092
rect 13412 22080 13418 22092
rect 13832 22080 13860 22120
rect 13909 22117 13921 22120
rect 13955 22117 13967 22151
rect 13909 22111 13967 22117
rect 16577 22151 16635 22157
rect 16577 22117 16589 22151
rect 16623 22148 16635 22151
rect 16942 22148 16948 22160
rect 16623 22120 16948 22148
rect 16623 22117 16635 22120
rect 16577 22111 16635 22117
rect 16942 22108 16948 22120
rect 17000 22108 17006 22160
rect 15286 22080 15292 22092
rect 13412 22052 13860 22080
rect 15247 22052 15292 22080
rect 13412 22040 13418 22052
rect 15286 22040 15292 22052
rect 15344 22040 15350 22092
rect 17497 22083 17555 22089
rect 17497 22049 17509 22083
rect 17543 22080 17555 22083
rect 17972 22080 18000 22179
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 18877 22219 18935 22225
rect 18877 22185 18889 22219
rect 18923 22216 18935 22219
rect 19242 22216 19248 22228
rect 18923 22188 19248 22216
rect 18923 22185 18935 22188
rect 18877 22179 18935 22185
rect 18892 22148 18920 22179
rect 19242 22176 19248 22188
rect 19300 22176 19306 22228
rect 22738 22216 22744 22228
rect 22699 22188 22744 22216
rect 22738 22176 22744 22188
rect 22796 22176 22802 22228
rect 20530 22148 20536 22160
rect 17543 22052 18000 22080
rect 18248 22120 18920 22148
rect 20491 22120 20536 22148
rect 17543 22049 17555 22052
rect 17497 22043 17555 22049
rect 13998 22012 14004 22024
rect 13959 21984 14004 22012
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 15562 22012 15568 22024
rect 15523 21984 15568 22012
rect 14093 21975 14151 21981
rect 13541 21947 13599 21953
rect 13541 21913 13553 21947
rect 13587 21944 13599 21947
rect 13722 21944 13728 21956
rect 13587 21916 13728 21944
rect 13587 21913 13599 21916
rect 13541 21907 13599 21913
rect 13722 21904 13728 21916
rect 13780 21904 13786 21956
rect 9309 21879 9367 21885
rect 9309 21845 9321 21879
rect 9355 21876 9367 21879
rect 9950 21876 9956 21888
rect 9355 21848 9956 21876
rect 9355 21845 9367 21848
rect 9309 21839 9367 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 10873 21879 10931 21885
rect 10873 21845 10885 21879
rect 10919 21876 10931 21879
rect 11238 21876 11244 21888
rect 10919 21848 11244 21876
rect 10919 21845 10931 21848
rect 10873 21839 10931 21845
rect 11238 21836 11244 21848
rect 11296 21836 11302 21888
rect 13446 21876 13452 21888
rect 13407 21848 13452 21876
rect 13446 21836 13452 21848
rect 13504 21876 13510 21888
rect 14108 21876 14136 21975
rect 15562 21972 15568 21984
rect 15620 21972 15626 22024
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 18049 22015 18107 22021
rect 18049 22012 18061 22015
rect 16724 21984 18061 22012
rect 16724 21972 16730 21984
rect 18049 21981 18061 21984
rect 18095 21981 18107 22015
rect 18049 21975 18107 21981
rect 18138 21972 18144 22024
rect 18196 22012 18202 22024
rect 18248 22012 18276 22120
rect 20530 22108 20536 22120
rect 20588 22108 20594 22160
rect 19153 22083 19211 22089
rect 19153 22049 19165 22083
rect 19199 22049 19211 22083
rect 19153 22043 19211 22049
rect 19429 22083 19487 22089
rect 19429 22049 19441 22083
rect 19475 22080 19487 22083
rect 20898 22080 20904 22092
rect 19475 22052 20904 22080
rect 19475 22049 19487 22052
rect 19429 22043 19487 22049
rect 18196 21984 18276 22012
rect 18196 21972 18202 21984
rect 15470 21904 15476 21956
rect 15528 21944 15534 21956
rect 15746 21944 15752 21956
rect 15528 21916 15752 21944
rect 15528 21904 15534 21916
rect 15746 21904 15752 21916
rect 15804 21904 15810 21956
rect 17589 21947 17647 21953
rect 17589 21913 17601 21947
rect 17635 21944 17647 21947
rect 19168 21944 19196 22043
rect 20898 22040 20904 22052
rect 20956 22040 20962 22092
rect 21266 22080 21272 22092
rect 21227 22052 21272 22080
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 23934 22040 23940 22092
rect 23992 22080 23998 22092
rect 24581 22083 24639 22089
rect 24581 22080 24593 22083
rect 23992 22052 24593 22080
rect 23992 22040 23998 22052
rect 24581 22049 24593 22052
rect 24627 22049 24639 22083
rect 24581 22043 24639 22049
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 22830 22012 22836 22024
rect 22520 21984 22836 22012
rect 22520 21972 22526 21984
rect 22830 21972 22836 21984
rect 22888 21972 22894 22024
rect 23014 22012 23020 22024
rect 22975 21984 23020 22012
rect 23014 21972 23020 21984
rect 23072 21972 23078 22024
rect 19426 21944 19432 21956
rect 17635 21916 19432 21944
rect 17635 21913 17647 21916
rect 17589 21907 17647 21913
rect 19426 21904 19432 21916
rect 19484 21904 19490 21956
rect 21450 21944 21456 21956
rect 21411 21916 21456 21944
rect 21450 21904 21456 21916
rect 21508 21904 21514 21956
rect 14642 21876 14648 21888
rect 13504 21848 14136 21876
rect 14603 21848 14648 21876
rect 13504 21836 13510 21848
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 14826 21836 14832 21888
rect 14884 21876 14890 21888
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 14884 21848 16037 21876
rect 14884 21836 14890 21848
rect 16025 21845 16037 21848
rect 16071 21876 16083 21879
rect 16482 21876 16488 21888
rect 16071 21848 16488 21876
rect 16071 21845 16083 21848
rect 16025 21839 16083 21845
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 17126 21876 17132 21888
rect 17087 21848 17132 21876
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 22002 21876 22008 21888
rect 21963 21848 22008 21876
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 22373 21879 22431 21885
rect 22373 21845 22385 21879
rect 22419 21876 22431 21879
rect 22646 21876 22652 21888
rect 22419 21848 22652 21876
rect 22419 21845 22431 21848
rect 22373 21839 22431 21845
rect 22646 21836 22652 21848
rect 22704 21836 22710 21888
rect 24670 21836 24676 21888
rect 24728 21876 24734 21888
rect 24765 21879 24823 21885
rect 24765 21876 24777 21879
rect 24728 21848 24777 21876
rect 24728 21836 24734 21848
rect 24765 21845 24777 21848
rect 24811 21845 24823 21879
rect 24765 21839 24823 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 8386 21632 8392 21684
rect 8444 21672 8450 21684
rect 9033 21675 9091 21681
rect 9033 21672 9045 21675
rect 8444 21644 9045 21672
rect 8444 21632 8450 21644
rect 9033 21641 9045 21644
rect 9079 21672 9091 21675
rect 11790 21672 11796 21684
rect 9079 21644 9628 21672
rect 11751 21644 11796 21672
rect 9079 21641 9091 21644
rect 9033 21635 9091 21641
rect 9600 21477 9628 21644
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12158 21672 12164 21684
rect 12119 21644 12164 21672
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 13354 21672 13360 21684
rect 13315 21644 13360 21672
rect 13354 21632 13360 21644
rect 13412 21672 13418 21684
rect 13412 21644 13492 21672
rect 13412 21632 13418 21644
rect 9861 21539 9919 21545
rect 9861 21505 9873 21539
rect 9907 21536 9919 21539
rect 9950 21536 9956 21548
rect 9907 21508 9956 21536
rect 9907 21505 9919 21508
rect 9861 21499 9919 21505
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21536 10747 21539
rect 11146 21536 11152 21548
rect 10735 21508 11152 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 11146 21496 11152 21508
rect 11204 21536 11210 21548
rect 13464 21545 13492 21644
rect 13814 21632 13820 21684
rect 13872 21672 13878 21684
rect 14277 21675 14335 21681
rect 14277 21672 14289 21675
rect 13872 21644 14289 21672
rect 13872 21632 13878 21644
rect 14277 21641 14289 21644
rect 14323 21641 14335 21675
rect 14277 21635 14335 21641
rect 14461 21675 14519 21681
rect 14461 21641 14473 21675
rect 14507 21672 14519 21675
rect 14826 21672 14832 21684
rect 14507 21644 14832 21672
rect 14507 21641 14519 21644
rect 14461 21635 14519 21641
rect 11333 21539 11391 21545
rect 11333 21536 11345 21539
rect 11204 21508 11345 21536
rect 11204 21496 11210 21508
rect 11333 21505 11345 21508
rect 11379 21505 11391 21539
rect 11333 21499 11391 21505
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21505 13507 21539
rect 14292 21536 14320 21635
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 15286 21632 15292 21684
rect 15344 21672 15350 21684
rect 15473 21675 15531 21681
rect 15473 21672 15485 21675
rect 15344 21644 15485 21672
rect 15344 21632 15350 21644
rect 15473 21641 15485 21644
rect 15519 21641 15531 21675
rect 15473 21635 15531 21641
rect 16666 21632 16672 21684
rect 16724 21672 16730 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16724 21644 17049 21672
rect 16724 21632 16730 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 17037 21635 17095 21641
rect 17126 21632 17132 21684
rect 17184 21672 17190 21684
rect 18049 21675 18107 21681
rect 18049 21672 18061 21675
rect 17184 21644 18061 21672
rect 17184 21632 17190 21644
rect 18049 21641 18061 21644
rect 18095 21641 18107 21675
rect 19426 21672 19432 21684
rect 19387 21644 19432 21672
rect 18049 21635 18107 21641
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 22833 21675 22891 21681
rect 22833 21672 22845 21675
rect 22796 21644 22845 21672
rect 22796 21632 22802 21644
rect 22833 21641 22845 21644
rect 22879 21641 22891 21675
rect 22833 21635 22891 21641
rect 23014 21632 23020 21684
rect 23072 21672 23078 21684
rect 23201 21675 23259 21681
rect 23201 21672 23213 21675
rect 23072 21644 23213 21672
rect 23072 21632 23078 21644
rect 23201 21641 23213 21644
rect 23247 21641 23259 21675
rect 23201 21635 23259 21641
rect 23934 21632 23940 21684
rect 23992 21672 23998 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 23992 21644 25053 21672
rect 23992 21632 23998 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 14642 21564 14648 21616
rect 14700 21604 14706 21616
rect 14700 21576 15056 21604
rect 14700 21564 14706 21576
rect 15028 21545 15056 21576
rect 15930 21564 15936 21616
rect 15988 21604 15994 21616
rect 15988 21576 16620 21604
rect 15988 21564 15994 21576
rect 14921 21539 14979 21545
rect 14921 21536 14933 21539
rect 14292 21508 14933 21536
rect 13449 21499 13507 21505
rect 14921 21505 14933 21508
rect 14967 21505 14979 21539
rect 14921 21499 14979 21505
rect 15013 21539 15071 21545
rect 15013 21505 15025 21539
rect 15059 21536 15071 21539
rect 15378 21536 15384 21548
rect 15059 21508 15384 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 15378 21496 15384 21508
rect 15436 21496 15442 21548
rect 16482 21536 16488 21548
rect 16443 21508 16488 21536
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 16592 21545 16620 21576
rect 16577 21539 16635 21545
rect 16577 21505 16589 21539
rect 16623 21505 16635 21539
rect 18598 21536 18604 21548
rect 18559 21508 18604 21536
rect 16577 21499 16635 21505
rect 18598 21496 18604 21508
rect 18656 21536 18662 21548
rect 19061 21539 19119 21545
rect 19061 21536 19073 21539
rect 18656 21508 19073 21536
rect 18656 21496 18662 21508
rect 19061 21505 19073 21508
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 9585 21471 9643 21477
rect 9585 21437 9597 21471
rect 9631 21437 9643 21471
rect 9585 21431 9643 21437
rect 16393 21471 16451 21477
rect 16393 21437 16405 21471
rect 16439 21468 16451 21471
rect 17126 21468 17132 21480
rect 16439 21440 17132 21468
rect 16439 21437 16451 21440
rect 16393 21431 16451 21437
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 20530 21468 20536 21480
rect 20443 21440 20536 21468
rect 20530 21428 20536 21440
rect 20588 21468 20594 21480
rect 22002 21468 22008 21480
rect 20588 21440 22008 21468
rect 20588 21428 20594 21440
rect 22002 21428 22008 21440
rect 22060 21428 22066 21480
rect 24305 21471 24363 21477
rect 24305 21468 24317 21471
rect 24136 21440 24317 21468
rect 10321 21403 10379 21409
rect 10321 21369 10333 21403
rect 10367 21400 10379 21403
rect 10686 21400 10692 21412
rect 10367 21372 10692 21400
rect 10367 21369 10379 21372
rect 10321 21363 10379 21369
rect 10686 21360 10692 21372
rect 10744 21400 10750 21412
rect 11149 21403 11207 21409
rect 11149 21400 11161 21403
rect 10744 21372 11161 21400
rect 10744 21360 10750 21372
rect 11149 21369 11161 21372
rect 11195 21369 11207 21403
rect 15930 21400 15936 21412
rect 15891 21372 15936 21400
rect 11149 21363 11207 21369
rect 15930 21360 15936 21372
rect 15988 21360 15994 21412
rect 16574 21360 16580 21412
rect 16632 21400 16638 21412
rect 17773 21403 17831 21409
rect 17773 21400 17785 21403
rect 16632 21372 17785 21400
rect 16632 21360 16638 21372
rect 17773 21369 17785 21372
rect 17819 21400 17831 21403
rect 18509 21403 18567 21409
rect 18509 21400 18521 21403
rect 17819 21372 18521 21400
rect 17819 21369 17831 21372
rect 17773 21363 17831 21369
rect 18509 21369 18521 21372
rect 18555 21369 18567 21403
rect 20778 21403 20836 21409
rect 20778 21400 20790 21403
rect 18509 21363 18567 21369
rect 20456 21372 20790 21400
rect 20456 21344 20484 21372
rect 20778 21369 20790 21372
rect 20824 21369 20836 21403
rect 23014 21400 23020 21412
rect 20778 21363 20836 21369
rect 22296 21372 23020 21400
rect 22296 21344 22324 21372
rect 23014 21360 23020 21372
rect 23072 21360 23078 21412
rect 9214 21332 9220 21344
rect 9175 21304 9220 21332
rect 9214 21292 9220 21304
rect 9272 21292 9278 21344
rect 9306 21292 9312 21344
rect 9364 21332 9370 21344
rect 9677 21335 9735 21341
rect 9677 21332 9689 21335
rect 9364 21304 9689 21332
rect 9364 21292 9370 21304
rect 9677 21301 9689 21304
rect 9723 21301 9735 21335
rect 9677 21295 9735 21301
rect 10781 21335 10839 21341
rect 10781 21301 10793 21335
rect 10827 21332 10839 21335
rect 10962 21332 10968 21344
rect 10827 21304 10968 21332
rect 10827 21301 10839 21304
rect 10781 21295 10839 21301
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11238 21332 11244 21344
rect 11199 21304 11244 21332
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 12437 21335 12495 21341
rect 12437 21301 12449 21335
rect 12483 21332 12495 21335
rect 12526 21332 12532 21344
rect 12483 21304 12532 21332
rect 12483 21301 12495 21304
rect 12437 21295 12495 21301
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 13998 21332 14004 21344
rect 13959 21304 14004 21332
rect 13998 21292 14004 21304
rect 14056 21292 14062 21344
rect 14642 21292 14648 21344
rect 14700 21332 14706 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 14700 21304 14841 21332
rect 14700 21292 14706 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 16022 21332 16028 21344
rect 15983 21304 16028 21332
rect 14829 21295 14887 21301
rect 16022 21292 16028 21304
rect 16080 21292 16086 21344
rect 17402 21332 17408 21344
rect 17363 21304 17408 21332
rect 17402 21292 17408 21304
rect 17460 21332 17466 21344
rect 18417 21335 18475 21341
rect 18417 21332 18429 21335
rect 17460 21304 18429 21332
rect 17460 21292 17466 21304
rect 18417 21301 18429 21304
rect 18463 21301 18475 21335
rect 18417 21295 18475 21301
rect 19518 21292 19524 21344
rect 19576 21332 19582 21344
rect 19797 21335 19855 21341
rect 19797 21332 19809 21335
rect 19576 21304 19809 21332
rect 19576 21292 19582 21304
rect 19797 21301 19809 21304
rect 19843 21301 19855 21335
rect 20438 21332 20444 21344
rect 20399 21304 20444 21332
rect 19797 21295 19855 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21913 21335 21971 21341
rect 21913 21301 21925 21335
rect 21959 21332 21971 21335
rect 22278 21332 22284 21344
rect 21959 21304 22284 21332
rect 21959 21301 21971 21304
rect 21913 21295 21971 21301
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 22462 21332 22468 21344
rect 22423 21304 22468 21332
rect 22462 21292 22468 21304
rect 22520 21292 22526 21344
rect 23934 21292 23940 21344
rect 23992 21332 23998 21344
rect 24136 21341 24164 21440
rect 24305 21437 24317 21440
rect 24351 21437 24363 21471
rect 24305 21431 24363 21437
rect 24578 21400 24584 21412
rect 24539 21372 24584 21400
rect 24578 21360 24584 21372
rect 24636 21360 24642 21412
rect 24121 21335 24179 21341
rect 24121 21332 24133 21335
rect 23992 21304 24133 21332
rect 23992 21292 23998 21304
rect 24121 21301 24133 21304
rect 24167 21301 24179 21335
rect 24121 21295 24179 21301
rect 24854 21292 24860 21344
rect 24912 21332 24918 21344
rect 25593 21335 25651 21341
rect 25593 21332 25605 21335
rect 24912 21304 25605 21332
rect 24912 21292 24918 21304
rect 25593 21301 25605 21304
rect 25639 21301 25651 21335
rect 25593 21295 25651 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 11238 21088 11244 21140
rect 11296 21128 11302 21140
rect 12529 21131 12587 21137
rect 12529 21128 12541 21131
rect 11296 21100 12541 21128
rect 11296 21088 11302 21100
rect 12529 21097 12541 21100
rect 12575 21097 12587 21131
rect 12529 21091 12587 21097
rect 13446 21088 13452 21140
rect 13504 21128 13510 21140
rect 13541 21131 13599 21137
rect 13541 21128 13553 21131
rect 13504 21100 13553 21128
rect 13504 21088 13510 21100
rect 13541 21097 13553 21100
rect 13587 21097 13599 21131
rect 13541 21091 13599 21097
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 16850 21128 16856 21140
rect 16080 21100 16856 21128
rect 16080 21088 16086 21100
rect 16850 21088 16856 21100
rect 16908 21128 16914 21140
rect 17221 21131 17279 21137
rect 17221 21128 17233 21131
rect 16908 21100 17233 21128
rect 16908 21088 16914 21100
rect 17221 21097 17233 21100
rect 17267 21097 17279 21131
rect 17221 21091 17279 21097
rect 17681 21131 17739 21137
rect 17681 21097 17693 21131
rect 17727 21128 17739 21131
rect 18138 21128 18144 21140
rect 17727 21100 18144 21128
rect 17727 21097 17739 21100
rect 17681 21091 17739 21097
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 19889 21131 19947 21137
rect 19889 21097 19901 21131
rect 19935 21128 19947 21131
rect 19978 21128 19984 21140
rect 19935 21100 19984 21128
rect 19935 21097 19947 21100
rect 19889 21091 19947 21097
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 21266 21088 21272 21140
rect 21324 21128 21330 21140
rect 21818 21128 21824 21140
rect 21324 21100 21824 21128
rect 21324 21088 21330 21100
rect 21818 21088 21824 21100
rect 21876 21088 21882 21140
rect 13170 21020 13176 21072
rect 13228 21060 13234 21072
rect 13906 21060 13912 21072
rect 13228 21032 13912 21060
rect 13228 21020 13234 21032
rect 13906 21020 13912 21032
rect 13964 21060 13970 21072
rect 13964 21032 15332 21060
rect 13964 21020 13970 21032
rect 9950 20952 9956 21004
rect 10008 20992 10014 21004
rect 10301 20995 10359 21001
rect 10301 20992 10313 20995
rect 10008 20964 10313 20992
rect 10008 20952 10014 20964
rect 10301 20961 10313 20964
rect 10347 20961 10359 20995
rect 10301 20955 10359 20961
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 12897 20995 12955 21001
rect 12492 20964 12537 20992
rect 12492 20952 12498 20964
rect 12897 20961 12909 20995
rect 12943 20992 12955 20995
rect 13354 20992 13360 21004
rect 12943 20964 13360 20992
rect 12943 20961 12955 20964
rect 12897 20955 12955 20961
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 15304 21001 15332 21032
rect 15378 21020 15384 21072
rect 15436 21060 15442 21072
rect 22278 21069 22284 21072
rect 15534 21063 15592 21069
rect 15534 21060 15546 21063
rect 15436 21032 15546 21060
rect 15436 21020 15442 21032
rect 15534 21029 15546 21032
rect 15580 21029 15592 21063
rect 22272 21060 22284 21069
rect 22239 21032 22284 21060
rect 15534 21023 15592 21029
rect 22272 21023 22284 21032
rect 22278 21020 22284 21023
rect 22336 21020 22342 21072
rect 24762 21060 24768 21072
rect 24723 21032 24768 21060
rect 24762 21020 24768 21032
rect 24820 21020 24826 21072
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20961 15347 20995
rect 18138 20992 18144 21004
rect 18099 20964 18144 20992
rect 15289 20955 15347 20961
rect 18138 20952 18144 20964
rect 18196 20952 18202 21004
rect 19518 20992 19524 21004
rect 19479 20964 19524 20992
rect 19518 20952 19524 20964
rect 19576 20952 19582 21004
rect 19705 20995 19763 21001
rect 19705 20961 19717 20995
rect 19751 20992 19763 20995
rect 20346 20992 20352 21004
rect 19751 20964 20352 20992
rect 19751 20961 19763 20964
rect 19705 20955 19763 20961
rect 20346 20952 20352 20964
rect 20404 20952 20410 21004
rect 20898 20992 20904 21004
rect 20859 20964 20904 20992
rect 20898 20952 20904 20964
rect 20956 20992 20962 21004
rect 21453 20995 21511 21001
rect 21453 20992 21465 20995
rect 20956 20964 21465 20992
rect 20956 20952 20962 20964
rect 21453 20961 21465 20964
rect 21499 20961 21511 20995
rect 22002 20992 22008 21004
rect 21963 20964 22008 20992
rect 21453 20955 21511 20961
rect 22002 20952 22008 20964
rect 22060 20952 22066 21004
rect 24118 20952 24124 21004
rect 24176 20992 24182 21004
rect 24489 20995 24547 21001
rect 24489 20992 24501 20995
rect 24176 20964 24501 20992
rect 24176 20952 24182 20964
rect 24489 20961 24501 20964
rect 24535 20961 24547 20995
rect 24489 20955 24547 20961
rect 10042 20924 10048 20936
rect 10003 20896 10048 20924
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 12452 20924 12480 20952
rect 12989 20927 13047 20933
rect 12989 20924 13001 20927
rect 12452 20896 13001 20924
rect 12989 20893 13001 20896
rect 13035 20893 13047 20927
rect 12989 20887 13047 20893
rect 13081 20927 13139 20933
rect 13081 20893 13093 20927
rect 13127 20893 13139 20927
rect 13081 20887 13139 20893
rect 11425 20859 11483 20865
rect 11425 20825 11437 20859
rect 11471 20856 11483 20859
rect 11790 20856 11796 20868
rect 11471 20828 11796 20856
rect 11471 20825 11483 20828
rect 11425 20819 11483 20825
rect 11790 20816 11796 20828
rect 11848 20856 11854 20868
rect 13096 20856 13124 20887
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 18012 20896 18245 20924
rect 18012 20884 18018 20896
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 18325 20927 18383 20933
rect 18325 20893 18337 20927
rect 18371 20893 18383 20927
rect 18325 20887 18383 20893
rect 18340 20856 18368 20887
rect 23658 20856 23664 20868
rect 11848 20828 13124 20856
rect 16684 20828 18368 20856
rect 23216 20828 23664 20856
rect 11848 20816 11854 20828
rect 7650 20788 7656 20800
rect 7611 20760 7656 20788
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 9306 20788 9312 20800
rect 9267 20760 9312 20788
rect 9306 20748 9312 20760
rect 9364 20748 9370 20800
rect 14553 20791 14611 20797
rect 14553 20757 14565 20791
rect 14599 20788 14611 20791
rect 14642 20788 14648 20800
rect 14599 20760 14648 20788
rect 14599 20757 14611 20760
rect 14553 20751 14611 20757
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 16684 20797 16712 20828
rect 16669 20791 16727 20797
rect 16669 20788 16681 20791
rect 15988 20760 16681 20788
rect 15988 20748 15994 20760
rect 16669 20757 16681 20760
rect 16715 20757 16727 20791
rect 16669 20751 16727 20757
rect 16758 20748 16764 20800
rect 16816 20788 16822 20800
rect 17773 20791 17831 20797
rect 17773 20788 17785 20791
rect 16816 20760 17785 20788
rect 16816 20748 16822 20760
rect 17773 20757 17785 20760
rect 17819 20757 17831 20791
rect 18782 20788 18788 20800
rect 18743 20760 18788 20788
rect 17773 20751 17831 20757
rect 18782 20748 18788 20760
rect 18840 20748 18846 20800
rect 19150 20788 19156 20800
rect 19111 20760 19156 20788
rect 19150 20748 19156 20760
rect 19208 20748 19214 20800
rect 19334 20788 19340 20800
rect 19295 20760 19340 20788
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 21082 20788 21088 20800
rect 21043 20760 21088 20788
rect 21082 20748 21088 20760
rect 21140 20748 21146 20800
rect 22002 20748 22008 20800
rect 22060 20788 22066 20800
rect 23216 20788 23244 20828
rect 23658 20816 23664 20828
rect 23716 20856 23722 20868
rect 23937 20859 23995 20865
rect 23937 20856 23949 20859
rect 23716 20828 23949 20856
rect 23716 20816 23722 20828
rect 23937 20825 23949 20828
rect 23983 20825 23995 20859
rect 23937 20819 23995 20825
rect 22060 20760 23244 20788
rect 22060 20748 22066 20760
rect 23290 20748 23296 20800
rect 23348 20788 23354 20800
rect 23385 20791 23443 20797
rect 23385 20788 23397 20791
rect 23348 20760 23397 20788
rect 23348 20748 23354 20760
rect 23385 20757 23397 20760
rect 23431 20757 23443 20791
rect 23385 20751 23443 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 9585 20587 9643 20593
rect 9585 20553 9597 20587
rect 9631 20584 9643 20587
rect 9674 20584 9680 20596
rect 9631 20556 9680 20584
rect 9631 20553 9643 20556
rect 9585 20547 9643 20553
rect 9674 20544 9680 20556
rect 9732 20584 9738 20596
rect 10042 20584 10048 20596
rect 9732 20556 10048 20584
rect 9732 20544 9738 20556
rect 10042 20544 10048 20556
rect 10100 20544 10106 20596
rect 10686 20544 10692 20596
rect 10744 20584 10750 20596
rect 10781 20587 10839 20593
rect 10781 20584 10793 20587
rect 10744 20556 10793 20584
rect 10744 20544 10750 20556
rect 10781 20553 10793 20556
rect 10827 20553 10839 20587
rect 11790 20584 11796 20596
rect 11751 20556 11796 20584
rect 10781 20547 10839 20553
rect 11790 20544 11796 20556
rect 11848 20584 11854 20596
rect 12161 20587 12219 20593
rect 12161 20584 12173 20587
rect 11848 20556 12173 20584
rect 11848 20544 11854 20556
rect 12161 20553 12173 20556
rect 12207 20553 12219 20587
rect 12161 20547 12219 20553
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 15378 20584 15384 20596
rect 15335 20556 15384 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 15378 20544 15384 20556
rect 15436 20584 15442 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 15436 20556 15853 20584
rect 15436 20544 15442 20556
rect 15841 20553 15853 20556
rect 15887 20584 15899 20587
rect 16022 20584 16028 20596
rect 15887 20556 16028 20584
rect 15887 20553 15899 20556
rect 15841 20547 15899 20553
rect 16022 20544 16028 20556
rect 16080 20544 16086 20596
rect 16206 20544 16212 20596
rect 16264 20584 16270 20596
rect 17497 20587 17555 20593
rect 16264 20556 16896 20584
rect 16264 20544 16270 20556
rect 11425 20451 11483 20457
rect 11425 20417 11437 20451
rect 11471 20448 11483 20451
rect 11808 20448 11836 20544
rect 16393 20519 16451 20525
rect 16393 20485 16405 20519
rect 16439 20485 16451 20519
rect 16868 20516 16896 20556
rect 17497 20553 17509 20587
rect 17543 20584 17555 20587
rect 17862 20584 17868 20596
rect 17543 20556 17868 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 23014 20584 23020 20596
rect 22975 20556 23020 20584
rect 23014 20544 23020 20556
rect 23072 20544 23078 20596
rect 16868 20488 16988 20516
rect 16393 20479 16451 20485
rect 12710 20448 12716 20460
rect 11471 20420 11836 20448
rect 12671 20420 12716 20448
rect 11471 20417 11483 20420
rect 11425 20411 11483 20417
rect 12710 20408 12716 20420
rect 12768 20408 12774 20460
rect 13906 20448 13912 20460
rect 13867 20420 13912 20448
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 7561 20383 7619 20389
rect 7561 20349 7573 20383
rect 7607 20380 7619 20383
rect 7650 20380 7656 20392
rect 7607 20352 7656 20380
rect 7607 20349 7619 20352
rect 7561 20343 7619 20349
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 12158 20340 12164 20392
rect 12216 20380 12222 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12216 20352 12449 20380
rect 12216 20340 12222 20352
rect 12437 20349 12449 20352
rect 12483 20349 12495 20383
rect 16408 20380 16436 20479
rect 16850 20448 16856 20460
rect 16811 20420 16856 20448
rect 16850 20408 16856 20420
rect 16908 20408 16914 20460
rect 16960 20457 16988 20488
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20448 17003 20451
rect 17218 20448 17224 20460
rect 16991 20420 17224 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 21545 20451 21603 20457
rect 21545 20417 21557 20451
rect 21591 20448 21603 20451
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 21591 20420 22661 20448
rect 21591 20417 21603 20420
rect 21545 20411 21603 20417
rect 22649 20417 22661 20420
rect 22695 20448 22707 20451
rect 23032 20448 23060 20544
rect 23658 20448 23664 20460
rect 22695 20420 23060 20448
rect 23619 20420 23664 20448
rect 22695 20417 22707 20420
rect 22649 20411 22707 20417
rect 23658 20408 23664 20420
rect 23716 20408 23722 20460
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 16408 20352 18061 20380
rect 12437 20343 12495 20349
rect 18049 20349 18061 20352
rect 18095 20380 18107 20383
rect 18782 20380 18788 20392
rect 18095 20352 18788 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 19392 20352 19533 20380
rect 19392 20340 19398 20352
rect 19521 20349 19533 20352
rect 19567 20380 19579 20383
rect 20530 20380 20536 20392
rect 19567 20352 20536 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 7834 20321 7840 20324
rect 7469 20315 7527 20321
rect 7469 20281 7481 20315
rect 7515 20312 7527 20315
rect 7828 20312 7840 20321
rect 7515 20284 7840 20312
rect 7515 20281 7527 20284
rect 7469 20275 7527 20281
rect 7828 20275 7840 20284
rect 7834 20272 7840 20275
rect 7892 20272 7898 20324
rect 10321 20315 10379 20321
rect 10321 20281 10333 20315
rect 10367 20312 10379 20315
rect 11149 20315 11207 20321
rect 11149 20312 11161 20315
rect 10367 20284 11161 20312
rect 10367 20281 10379 20284
rect 10321 20275 10379 20281
rect 11149 20281 11161 20284
rect 11195 20312 11207 20315
rect 12342 20312 12348 20324
rect 11195 20284 12348 20312
rect 11195 20281 11207 20284
rect 11149 20275 11207 20281
rect 12342 20272 12348 20284
rect 12400 20272 12406 20324
rect 14182 20321 14188 20324
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20312 13875 20315
rect 14165 20315 14188 20321
rect 14165 20312 14177 20315
rect 13863 20284 14177 20312
rect 13863 20281 13875 20284
rect 13817 20275 13875 20281
rect 14165 20281 14177 20284
rect 14165 20275 14188 20281
rect 14182 20272 14188 20275
rect 14240 20272 14246 20324
rect 16206 20312 16212 20324
rect 16167 20284 16212 20312
rect 16206 20272 16212 20284
rect 16264 20272 16270 20324
rect 16758 20312 16764 20324
rect 16719 20284 16764 20312
rect 16758 20272 16764 20284
rect 16816 20272 16822 20324
rect 18322 20312 18328 20324
rect 18283 20284 18328 20312
rect 18322 20272 18328 20284
rect 18380 20272 18386 20324
rect 19429 20315 19487 20321
rect 19429 20281 19441 20315
rect 19475 20312 19487 20315
rect 19788 20315 19846 20321
rect 19788 20312 19800 20315
rect 19475 20284 19800 20312
rect 19475 20281 19487 20284
rect 19429 20275 19487 20281
rect 19788 20281 19800 20284
rect 19834 20312 19846 20315
rect 20070 20312 20076 20324
rect 19834 20284 20076 20312
rect 19834 20281 19846 20284
rect 19788 20275 19846 20281
rect 20070 20272 20076 20284
rect 20128 20272 20134 20324
rect 20806 20272 20812 20324
rect 20864 20312 20870 20324
rect 21821 20315 21879 20321
rect 21821 20312 21833 20315
rect 20864 20284 21833 20312
rect 20864 20272 20870 20284
rect 21821 20281 21833 20284
rect 21867 20312 21879 20315
rect 22465 20315 22523 20321
rect 22465 20312 22477 20315
rect 21867 20284 22477 20312
rect 21867 20281 21879 20284
rect 21821 20275 21879 20281
rect 22465 20281 22477 20284
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 22922 20272 22928 20324
rect 22980 20312 22986 20324
rect 23290 20312 23296 20324
rect 22980 20284 23296 20312
rect 22980 20272 22986 20284
rect 23290 20272 23296 20284
rect 23348 20312 23354 20324
rect 23385 20315 23443 20321
rect 23385 20312 23397 20315
rect 23348 20284 23397 20312
rect 23348 20272 23354 20284
rect 23385 20281 23397 20284
rect 23431 20312 23443 20315
rect 23906 20315 23964 20321
rect 23906 20312 23918 20315
rect 23431 20284 23918 20312
rect 23431 20281 23443 20284
rect 23385 20275 23443 20281
rect 23906 20281 23918 20284
rect 23952 20281 23964 20315
rect 23906 20275 23964 20281
rect 8018 20204 8024 20256
rect 8076 20244 8082 20256
rect 8941 20247 8999 20253
rect 8941 20244 8953 20247
rect 8076 20216 8953 20244
rect 8076 20204 8082 20216
rect 8941 20213 8953 20216
rect 8987 20213 8999 20247
rect 9950 20244 9956 20256
rect 9911 20216 9956 20244
rect 8941 20207 8999 20213
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 10689 20247 10747 20253
rect 10689 20213 10701 20247
rect 10735 20244 10747 20247
rect 10778 20244 10784 20256
rect 10735 20216 10784 20244
rect 10735 20213 10747 20216
rect 10689 20207 10747 20213
rect 10778 20204 10784 20216
rect 10836 20244 10842 20256
rect 11238 20244 11244 20256
rect 10836 20216 11244 20244
rect 10836 20204 10842 20216
rect 11238 20204 11244 20216
rect 11296 20204 11302 20256
rect 13265 20247 13323 20253
rect 13265 20213 13277 20247
rect 13311 20244 13323 20247
rect 13354 20244 13360 20256
rect 13311 20216 13360 20244
rect 13311 20213 13323 20216
rect 13265 20207 13323 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 15930 20204 15936 20256
rect 15988 20244 15994 20256
rect 17773 20247 17831 20253
rect 17773 20244 17785 20247
rect 15988 20216 17785 20244
rect 15988 20204 15994 20216
rect 17773 20213 17785 20216
rect 17819 20213 17831 20247
rect 18782 20244 18788 20256
rect 18743 20216 18788 20244
rect 17773 20207 17831 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 19978 20204 19984 20256
rect 20036 20244 20042 20256
rect 20438 20244 20444 20256
rect 20036 20216 20444 20244
rect 20036 20204 20042 20216
rect 20438 20204 20444 20216
rect 20496 20244 20502 20256
rect 20901 20247 20959 20253
rect 20901 20244 20913 20247
rect 20496 20216 20913 20244
rect 20496 20204 20502 20216
rect 20901 20213 20913 20216
rect 20947 20213 20959 20247
rect 22002 20244 22008 20256
rect 21963 20216 22008 20244
rect 20901 20207 20959 20213
rect 22002 20204 22008 20216
rect 22060 20204 22066 20256
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 22373 20247 22431 20253
rect 22373 20244 22385 20247
rect 22152 20216 22385 20244
rect 22152 20204 22158 20216
rect 22373 20213 22385 20216
rect 22419 20213 22431 20247
rect 22373 20207 22431 20213
rect 24578 20204 24584 20256
rect 24636 20244 24642 20256
rect 25041 20247 25099 20253
rect 25041 20244 25053 20247
rect 24636 20216 25053 20244
rect 24636 20204 24642 20216
rect 25041 20213 25053 20216
rect 25087 20213 25099 20247
rect 25041 20207 25099 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 7834 20040 7840 20052
rect 7795 20012 7840 20040
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 11057 20043 11115 20049
rect 11057 20040 11069 20043
rect 10008 20012 11069 20040
rect 10008 20000 10014 20012
rect 11057 20009 11069 20012
rect 11103 20009 11115 20043
rect 11057 20003 11115 20009
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 12713 20043 12771 20049
rect 12713 20040 12725 20043
rect 12676 20012 12725 20040
rect 12676 20000 12682 20012
rect 12713 20009 12725 20012
rect 12759 20009 12771 20043
rect 13906 20040 13912 20052
rect 13867 20012 13912 20040
rect 12713 20003 12771 20009
rect 13906 20000 13912 20012
rect 13964 20040 13970 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 13964 20012 15025 20040
rect 13964 20000 13970 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 15749 20043 15807 20049
rect 15749 20009 15761 20043
rect 15795 20040 15807 20043
rect 16758 20040 16764 20052
rect 15795 20012 16764 20040
rect 15795 20009 15807 20012
rect 15749 20003 15807 20009
rect 16758 20000 16764 20012
rect 16816 20000 16822 20052
rect 17218 20040 17224 20052
rect 17179 20012 17224 20040
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 18325 20043 18383 20049
rect 18325 20009 18337 20043
rect 18371 20040 18383 20043
rect 19518 20040 19524 20052
rect 18371 20012 19524 20040
rect 18371 20009 18383 20012
rect 18325 20003 18383 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 20530 20000 20536 20052
rect 20588 20040 20594 20052
rect 20625 20043 20683 20049
rect 20625 20040 20637 20043
rect 20588 20012 20637 20040
rect 20588 20000 20594 20012
rect 20625 20009 20637 20012
rect 20671 20009 20683 20043
rect 20625 20003 20683 20009
rect 22002 20000 22008 20052
rect 22060 20040 22066 20052
rect 22833 20043 22891 20049
rect 22833 20040 22845 20043
rect 22060 20012 22845 20040
rect 22060 20000 22066 20012
rect 22833 20009 22845 20012
rect 22879 20009 22891 20043
rect 22833 20003 22891 20009
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 23937 20043 23995 20049
rect 23937 20040 23949 20043
rect 23348 20012 23949 20040
rect 23348 20000 23354 20012
rect 23937 20009 23949 20012
rect 23983 20009 23995 20043
rect 23937 20003 23995 20009
rect 24305 20043 24363 20049
rect 24305 20009 24317 20043
rect 24351 20040 24363 20043
rect 24762 20040 24768 20052
rect 24351 20012 24768 20040
rect 24351 20009 24363 20012
rect 24305 20003 24363 20009
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 18598 19932 18604 19984
rect 18656 19972 18662 19984
rect 18785 19975 18843 19981
rect 18785 19972 18797 19975
rect 18656 19944 18797 19972
rect 18656 19932 18662 19944
rect 18785 19941 18797 19944
rect 18831 19941 18843 19975
rect 21174 19972 21180 19984
rect 21135 19944 21180 19972
rect 18785 19935 18843 19941
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 22152 19944 22197 19972
rect 22152 19932 22158 19944
rect 7742 19904 7748 19916
rect 7703 19876 7748 19904
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 9674 19904 9680 19916
rect 9635 19876 9680 19904
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 9950 19913 9956 19916
rect 9944 19867 9956 19913
rect 10008 19904 10014 19916
rect 10008 19876 10044 19904
rect 9950 19864 9956 19867
rect 10008 19864 10014 19876
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 12158 19904 12164 19916
rect 11112 19876 12164 19904
rect 11112 19864 11118 19876
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 14093 19907 14151 19913
rect 14093 19873 14105 19907
rect 14139 19904 14151 19907
rect 14274 19904 14280 19916
rect 14139 19876 14280 19904
rect 14139 19873 14151 19876
rect 14093 19867 14151 19873
rect 14274 19864 14280 19876
rect 14332 19864 14338 19916
rect 15930 19864 15936 19916
rect 15988 19904 15994 19916
rect 16097 19907 16155 19913
rect 16097 19904 16109 19907
rect 15988 19876 16109 19904
rect 15988 19864 15994 19876
rect 16097 19873 16109 19876
rect 16143 19873 16155 19907
rect 16097 19867 16155 19873
rect 18046 19864 18052 19916
rect 18104 19904 18110 19916
rect 18509 19907 18567 19913
rect 18509 19904 18521 19907
rect 18104 19876 18521 19904
rect 18104 19864 18110 19876
rect 18509 19873 18521 19876
rect 18555 19904 18567 19907
rect 19150 19904 19156 19916
rect 18555 19876 19156 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 19610 19904 19616 19916
rect 19523 19876 19616 19904
rect 19610 19864 19616 19876
rect 19668 19904 19674 19916
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 19668 19876 20269 19904
rect 19668 19864 19674 19876
rect 20257 19873 20269 19876
rect 20303 19873 20315 19907
rect 20257 19867 20315 19873
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19873 20959 19907
rect 22738 19904 22744 19916
rect 22699 19876 22744 19904
rect 20901 19867 20959 19873
rect 8018 19836 8024 19848
rect 7979 19808 8024 19836
rect 8018 19796 8024 19808
rect 8076 19796 8082 19848
rect 12802 19836 12808 19848
rect 12763 19808 12808 19836
rect 12802 19796 12808 19808
rect 12860 19796 12866 19848
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19836 14795 19839
rect 15562 19836 15568 19848
rect 14783 19808 15568 19836
rect 14783 19805 14795 19808
rect 14737 19799 14795 19805
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 12912 19768 12940 19799
rect 15562 19796 15568 19808
rect 15620 19836 15626 19848
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 15620 19808 15853 19836
rect 15620 19796 15626 19808
rect 15841 19805 15853 19808
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 19518 19796 19524 19848
rect 19576 19836 19582 19848
rect 19705 19839 19763 19845
rect 19705 19836 19717 19839
rect 19576 19808 19717 19836
rect 19576 19796 19582 19808
rect 19705 19805 19717 19808
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 19978 19836 19984 19848
rect 19935 19808 19984 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 11940 19740 12940 19768
rect 19245 19771 19303 19777
rect 11940 19728 11946 19740
rect 19245 19737 19257 19771
rect 19291 19768 19303 19771
rect 20916 19768 20944 19867
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 24394 19904 24400 19916
rect 24355 19876 24400 19904
rect 24394 19864 24400 19876
rect 24452 19864 24458 19916
rect 22922 19836 22928 19848
rect 22883 19808 22928 19836
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 24578 19836 24584 19848
rect 24539 19808 24584 19836
rect 24578 19796 24584 19808
rect 24636 19836 24642 19848
rect 24854 19836 24860 19848
rect 24636 19808 24860 19836
rect 24636 19796 24642 19808
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 21637 19771 21695 19777
rect 21637 19768 21649 19771
rect 19291 19740 21649 19768
rect 19291 19737 19303 19740
rect 19245 19731 19303 19737
rect 21637 19737 21649 19740
rect 21683 19737 21695 19771
rect 21637 19731 21695 19737
rect 22373 19771 22431 19777
rect 22373 19737 22385 19771
rect 22419 19768 22431 19771
rect 24118 19768 24124 19780
rect 22419 19740 24124 19768
rect 22419 19737 22431 19740
rect 22373 19731 22431 19737
rect 24118 19728 24124 19740
rect 24176 19768 24182 19780
rect 24949 19771 25007 19777
rect 24949 19768 24961 19771
rect 24176 19740 24961 19768
rect 24176 19728 24182 19740
rect 24949 19737 24961 19740
rect 24995 19737 25007 19771
rect 24949 19731 25007 19737
rect 7377 19703 7435 19709
rect 7377 19669 7389 19703
rect 7423 19700 7435 19703
rect 8202 19700 8208 19712
rect 7423 19672 8208 19700
rect 7423 19669 7435 19672
rect 7377 19663 7435 19669
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 12250 19660 12256 19712
rect 12308 19700 12314 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 12308 19672 12357 19700
rect 12308 19660 12314 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 13354 19700 13360 19712
rect 13315 19672 13360 19700
rect 12345 19663 12403 19669
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13814 19700 13820 19712
rect 13775 19672 13820 19700
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 18141 19703 18199 19709
rect 18141 19669 18153 19703
rect 18187 19700 18199 19703
rect 18414 19700 18420 19712
rect 18187 19672 18420 19700
rect 18187 19669 18199 19672
rect 18141 19663 18199 19669
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 23658 19700 23664 19712
rect 23619 19672 23664 19700
rect 23658 19660 23664 19672
rect 23716 19660 23722 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 7469 19499 7527 19505
rect 7469 19465 7481 19499
rect 7515 19496 7527 19499
rect 7834 19496 7840 19508
rect 7515 19468 7840 19496
rect 7515 19465 7527 19468
rect 7469 19459 7527 19465
rect 7834 19456 7840 19468
rect 7892 19456 7898 19508
rect 9950 19496 9956 19508
rect 9911 19468 9956 19496
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 11882 19496 11888 19508
rect 11843 19468 11888 19496
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 16390 19496 16396 19508
rect 16351 19468 16396 19496
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 19610 19456 19616 19508
rect 19668 19496 19674 19508
rect 19705 19499 19763 19505
rect 19705 19496 19717 19499
rect 19668 19468 19717 19496
rect 19668 19456 19674 19468
rect 19705 19465 19717 19468
rect 19751 19465 19763 19499
rect 19705 19459 19763 19465
rect 22465 19499 22523 19505
rect 22465 19465 22477 19499
rect 22511 19496 22523 19499
rect 22922 19496 22928 19508
rect 22511 19468 22928 19496
rect 22511 19465 22523 19468
rect 22465 19459 22523 19465
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 23658 19456 23664 19508
rect 23716 19496 23722 19508
rect 23716 19468 23796 19496
rect 23716 19456 23722 19468
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19360 7159 19363
rect 11425 19363 11483 19369
rect 7147 19332 8156 19360
rect 7147 19329 7159 19332
rect 7101 19323 7159 19329
rect 8128 19304 8156 19332
rect 11425 19329 11437 19363
rect 11471 19360 11483 19363
rect 11900 19360 11928 19456
rect 22186 19428 22192 19440
rect 19260 19400 22192 19428
rect 12618 19360 12624 19372
rect 11471 19332 11928 19360
rect 12360 19332 12624 19360
rect 11471 19329 11483 19332
rect 11425 19323 11483 19329
rect 7558 19252 7564 19304
rect 7616 19292 7622 19304
rect 8021 19295 8079 19301
rect 8021 19292 8033 19295
rect 7616 19264 8033 19292
rect 7616 19252 7622 19264
rect 8021 19261 8033 19264
rect 8067 19261 8079 19295
rect 8021 19255 8079 19261
rect 7834 19224 7840 19236
rect 7795 19196 7840 19224
rect 7834 19184 7840 19196
rect 7892 19184 7898 19236
rect 8036 19224 8064 19255
rect 8110 19252 8116 19304
rect 8168 19292 8174 19304
rect 8277 19295 8335 19301
rect 8277 19292 8289 19295
rect 8168 19264 8289 19292
rect 8168 19252 8174 19264
rect 8277 19261 8289 19264
rect 8323 19261 8335 19295
rect 8277 19255 8335 19261
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12360 19292 12388 19332
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 16022 19320 16028 19372
rect 16080 19360 16086 19372
rect 16945 19363 17003 19369
rect 16945 19360 16957 19363
rect 16080 19332 16957 19360
rect 16080 19320 16086 19332
rect 16945 19329 16957 19332
rect 16991 19360 17003 19363
rect 17405 19363 17463 19369
rect 17405 19360 17417 19363
rect 16991 19332 17417 19360
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17405 19329 17417 19332
rect 17451 19360 17463 19363
rect 18598 19360 18604 19372
rect 17451 19332 18604 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 19260 19304 19288 19400
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 23768 19428 23796 19468
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24673 19499 24731 19505
rect 24673 19496 24685 19499
rect 24084 19468 24685 19496
rect 24084 19456 24090 19468
rect 24673 19465 24685 19468
rect 24719 19465 24731 19499
rect 24673 19459 24731 19465
rect 23768 19400 24072 19428
rect 24044 19372 24072 19400
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 20128 19332 20269 19360
rect 20128 19320 20134 19332
rect 20257 19329 20269 19332
rect 20303 19329 20315 19363
rect 21818 19360 21824 19372
rect 21779 19332 21824 19360
rect 20257 19323 20315 19329
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 24026 19320 24032 19372
rect 24084 19320 24090 19372
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19360 24363 19363
rect 24486 19360 24492 19372
rect 24351 19332 24492 19360
rect 24351 19329 24363 19332
rect 24305 19323 24363 19329
rect 12299 19264 12388 19292
rect 12805 19295 12863 19301
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12805 19261 12817 19295
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 13072 19295 13130 19301
rect 13072 19261 13084 19295
rect 13118 19292 13130 19295
rect 13354 19292 13360 19304
rect 13118 19264 13360 19292
rect 13118 19261 13130 19264
rect 13072 19255 13130 19261
rect 8386 19224 8392 19236
rect 8036 19196 8392 19224
rect 8386 19184 8392 19196
rect 8444 19184 8450 19236
rect 10594 19224 10600 19236
rect 10555 19196 10600 19224
rect 10594 19184 10600 19196
rect 10652 19224 10658 19236
rect 11241 19227 11299 19233
rect 11241 19224 11253 19227
rect 10652 19196 11253 19224
rect 10652 19184 10658 19196
rect 11241 19193 11253 19196
rect 11287 19193 11299 19227
rect 12820 19224 12848 19255
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 15933 19295 15991 19301
rect 15933 19261 15945 19295
rect 15979 19292 15991 19295
rect 16761 19295 16819 19301
rect 16761 19292 16773 19295
rect 15979 19264 16773 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 16761 19261 16773 19264
rect 16807 19292 16819 19295
rect 16850 19292 16856 19304
rect 16807 19264 16856 19292
rect 16807 19261 16819 19264
rect 16761 19255 16819 19261
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 18138 19292 18144 19304
rect 17911 19264 18144 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 18414 19292 18420 19304
rect 18375 19264 18420 19292
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 19242 19252 19248 19304
rect 19300 19252 19306 19304
rect 21174 19292 21180 19304
rect 21135 19264 21180 19292
rect 21174 19252 21180 19264
rect 21232 19292 21238 19304
rect 21729 19295 21787 19301
rect 21729 19292 21741 19295
rect 21232 19264 21741 19292
rect 21232 19252 21238 19264
rect 21729 19261 21741 19264
rect 21775 19261 21787 19295
rect 23106 19292 23112 19304
rect 23019 19264 23112 19292
rect 21729 19255 21787 19261
rect 23106 19252 23112 19264
rect 23164 19292 23170 19304
rect 24320 19292 24348 19323
rect 24486 19320 24492 19332
rect 24544 19360 24550 19372
rect 24854 19360 24860 19372
rect 24544 19332 24860 19360
rect 24544 19320 24550 19332
rect 24854 19320 24860 19332
rect 24912 19320 24918 19372
rect 25038 19292 25044 19304
rect 23164 19264 24348 19292
rect 24999 19264 25044 19292
rect 23164 19252 23170 19264
rect 25038 19252 25044 19264
rect 25096 19252 25102 19304
rect 25222 19292 25228 19304
rect 25183 19264 25228 19292
rect 25222 19252 25228 19264
rect 25280 19292 25286 19304
rect 25961 19295 26019 19301
rect 25961 19292 25973 19295
rect 25280 19264 25973 19292
rect 25280 19252 25286 19264
rect 25961 19261 25973 19264
rect 26007 19261 26019 19295
rect 25961 19255 26019 19261
rect 13814 19224 13820 19236
rect 12820 19196 13820 19224
rect 11241 19187 11299 19193
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 15381 19227 15439 19233
rect 15381 19193 15393 19227
rect 15427 19224 15439 19227
rect 19153 19227 19211 19233
rect 19153 19224 19165 19227
rect 15427 19196 19165 19224
rect 15427 19193 15439 19196
rect 15381 19187 15439 19193
rect 19153 19193 19165 19196
rect 19199 19224 19211 19227
rect 20073 19227 20131 19233
rect 20073 19224 20085 19227
rect 19199 19196 20085 19224
rect 19199 19193 19211 19196
rect 19153 19187 19211 19193
rect 20073 19193 20085 19196
rect 20119 19193 20131 19227
rect 20073 19187 20131 19193
rect 20809 19227 20867 19233
rect 20809 19193 20821 19227
rect 20855 19224 20867 19227
rect 21637 19227 21695 19233
rect 21637 19224 21649 19227
rect 20855 19196 21649 19224
rect 20855 19193 20867 19196
rect 20809 19187 20867 19193
rect 21637 19193 21649 19196
rect 21683 19224 21695 19227
rect 21910 19224 21916 19236
rect 21683 19196 21916 19224
rect 21683 19193 21695 19196
rect 21637 19187 21695 19193
rect 21910 19184 21916 19196
rect 21968 19184 21974 19236
rect 23474 19224 23480 19236
rect 23387 19196 23480 19224
rect 23474 19184 23480 19196
rect 23532 19224 23538 19236
rect 25498 19224 25504 19236
rect 23532 19196 24164 19224
rect 25459 19196 25504 19224
rect 23532 19184 23538 19196
rect 9398 19156 9404 19168
rect 9359 19128 9404 19156
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 10781 19159 10839 19165
rect 10781 19125 10793 19159
rect 10827 19156 10839 19159
rect 10870 19156 10876 19168
rect 10827 19128 10876 19156
rect 10827 19125 10839 19128
rect 10781 19119 10839 19125
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 11146 19156 11152 19168
rect 11107 19128 11152 19156
rect 11146 19116 11152 19128
rect 11204 19156 11210 19168
rect 12066 19156 12072 19168
rect 11204 19128 12072 19156
rect 11204 19116 11210 19128
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12713 19159 12771 19165
rect 12713 19125 12725 19159
rect 12759 19156 12771 19159
rect 12802 19156 12808 19168
rect 12759 19128 12808 19156
rect 12759 19125 12771 19128
rect 12713 19119 12771 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 14182 19156 14188 19168
rect 14143 19128 14188 19156
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14332 19128 14749 19156
rect 14332 19116 14338 19128
rect 14737 19125 14749 19128
rect 14783 19125 14795 19159
rect 14737 19119 14795 19125
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15562 19156 15568 19168
rect 15335 19128 15568 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16301 19159 16359 19165
rect 16301 19125 16313 19159
rect 16347 19156 16359 19159
rect 16853 19159 16911 19165
rect 16853 19156 16865 19159
rect 16347 19128 16865 19156
rect 16347 19125 16359 19128
rect 16301 19119 16359 19125
rect 16853 19125 16865 19128
rect 16899 19156 16911 19159
rect 17126 19156 17132 19168
rect 16899 19128 17132 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 17126 19116 17132 19128
rect 17184 19116 17190 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18049 19159 18107 19165
rect 18049 19156 18061 19159
rect 18012 19128 18061 19156
rect 18012 19116 18018 19128
rect 18049 19125 18061 19128
rect 18095 19125 18107 19159
rect 18049 19119 18107 19125
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18509 19159 18567 19165
rect 18509 19156 18521 19159
rect 18196 19128 18521 19156
rect 18196 19116 18202 19128
rect 18509 19125 18521 19128
rect 18555 19156 18567 19159
rect 19242 19156 19248 19168
rect 18555 19128 19248 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 19334 19116 19340 19168
rect 19392 19156 19398 19168
rect 19521 19159 19579 19165
rect 19521 19156 19533 19159
rect 19392 19128 19533 19156
rect 19392 19116 19398 19128
rect 19521 19125 19533 19128
rect 19567 19156 19579 19159
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 19567 19128 20177 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 20165 19125 20177 19128
rect 20211 19156 20223 19159
rect 20714 19156 20720 19168
rect 20211 19128 20720 19156
rect 20211 19125 20223 19128
rect 20165 19119 20223 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 23661 19159 23719 19165
rect 23661 19156 23673 19159
rect 22520 19128 23673 19156
rect 22520 19116 22526 19128
rect 23661 19125 23673 19128
rect 23707 19125 23719 19159
rect 24026 19156 24032 19168
rect 23987 19128 24032 19156
rect 23661 19119 23719 19125
rect 24026 19116 24032 19128
rect 24084 19116 24090 19168
rect 24136 19165 24164 19196
rect 25498 19184 25504 19196
rect 25556 19184 25562 19236
rect 24121 19159 24179 19165
rect 24121 19125 24133 19159
rect 24167 19156 24179 19159
rect 24210 19156 24216 19168
rect 24167 19128 24216 19156
rect 24167 19125 24179 19128
rect 24121 19119 24179 19125
rect 24210 19116 24216 19128
rect 24268 19116 24274 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 8018 18952 8024 18964
rect 7979 18924 8024 18952
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 8386 18952 8392 18964
rect 8347 18924 8392 18952
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9306 18952 9312 18964
rect 9219 18924 9312 18952
rect 9306 18912 9312 18924
rect 9364 18952 9370 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 9364 18924 11621 18952
rect 9364 18912 9370 18924
rect 11609 18921 11621 18924
rect 11655 18952 11667 18955
rect 11790 18952 11796 18964
rect 11655 18924 11796 18952
rect 11655 18921 11667 18924
rect 11609 18915 11667 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 13173 18955 13231 18961
rect 13173 18921 13185 18955
rect 13219 18952 13231 18955
rect 13354 18952 13360 18964
rect 13219 18924 13360 18952
rect 13219 18921 13231 18924
rect 13173 18915 13231 18921
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 15930 18952 15936 18964
rect 15891 18924 15936 18952
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 19518 18912 19524 18964
rect 19576 18952 19582 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19576 18924 19717 18952
rect 19576 18912 19582 18924
rect 19705 18921 19717 18924
rect 19751 18952 19763 18955
rect 21266 18952 21272 18964
rect 19751 18924 21272 18952
rect 19751 18921 19763 18924
rect 19705 18915 19763 18921
rect 21266 18912 21272 18924
rect 21324 18912 21330 18964
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 24213 18955 24271 18961
rect 22152 18924 22197 18952
rect 22152 18912 22158 18924
rect 24213 18921 24225 18955
rect 24259 18952 24271 18955
rect 24762 18952 24768 18964
rect 24259 18924 24768 18952
rect 24259 18921 24271 18924
rect 24213 18915 24271 18921
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 10134 18844 10140 18896
rect 10192 18884 10198 18896
rect 10781 18887 10839 18893
rect 10781 18884 10793 18887
rect 10192 18856 10793 18884
rect 10192 18844 10198 18856
rect 10781 18853 10793 18856
rect 10827 18884 10839 18887
rect 11146 18884 11152 18896
rect 10827 18856 11152 18884
rect 10827 18853 10839 18856
rect 10781 18847 10839 18853
rect 11146 18844 11152 18856
rect 11204 18844 11210 18896
rect 11241 18887 11299 18893
rect 11241 18853 11253 18887
rect 11287 18884 11299 18887
rect 11882 18884 11888 18896
rect 11287 18856 11888 18884
rect 11287 18853 11299 18856
rect 11241 18847 11299 18853
rect 11882 18844 11888 18856
rect 11940 18884 11946 18896
rect 12038 18887 12096 18893
rect 12038 18884 12050 18887
rect 11940 18856 12050 18884
rect 11940 18844 11946 18856
rect 12038 18853 12050 18856
rect 12084 18884 12096 18887
rect 12342 18884 12348 18896
rect 12084 18856 12348 18884
rect 12084 18853 12096 18856
rect 12038 18847 12096 18853
rect 12342 18844 12348 18856
rect 12400 18844 12406 18896
rect 17954 18844 17960 18896
rect 18012 18884 18018 18896
rect 18509 18887 18567 18893
rect 18509 18884 18521 18887
rect 18012 18856 18521 18884
rect 18012 18844 18018 18856
rect 18509 18853 18521 18856
rect 18555 18853 18567 18887
rect 18509 18847 18567 18853
rect 19337 18887 19395 18893
rect 19337 18853 19349 18887
rect 19383 18884 19395 18887
rect 19978 18884 19984 18896
rect 19383 18856 19984 18884
rect 19383 18853 19395 18856
rect 19337 18847 19395 18853
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 20070 18844 20076 18896
rect 20128 18884 20134 18896
rect 20257 18887 20315 18893
rect 20257 18884 20269 18887
rect 20128 18856 20269 18884
rect 20128 18844 20134 18856
rect 20257 18853 20269 18856
rect 20303 18884 20315 18887
rect 21637 18887 21695 18893
rect 21637 18884 21649 18887
rect 20303 18856 21649 18884
rect 20303 18853 20315 18856
rect 20257 18847 20315 18853
rect 21637 18853 21649 18856
rect 21683 18884 21695 18887
rect 21818 18884 21824 18896
rect 21683 18856 21824 18884
rect 21683 18853 21695 18856
rect 21637 18847 21695 18853
rect 21818 18844 21824 18856
rect 21876 18844 21882 18896
rect 22456 18887 22514 18893
rect 22456 18853 22468 18887
rect 22502 18884 22514 18887
rect 23106 18884 23112 18896
rect 22502 18856 23112 18884
rect 22502 18853 22514 18856
rect 22456 18847 22514 18853
rect 23106 18844 23112 18856
rect 23164 18844 23170 18896
rect 24486 18884 24492 18896
rect 24447 18856 24492 18884
rect 24486 18844 24492 18856
rect 24544 18844 24550 18896
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 8754 18816 8760 18828
rect 8444 18788 8760 18816
rect 8444 18776 8450 18788
rect 8754 18776 8760 18788
rect 8812 18816 8818 18828
rect 9309 18819 9367 18825
rect 9309 18816 9321 18819
rect 8812 18788 9321 18816
rect 8812 18776 8818 18788
rect 9309 18785 9321 18788
rect 9355 18816 9367 18819
rect 9401 18819 9459 18825
rect 9401 18816 9413 18819
rect 9355 18788 9413 18816
rect 9355 18785 9367 18788
rect 9309 18779 9367 18785
rect 9401 18785 9413 18788
rect 9447 18785 9459 18819
rect 10042 18816 10048 18828
rect 9955 18788 10048 18816
rect 9401 18779 9459 18785
rect 10042 18776 10048 18788
rect 10100 18816 10106 18828
rect 11422 18816 11428 18828
rect 10100 18788 11428 18816
rect 10100 18776 10106 18788
rect 11422 18776 11428 18788
rect 11480 18776 11486 18828
rect 11790 18816 11796 18828
rect 11751 18788 11796 18816
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 14185 18819 14243 18825
rect 14185 18785 14197 18819
rect 14231 18816 14243 18819
rect 14461 18819 14519 18825
rect 14461 18816 14473 18819
rect 14231 18788 14473 18816
rect 14231 18785 14243 18788
rect 14185 18779 14243 18785
rect 14461 18785 14473 18788
rect 14507 18816 14519 18819
rect 14826 18816 14832 18828
rect 14507 18788 14832 18816
rect 14507 18785 14519 18788
rect 14461 18779 14519 18785
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 16853 18819 16911 18825
rect 16853 18816 16865 18819
rect 16080 18788 16865 18816
rect 16080 18776 16086 18788
rect 16853 18785 16865 18788
rect 16899 18816 16911 18819
rect 17402 18816 17408 18828
rect 16899 18788 17408 18816
rect 16899 18785 16911 18788
rect 16853 18779 16911 18785
rect 17402 18776 17408 18788
rect 17460 18776 17466 18828
rect 17589 18819 17647 18825
rect 17589 18785 17601 18819
rect 17635 18816 17647 18819
rect 18414 18816 18420 18828
rect 17635 18788 18420 18816
rect 17635 18785 17647 18788
rect 17589 18779 17647 18785
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 21082 18816 21088 18828
rect 21043 18788 21088 18816
rect 21082 18776 21088 18788
rect 21140 18776 21146 18828
rect 21358 18776 21364 18828
rect 21416 18816 21422 18828
rect 25038 18816 25044 18828
rect 21416 18788 25044 18816
rect 21416 18776 21422 18788
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 25130 18776 25136 18828
rect 25188 18816 25194 18828
rect 25406 18816 25412 18828
rect 25188 18788 25412 18816
rect 25188 18776 25194 18788
rect 25406 18776 25412 18788
rect 25464 18776 25470 18828
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10134 18748 10140 18760
rect 9732 18720 10140 18748
rect 9732 18708 9738 18720
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18717 10287 18751
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 10229 18711 10287 18717
rect 9950 18640 9956 18692
rect 10008 18680 10014 18692
rect 10244 18680 10272 18711
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16632 18720 16957 18748
rect 16632 18708 16638 18720
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 17494 18748 17500 18760
rect 17175 18720 17500 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 10008 18652 10272 18680
rect 16960 18680 16988 18711
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 18598 18708 18604 18760
rect 18656 18748 18662 18760
rect 19797 18751 19855 18757
rect 18656 18720 18701 18748
rect 18656 18708 18662 18720
rect 19797 18717 19809 18751
rect 19843 18748 19855 18751
rect 20622 18748 20628 18760
rect 19843 18720 20628 18748
rect 19843 18717 19855 18720
rect 19797 18711 19855 18717
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18748 20775 18751
rect 22094 18748 22100 18760
rect 20763 18720 22100 18748
rect 20763 18717 20775 18720
rect 20717 18711 20775 18717
rect 22094 18708 22100 18720
rect 22152 18748 22158 18760
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 22152 18720 22201 18748
rect 22152 18708 22158 18720
rect 22189 18717 22201 18720
rect 22235 18717 22247 18751
rect 25222 18748 25228 18760
rect 25183 18720 25228 18748
rect 22189 18711 22247 18717
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 17402 18680 17408 18692
rect 16960 18652 17408 18680
rect 10008 18640 10014 18652
rect 17402 18640 17408 18652
rect 17460 18640 17466 18692
rect 17957 18683 18015 18689
rect 17957 18649 17969 18683
rect 18003 18680 18015 18683
rect 18616 18680 18644 18708
rect 18003 18652 18644 18680
rect 18003 18649 18015 18652
rect 17957 18643 18015 18649
rect 9674 18612 9680 18624
rect 9635 18584 9680 18612
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 13722 18612 13728 18624
rect 13683 18584 13728 18612
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 14274 18612 14280 18624
rect 14235 18584 14280 18612
rect 14274 18572 14280 18584
rect 14332 18572 14338 18624
rect 15013 18615 15071 18621
rect 15013 18581 15025 18615
rect 15059 18612 15071 18615
rect 15470 18612 15476 18624
rect 15059 18584 15476 18612
rect 15059 18581 15071 18584
rect 15013 18575 15071 18581
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 16206 18612 16212 18624
rect 16167 18584 16212 18612
rect 16206 18572 16212 18584
rect 16264 18572 16270 18624
rect 16482 18612 16488 18624
rect 16443 18584 16488 18612
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 18046 18612 18052 18624
rect 18007 18584 18052 18612
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 21266 18612 21272 18624
rect 21227 18584 21272 18612
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 23569 18615 23627 18621
rect 23569 18612 23581 18615
rect 23532 18584 23581 18612
rect 23532 18572 23538 18584
rect 23569 18581 23581 18584
rect 23615 18581 23627 18615
rect 24670 18612 24676 18624
rect 24631 18584 24676 18612
rect 23569 18575 23627 18581
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 10137 18411 10195 18417
rect 10137 18408 10149 18411
rect 10008 18380 10149 18408
rect 10008 18368 10014 18380
rect 10137 18377 10149 18380
rect 10183 18408 10195 18411
rect 10689 18411 10747 18417
rect 10689 18408 10701 18411
rect 10183 18380 10701 18408
rect 10183 18377 10195 18380
rect 10137 18371 10195 18377
rect 10689 18377 10701 18380
rect 10735 18377 10747 18411
rect 11422 18408 11428 18420
rect 11383 18380 11428 18408
rect 10689 18371 10747 18377
rect 11422 18368 11428 18380
rect 11480 18368 11486 18420
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 13906 18408 13912 18420
rect 12400 18380 13912 18408
rect 12400 18368 12406 18380
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 14090 18368 14096 18420
rect 14148 18408 14154 18420
rect 14737 18411 14795 18417
rect 14737 18408 14749 18411
rect 14148 18380 14749 18408
rect 14148 18368 14154 18380
rect 14737 18377 14749 18380
rect 14783 18408 14795 18411
rect 14826 18408 14832 18420
rect 14783 18380 14832 18408
rect 14783 18377 14795 18380
rect 14737 18371 14795 18377
rect 14826 18368 14832 18380
rect 14884 18368 14890 18420
rect 20346 18368 20352 18420
rect 20404 18408 20410 18420
rect 20530 18408 20536 18420
rect 20404 18380 20536 18408
rect 20404 18368 20410 18380
rect 20530 18368 20536 18380
rect 20588 18368 20594 18420
rect 21082 18408 21088 18420
rect 21043 18380 21088 18408
rect 21082 18368 21088 18380
rect 21140 18368 21146 18420
rect 22002 18408 22008 18420
rect 21963 18380 22008 18408
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 23106 18408 23112 18420
rect 23067 18380 23112 18408
rect 23106 18368 23112 18380
rect 23164 18368 23170 18420
rect 25041 18411 25099 18417
rect 25041 18377 25053 18411
rect 25087 18408 25099 18411
rect 25222 18408 25228 18420
rect 25087 18380 25228 18408
rect 25087 18377 25099 18380
rect 25041 18371 25099 18377
rect 25222 18368 25228 18380
rect 25280 18368 25286 18420
rect 14921 18343 14979 18349
rect 14921 18309 14933 18343
rect 14967 18340 14979 18343
rect 15378 18340 15384 18352
rect 14967 18312 15384 18340
rect 14967 18309 14979 18312
rect 14921 18303 14979 18309
rect 15378 18300 15384 18312
rect 15436 18300 15442 18352
rect 20809 18343 20867 18349
rect 20809 18309 20821 18343
rect 20855 18340 20867 18343
rect 20990 18340 20996 18352
rect 20855 18312 20996 18340
rect 20855 18309 20867 18312
rect 20809 18303 20867 18309
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 8754 18272 8760 18284
rect 8715 18244 8760 18272
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 11057 18275 11115 18281
rect 11057 18272 11069 18275
rect 10192 18244 11069 18272
rect 10192 18232 10198 18244
rect 11057 18241 11069 18244
rect 11103 18241 11115 18275
rect 11057 18235 11115 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13817 18275 13875 18281
rect 13817 18272 13829 18275
rect 13219 18244 13829 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13817 18241 13829 18244
rect 13863 18272 13875 18275
rect 14182 18272 14188 18284
rect 13863 18244 14188 18272
rect 13863 18241 13875 18244
rect 13817 18235 13875 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 15470 18272 15476 18284
rect 15431 18244 15476 18272
rect 15470 18232 15476 18244
rect 15528 18232 15534 18284
rect 15562 18232 15568 18284
rect 15620 18272 15626 18284
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 15620 18244 18337 18272
rect 15620 18232 15626 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 20346 18272 20352 18284
rect 20307 18244 20352 18272
rect 18325 18235 18383 18241
rect 20346 18232 20352 18244
rect 20404 18272 20410 18284
rect 21913 18275 21971 18281
rect 20404 18244 20944 18272
rect 20404 18232 20410 18244
rect 9024 18207 9082 18213
rect 9024 18204 9036 18207
rect 8956 18176 9036 18204
rect 8665 18139 8723 18145
rect 8665 18105 8677 18139
rect 8711 18136 8723 18139
rect 8956 18136 8984 18176
rect 9024 18173 9036 18176
rect 9070 18204 9082 18207
rect 9398 18204 9404 18216
rect 9070 18176 9404 18204
rect 9070 18173 9082 18176
rect 9024 18167 9082 18173
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 13633 18207 13691 18213
rect 13633 18173 13645 18207
rect 13679 18204 13691 18207
rect 13722 18204 13728 18216
rect 13679 18176 13728 18204
rect 13679 18173 13691 18176
rect 13633 18167 13691 18173
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 16390 18164 16396 18216
rect 16448 18204 16454 18216
rect 16485 18207 16543 18213
rect 16485 18204 16497 18207
rect 16448 18176 16497 18204
rect 16448 18164 16454 18176
rect 16485 18173 16497 18176
rect 16531 18204 16543 18207
rect 16574 18204 16580 18216
rect 16531 18176 16580 18204
rect 16531 18173 16543 18176
rect 16485 18167 16543 18173
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 20916 18213 20944 18244
rect 21913 18241 21925 18275
rect 21959 18272 21971 18275
rect 22557 18275 22615 18281
rect 22557 18272 22569 18275
rect 21959 18244 22569 18272
rect 21959 18241 21971 18244
rect 21913 18235 21971 18241
rect 22557 18241 22569 18244
rect 22603 18272 22615 18275
rect 23385 18275 23443 18281
rect 23385 18272 23397 18275
rect 22603 18244 23397 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 23385 18241 23397 18244
rect 23431 18272 23443 18275
rect 23474 18272 23480 18284
rect 23431 18244 23480 18272
rect 23431 18241 23443 18244
rect 23385 18235 23443 18241
rect 23474 18232 23480 18244
rect 23532 18272 23538 18284
rect 23532 18244 23796 18272
rect 23532 18232 23538 18244
rect 20901 18207 20959 18213
rect 20901 18173 20913 18207
rect 20947 18173 20959 18207
rect 20901 18167 20959 18173
rect 21545 18207 21603 18213
rect 21545 18173 21557 18207
rect 21591 18204 21603 18207
rect 22462 18204 22468 18216
rect 21591 18176 22468 18204
rect 21591 18173 21603 18176
rect 21545 18167 21603 18173
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 23290 18164 23296 18216
rect 23348 18204 23354 18216
rect 23661 18207 23719 18213
rect 23661 18204 23673 18207
rect 23348 18176 23673 18204
rect 23348 18164 23354 18176
rect 23661 18173 23673 18176
rect 23707 18173 23719 18207
rect 23768 18204 23796 18244
rect 23917 18207 23975 18213
rect 23917 18204 23929 18207
rect 23768 18176 23929 18204
rect 23661 18167 23719 18173
rect 23917 18173 23929 18176
rect 23963 18173 23975 18207
rect 23917 18167 23975 18173
rect 8711 18108 8984 18136
rect 8711 18105 8723 18108
rect 8665 18099 8723 18105
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 12805 18139 12863 18145
rect 12805 18136 12817 18139
rect 12400 18108 12817 18136
rect 12400 18096 12406 18108
rect 12805 18105 12817 18108
rect 12851 18136 12863 18139
rect 12851 18108 13768 18136
rect 12851 18105 12863 18108
rect 12805 18099 12863 18105
rect 13265 18071 13323 18077
rect 13265 18037 13277 18071
rect 13311 18068 13323 18071
rect 13630 18068 13636 18080
rect 13311 18040 13636 18068
rect 13311 18037 13323 18040
rect 13265 18031 13323 18037
rect 13630 18028 13636 18040
rect 13688 18028 13694 18080
rect 13740 18077 13768 18108
rect 14826 18096 14832 18148
rect 14884 18136 14890 18148
rect 15381 18139 15439 18145
rect 15381 18136 15393 18139
rect 14884 18108 15393 18136
rect 14884 18096 14890 18108
rect 15381 18105 15393 18108
rect 15427 18105 15439 18139
rect 15381 18099 15439 18105
rect 16761 18139 16819 18145
rect 16761 18105 16773 18139
rect 16807 18136 16819 18139
rect 17678 18136 17684 18148
rect 16807 18108 17684 18136
rect 16807 18105 16819 18108
rect 16761 18099 16819 18105
rect 17678 18096 17684 18108
rect 17736 18096 17742 18148
rect 18598 18145 18604 18148
rect 17865 18139 17923 18145
rect 17865 18105 17877 18139
rect 17911 18136 17923 18139
rect 18592 18136 18604 18145
rect 17911 18108 18604 18136
rect 17911 18105 17923 18108
rect 17865 18099 17923 18105
rect 18592 18099 18604 18108
rect 18656 18136 18662 18148
rect 19150 18136 19156 18148
rect 18656 18108 19156 18136
rect 18598 18096 18604 18099
rect 18656 18096 18662 18108
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 22373 18139 22431 18145
rect 22373 18105 22385 18139
rect 22419 18136 22431 18139
rect 23198 18136 23204 18148
rect 22419 18108 23204 18136
rect 22419 18105 22431 18108
rect 22373 18099 22431 18105
rect 23198 18096 23204 18108
rect 23256 18096 23262 18148
rect 13725 18071 13783 18077
rect 13725 18037 13737 18071
rect 13771 18037 13783 18071
rect 14274 18068 14280 18080
rect 14235 18040 14280 18068
rect 13725 18031 13783 18037
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 14918 18068 14924 18080
rect 14792 18040 14924 18068
rect 14792 18028 14798 18040
rect 14918 18028 14924 18040
rect 14976 18068 14982 18080
rect 15289 18071 15347 18077
rect 15289 18068 15301 18071
rect 14976 18040 15301 18068
rect 14976 18028 14982 18040
rect 15289 18037 15301 18040
rect 15335 18037 15347 18071
rect 15289 18031 15347 18037
rect 15562 18028 15568 18080
rect 15620 18068 15626 18080
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 15620 18040 15945 18068
rect 15620 18028 15626 18040
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 16022 18028 16028 18080
rect 16080 18068 16086 18080
rect 16301 18071 16359 18077
rect 16301 18068 16313 18071
rect 16080 18040 16313 18068
rect 16080 18028 16086 18040
rect 16301 18037 16313 18040
rect 16347 18037 16359 18071
rect 16301 18031 16359 18037
rect 17313 18071 17371 18077
rect 17313 18037 17325 18071
rect 17359 18068 17371 18071
rect 17402 18068 17408 18080
rect 17359 18040 17408 18068
rect 17359 18037 17371 18040
rect 17313 18031 17371 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 19705 18071 19763 18077
rect 19705 18037 19717 18071
rect 19751 18068 19763 18071
rect 19978 18068 19984 18080
rect 19751 18040 19984 18068
rect 19751 18037 19763 18040
rect 19705 18031 19763 18037
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 23106 18028 23112 18080
rect 23164 18068 23170 18080
rect 24026 18068 24032 18080
rect 23164 18040 24032 18068
rect 23164 18028 23170 18040
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 25130 18028 25136 18080
rect 25188 18068 25194 18080
rect 25593 18071 25651 18077
rect 25593 18068 25605 18071
rect 25188 18040 25605 18068
rect 25188 18028 25194 18040
rect 25593 18037 25605 18040
rect 25639 18037 25651 18071
rect 25593 18031 25651 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 9125 17867 9183 17873
rect 9125 17864 9137 17867
rect 8352 17836 9137 17864
rect 8352 17824 8358 17836
rect 9125 17833 9137 17836
rect 9171 17864 9183 17867
rect 9582 17864 9588 17876
rect 9171 17836 9588 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10686 17864 10692 17876
rect 9732 17836 10692 17864
rect 9732 17824 9738 17836
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 10870 17824 10876 17876
rect 10928 17864 10934 17876
rect 11793 17867 11851 17873
rect 11793 17864 11805 17867
rect 10928 17836 11805 17864
rect 10928 17824 10934 17836
rect 11793 17833 11805 17836
rect 11839 17864 11851 17867
rect 11885 17867 11943 17873
rect 11885 17864 11897 17867
rect 11839 17836 11897 17864
rect 11839 17833 11851 17836
rect 11793 17827 11851 17833
rect 11885 17833 11897 17836
rect 11931 17833 11943 17867
rect 11885 17827 11943 17833
rect 12069 17867 12127 17873
rect 12069 17833 12081 17867
rect 12115 17864 12127 17867
rect 12342 17864 12348 17876
rect 12115 17836 12348 17864
rect 12115 17833 12127 17836
rect 12069 17827 12127 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 13722 17864 13728 17876
rect 13679 17836 13728 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14001 17867 14059 17873
rect 14001 17833 14013 17867
rect 14047 17864 14059 17867
rect 14274 17864 14280 17876
rect 14047 17836 14280 17864
rect 14047 17833 14059 17836
rect 14001 17827 14059 17833
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 16574 17824 16580 17876
rect 16632 17864 16638 17876
rect 17221 17867 17279 17873
rect 17221 17864 17233 17867
rect 16632 17836 17233 17864
rect 16632 17824 16638 17836
rect 17221 17833 17233 17836
rect 17267 17833 17279 17867
rect 17221 17827 17279 17833
rect 17681 17867 17739 17873
rect 17681 17833 17693 17867
rect 17727 17864 17739 17867
rect 17862 17864 17868 17876
rect 17727 17836 17868 17864
rect 17727 17833 17739 17836
rect 17681 17827 17739 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 19150 17864 19156 17876
rect 19111 17836 19156 17864
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 22925 17867 22983 17873
rect 22925 17833 22937 17867
rect 22971 17864 22983 17867
rect 23198 17864 23204 17876
rect 22971 17836 23204 17864
rect 22971 17833 22983 17836
rect 22925 17827 22983 17833
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 23934 17864 23940 17876
rect 23895 17836 23940 17864
rect 23934 17824 23940 17836
rect 23992 17824 23998 17876
rect 24397 17867 24455 17873
rect 24397 17833 24409 17867
rect 24443 17864 24455 17867
rect 24670 17864 24676 17876
rect 24443 17836 24676 17864
rect 24443 17833 24455 17836
rect 24397 17827 24455 17833
rect 24670 17824 24676 17836
rect 24728 17824 24734 17876
rect 25222 17824 25228 17876
rect 25280 17864 25286 17876
rect 25317 17867 25375 17873
rect 25317 17864 25329 17867
rect 25280 17836 25329 17864
rect 25280 17824 25286 17836
rect 25317 17833 25329 17836
rect 25363 17833 25375 17867
rect 25317 17827 25375 17833
rect 11609 17799 11667 17805
rect 11609 17765 11621 17799
rect 11655 17796 11667 17799
rect 12158 17796 12164 17808
rect 11655 17768 12164 17796
rect 11655 17765 11667 17768
rect 11609 17759 11667 17765
rect 12158 17756 12164 17768
rect 12216 17796 12222 17808
rect 12437 17799 12495 17805
rect 12437 17796 12449 17799
rect 12216 17768 12449 17796
rect 12216 17756 12222 17768
rect 12437 17765 12449 17768
rect 12483 17765 12495 17799
rect 12437 17759 12495 17765
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 16206 17796 16212 17808
rect 13872 17768 16212 17796
rect 13872 17756 13878 17768
rect 8573 17731 8631 17737
rect 8573 17697 8585 17731
rect 8619 17728 8631 17731
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 8619 17700 10057 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 10045 17697 10057 17700
rect 10091 17728 10103 17731
rect 10502 17728 10508 17740
rect 10091 17700 10508 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10502 17688 10508 17700
rect 10560 17688 10566 17740
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17728 11851 17731
rect 12529 17731 12587 17737
rect 12529 17728 12541 17731
rect 11839 17700 12541 17728
rect 11839 17697 11851 17700
rect 11793 17691 11851 17697
rect 12529 17697 12541 17700
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17728 13599 17731
rect 14090 17728 14096 17740
rect 13587 17700 14096 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 15304 17737 15332 17768
rect 16206 17756 16212 17768
rect 16264 17756 16270 17808
rect 22094 17796 22100 17808
rect 20916 17768 22100 17796
rect 15562 17737 15568 17740
rect 15289 17731 15347 17737
rect 15289 17697 15301 17731
rect 15335 17697 15347 17731
rect 15556 17728 15568 17737
rect 15523 17700 15568 17728
rect 15289 17691 15347 17697
rect 15556 17691 15568 17700
rect 15562 17688 15568 17691
rect 15620 17688 15626 17740
rect 18040 17731 18098 17737
rect 18040 17728 18052 17731
rect 16684 17700 18052 17728
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 10008 17632 10149 17660
rect 10008 17620 10014 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 12710 17660 12716 17672
rect 12623 17632 12716 17660
rect 10229 17623 10287 17629
rect 9677 17595 9735 17601
rect 9677 17561 9689 17595
rect 9723 17592 9735 17595
rect 10042 17592 10048 17604
rect 9723 17564 10048 17592
rect 9723 17561 9735 17564
rect 9677 17555 9735 17561
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 9398 17484 9404 17536
rect 9456 17524 9462 17536
rect 10244 17524 10272 17623
rect 12710 17620 12716 17632
rect 12768 17660 12774 17672
rect 13354 17660 13360 17672
rect 12768 17632 13360 17660
rect 12768 17620 12774 17632
rect 13354 17620 13360 17632
rect 13412 17660 13418 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13412 17632 14197 17660
rect 13412 17620 13418 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14918 17660 14924 17672
rect 14831 17632 14924 17660
rect 14185 17623 14243 17629
rect 14090 17552 14096 17604
rect 14148 17592 14154 17604
rect 14844 17592 14872 17632
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 16684 17604 16712 17700
rect 18040 17697 18052 17700
rect 18086 17728 18098 17731
rect 19058 17728 19064 17740
rect 18086 17700 19064 17728
rect 18086 17697 18098 17700
rect 18040 17691 18098 17697
rect 19058 17688 19064 17700
rect 19116 17688 19122 17740
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 20441 17731 20499 17737
rect 20441 17728 20453 17731
rect 19484 17700 20453 17728
rect 19484 17688 19490 17700
rect 20441 17697 20453 17700
rect 20487 17697 20499 17731
rect 20441 17691 20499 17697
rect 20916 17669 20944 17768
rect 22094 17756 22100 17768
rect 22152 17796 22158 17808
rect 22554 17796 22560 17808
rect 22152 17768 22560 17796
rect 22152 17756 22158 17768
rect 22554 17756 22560 17768
rect 22612 17756 22618 17808
rect 21174 17737 21180 17740
rect 21168 17728 21180 17737
rect 21135 17700 21180 17728
rect 21168 17691 21180 17700
rect 21174 17688 21180 17691
rect 21232 17688 21238 17740
rect 24026 17688 24032 17740
rect 24084 17728 24090 17740
rect 24305 17731 24363 17737
rect 24305 17728 24317 17731
rect 24084 17700 24317 17728
rect 24084 17688 24090 17700
rect 24305 17697 24317 17700
rect 24351 17728 24363 17731
rect 25590 17728 25596 17740
rect 24351 17700 25596 17728
rect 24351 17697 24363 17700
rect 24305 17691 24363 17697
rect 25590 17688 25596 17700
rect 25648 17688 25654 17740
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17629 17831 17663
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 17773 17623 17831 17629
rect 20272 17632 20913 17660
rect 16666 17592 16672 17604
rect 14148 17564 14872 17592
rect 16579 17564 16672 17592
rect 14148 17552 14154 17564
rect 16666 17552 16672 17564
rect 16724 17552 16730 17604
rect 13170 17524 13176 17536
rect 9456 17496 10272 17524
rect 13131 17496 13176 17524
rect 9456 17484 9462 17496
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 17788 17524 17816 17623
rect 19518 17524 19524 17536
rect 17788 17496 19524 17524
rect 19518 17484 19524 17496
rect 19576 17524 19582 17536
rect 20272 17533 20300 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 24210 17620 24216 17672
rect 24268 17660 24274 17672
rect 24489 17663 24547 17669
rect 24489 17660 24501 17663
rect 24268 17632 24501 17660
rect 24268 17620 24274 17632
rect 24489 17629 24501 17632
rect 24535 17629 24547 17663
rect 24489 17623 24547 17629
rect 25041 17595 25099 17601
rect 25041 17561 25053 17595
rect 25087 17592 25099 17595
rect 25406 17592 25412 17604
rect 25087 17564 25412 17592
rect 25087 17561 25099 17564
rect 25041 17555 25099 17561
rect 25406 17552 25412 17564
rect 25464 17552 25470 17604
rect 19797 17527 19855 17533
rect 19797 17524 19809 17527
rect 19576 17496 19809 17524
rect 19576 17484 19582 17496
rect 19797 17493 19809 17496
rect 19843 17524 19855 17527
rect 20257 17527 20315 17533
rect 20257 17524 20269 17527
rect 19843 17496 20269 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20257 17493 20269 17496
rect 20303 17493 20315 17527
rect 22278 17524 22284 17536
rect 22239 17496 22284 17524
rect 20257 17487 20315 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 23290 17524 23296 17536
rect 23203 17496 23296 17524
rect 23290 17484 23296 17496
rect 23348 17524 23354 17536
rect 23750 17524 23756 17536
rect 23348 17496 23756 17524
rect 23348 17484 23354 17496
rect 23750 17484 23756 17496
rect 23808 17484 23814 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9490 17320 9496 17332
rect 9171 17292 9496 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 9490 17280 9496 17292
rect 9548 17280 9554 17332
rect 10502 17320 10508 17332
rect 10463 17292 10508 17320
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 11609 17323 11667 17329
rect 11609 17289 11621 17323
rect 11655 17320 11667 17323
rect 12710 17320 12716 17332
rect 11655 17292 12716 17320
rect 11655 17289 11667 17292
rect 11609 17283 11667 17289
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 14093 17323 14151 17329
rect 14093 17289 14105 17323
rect 14139 17320 14151 17323
rect 14274 17320 14280 17332
rect 14139 17292 14280 17320
rect 14139 17289 14151 17292
rect 14093 17283 14151 17289
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 15197 17323 15255 17329
rect 15197 17289 15209 17323
rect 15243 17320 15255 17323
rect 15286 17320 15292 17332
rect 15243 17292 15292 17320
rect 15243 17289 15255 17292
rect 15197 17283 15255 17289
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 9456 17224 9720 17252
rect 9456 17212 9462 17224
rect 9582 17184 9588 17196
rect 9543 17156 9588 17184
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 9692 17193 9720 17224
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 12069 17255 12127 17261
rect 12069 17252 12081 17255
rect 11480 17224 12081 17252
rect 11480 17212 11486 17224
rect 12069 17221 12081 17224
rect 12115 17252 12127 17255
rect 13814 17252 13820 17264
rect 12115 17224 13820 17252
rect 12115 17221 12127 17224
rect 12069 17215 12127 17221
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 9677 17187 9735 17193
rect 9677 17153 9689 17187
rect 9723 17153 9735 17187
rect 10962 17184 10968 17196
rect 10923 17156 10968 17184
rect 9677 17147 9735 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 13170 17184 13176 17196
rect 13131 17156 13176 17184
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17184 14059 17187
rect 14550 17184 14556 17196
rect 14047 17156 14556 17184
rect 14047 17153 14059 17156
rect 14001 17147 14059 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 14734 17184 14740 17196
rect 14695 17156 14740 17184
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 10686 17116 10692 17128
rect 10647 17088 10692 17116
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 12250 17116 12256 17128
rect 12211 17088 12256 17116
rect 12250 17076 12256 17088
rect 12308 17076 12314 17128
rect 12894 17116 12900 17128
rect 12807 17088 12900 17116
rect 12894 17076 12900 17088
rect 12952 17116 12958 17128
rect 14461 17119 14519 17125
rect 12952 17088 13676 17116
rect 12952 17076 12958 17088
rect 9033 17051 9091 17057
rect 9033 17017 9045 17051
rect 9079 17048 9091 17051
rect 9490 17048 9496 17060
rect 9079 17020 9496 17048
rect 9079 17017 9091 17020
rect 9033 17011 9091 17017
rect 9490 17008 9496 17020
rect 9548 17008 9554 17060
rect 11977 17051 12035 17057
rect 11977 17017 11989 17051
rect 12023 17048 12035 17051
rect 12023 17020 13032 17048
rect 12023 17017 12035 17020
rect 11977 17011 12035 17017
rect 13004 16992 13032 17020
rect 13648 16992 13676 17088
rect 14461 17085 14473 17119
rect 14507 17116 14519 17119
rect 15212 17116 15240 17283
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 16117 17323 16175 17329
rect 16117 17289 16129 17323
rect 16163 17320 16175 17323
rect 17862 17320 17868 17332
rect 16163 17292 17868 17320
rect 16163 17289 16175 17292
rect 16117 17283 16175 17289
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19613 17323 19671 17329
rect 19613 17320 19625 17323
rect 19484 17292 19625 17320
rect 19484 17280 19490 17292
rect 19613 17289 19625 17292
rect 19659 17289 19671 17323
rect 19613 17283 19671 17289
rect 23109 17323 23167 17329
rect 23109 17289 23121 17323
rect 23155 17320 23167 17323
rect 24670 17320 24676 17332
rect 23155 17292 24676 17320
rect 23155 17289 23167 17292
rect 23109 17283 23167 17289
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 25590 17320 25596 17332
rect 25551 17292 25596 17320
rect 25590 17280 25596 17292
rect 25648 17280 25654 17332
rect 16025 17255 16083 17261
rect 16025 17221 16037 17255
rect 16071 17252 16083 17255
rect 16071 17224 16712 17252
rect 16071 17221 16083 17224
rect 16025 17215 16083 17221
rect 16684 17196 16712 17224
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16298 17184 16304 17196
rect 15436 17156 16304 17184
rect 15436 17144 15442 17156
rect 16298 17144 16304 17156
rect 16356 17184 16362 17196
rect 16577 17187 16635 17193
rect 16577 17184 16589 17187
rect 16356 17156 16589 17184
rect 16356 17144 16362 17156
rect 16577 17153 16589 17156
rect 16623 17153 16635 17187
rect 16577 17147 16635 17153
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 17494 17184 17500 17196
rect 16724 17156 16769 17184
rect 17407 17156 17500 17184
rect 16724 17144 16730 17156
rect 17494 17144 17500 17156
rect 17552 17184 17558 17196
rect 18690 17184 18696 17196
rect 17552 17156 18696 17184
rect 17552 17144 17558 17156
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 16482 17116 16488 17128
rect 14507 17088 15240 17116
rect 16443 17088 16488 17116
rect 14507 17085 14519 17088
rect 14461 17079 14519 17085
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17116 18475 17119
rect 18506 17116 18512 17128
rect 18463 17088 18512 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 19576 17088 20177 17116
rect 19576 17076 19582 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 22189 17119 22247 17125
rect 22189 17085 22201 17119
rect 22235 17116 22247 17119
rect 22554 17116 22560 17128
rect 22235 17088 22560 17116
rect 22235 17085 22247 17088
rect 22189 17079 22247 17085
rect 22554 17076 22560 17088
rect 22612 17116 22618 17128
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 22612 17088 23673 17116
rect 22612 17076 22618 17088
rect 23661 17085 23673 17088
rect 23707 17116 23719 17119
rect 23750 17116 23756 17128
rect 23707 17088 23756 17116
rect 23707 17085 23719 17088
rect 23661 17079 23719 17085
rect 23750 17076 23756 17088
rect 23808 17116 23814 17128
rect 25498 17116 25504 17128
rect 23808 17088 25504 17116
rect 23808 17076 23814 17088
rect 25498 17076 25504 17088
rect 25556 17076 25562 17128
rect 17865 17051 17923 17057
rect 17865 17017 17877 17051
rect 17911 17048 17923 17051
rect 18138 17048 18144 17060
rect 17911 17020 18144 17048
rect 17911 17017 17923 17020
rect 17865 17011 17923 17017
rect 18138 17008 18144 17020
rect 18196 17048 18202 17060
rect 19242 17048 19248 17060
rect 18196 17020 19248 17048
rect 18196 17008 18202 17020
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 10100 16952 10149 16980
rect 10100 16940 10106 16952
rect 10137 16949 10149 16952
rect 10183 16949 10195 16983
rect 10137 16943 10195 16949
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12529 16983 12587 16989
rect 12529 16980 12541 16983
rect 12492 16952 12541 16980
rect 12492 16940 12498 16952
rect 12529 16949 12541 16952
rect 12575 16949 12587 16983
rect 12986 16980 12992 16992
rect 12947 16952 12992 16980
rect 12529 16943 12587 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 13630 16980 13636 16992
rect 13591 16952 13636 16980
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 15562 16980 15568 16992
rect 15475 16952 15568 16980
rect 15562 16940 15568 16952
rect 15620 16980 15626 16992
rect 16206 16980 16212 16992
rect 15620 16952 16212 16980
rect 15620 16940 15626 16952
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 18046 16980 18052 16992
rect 18007 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 18524 16989 18552 17020
rect 19242 17008 19248 17020
rect 19300 17008 19306 17060
rect 20254 17008 20260 17060
rect 20312 17048 20318 17060
rect 23934 17057 23940 17060
rect 20410 17051 20468 17057
rect 20410 17048 20422 17051
rect 20312 17020 20422 17048
rect 20312 17008 20318 17020
rect 20410 17017 20422 17020
rect 20456 17017 20468 17051
rect 23928 17048 23940 17057
rect 23895 17020 23940 17048
rect 20410 17011 20468 17017
rect 23928 17011 23940 17020
rect 23934 17008 23940 17011
rect 23992 17008 23998 17060
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16949 18567 16983
rect 19058 16980 19064 16992
rect 19019 16952 19064 16980
rect 18509 16943 18567 16949
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 20070 16980 20076 16992
rect 20031 16952 20076 16980
rect 20070 16940 20076 16952
rect 20128 16980 20134 16992
rect 21174 16980 21180 16992
rect 20128 16952 21180 16980
rect 20128 16940 20134 16952
rect 21174 16940 21180 16952
rect 21232 16980 21238 16992
rect 21545 16983 21603 16989
rect 21545 16980 21557 16983
rect 21232 16952 21557 16980
rect 21232 16940 21238 16952
rect 21545 16949 21557 16952
rect 21591 16949 21603 16983
rect 23474 16980 23480 16992
rect 23435 16952 23480 16980
rect 21545 16943 21603 16949
rect 23474 16940 23480 16952
rect 23532 16980 23538 16992
rect 24210 16980 24216 16992
rect 23532 16952 24216 16980
rect 23532 16940 23538 16952
rect 24210 16940 24216 16952
rect 24268 16980 24274 16992
rect 25041 16983 25099 16989
rect 25041 16980 25053 16983
rect 24268 16952 25053 16980
rect 24268 16940 24274 16952
rect 25041 16949 25053 16952
rect 25087 16949 25099 16983
rect 25041 16943 25099 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 9217 16779 9275 16785
rect 9217 16745 9229 16779
rect 9263 16776 9275 16779
rect 9398 16776 9404 16788
rect 9263 16748 9404 16776
rect 9263 16745 9275 16748
rect 9217 16739 9275 16745
rect 9398 16736 9404 16748
rect 9456 16776 9462 16788
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9456 16748 9873 16776
rect 9456 16736 9462 16748
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 12805 16779 12863 16785
rect 12805 16776 12817 16779
rect 12768 16748 12817 16776
rect 12768 16736 12774 16748
rect 12805 16745 12817 16748
rect 12851 16745 12863 16779
rect 12805 16739 12863 16745
rect 13446 16736 13452 16788
rect 13504 16776 13510 16788
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13504 16748 13645 16776
rect 13504 16736 13510 16748
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 14734 16776 14740 16788
rect 14695 16748 14740 16776
rect 13633 16739 13691 16745
rect 14734 16736 14740 16748
rect 14792 16736 14798 16788
rect 16298 16776 16304 16788
rect 16259 16748 16304 16776
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16540 16748 16681 16776
rect 16540 16736 16546 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 16853 16779 16911 16785
rect 16853 16745 16865 16779
rect 16899 16776 16911 16779
rect 18138 16776 18144 16788
rect 16899 16748 18144 16776
rect 16899 16745 16911 16748
rect 16853 16739 16911 16745
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18414 16776 18420 16788
rect 18375 16748 18420 16776
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 20254 16776 20260 16788
rect 20215 16748 20260 16776
rect 20254 16736 20260 16748
rect 20312 16776 20318 16788
rect 21818 16776 21824 16788
rect 20312 16748 21824 16776
rect 20312 16736 20318 16748
rect 21818 16736 21824 16748
rect 21876 16776 21882 16788
rect 21913 16779 21971 16785
rect 21913 16776 21925 16779
rect 21876 16748 21925 16776
rect 21876 16736 21882 16748
rect 21913 16745 21925 16748
rect 21959 16745 21971 16779
rect 21913 16739 21971 16745
rect 22094 16736 22100 16788
rect 22152 16736 22158 16788
rect 22462 16776 22468 16788
rect 22423 16748 22468 16776
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 24026 16776 24032 16788
rect 23987 16748 24032 16776
rect 24026 16736 24032 16748
rect 24084 16736 24090 16788
rect 24486 16776 24492 16788
rect 24447 16748 24492 16776
rect 24486 16736 24492 16748
rect 24544 16736 24550 16788
rect 14185 16711 14243 16717
rect 14185 16677 14197 16711
rect 14231 16708 14243 16711
rect 14458 16708 14464 16720
rect 14231 16680 14464 16708
rect 14231 16677 14243 16680
rect 14185 16671 14243 16677
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 15105 16711 15163 16717
rect 15105 16677 15117 16711
rect 15151 16708 15163 16711
rect 17313 16711 17371 16717
rect 15151 16680 15792 16708
rect 15151 16677 15163 16680
rect 15105 16671 15163 16677
rect 15764 16652 15792 16680
rect 17313 16677 17325 16711
rect 17359 16708 17371 16711
rect 17586 16708 17592 16720
rect 17359 16680 17592 16708
rect 17359 16677 17371 16680
rect 17313 16671 17371 16677
rect 17586 16668 17592 16680
rect 17644 16668 17650 16720
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 18877 16711 18935 16717
rect 18877 16708 18889 16711
rect 18104 16680 18889 16708
rect 18104 16668 18110 16680
rect 18877 16677 18889 16680
rect 18923 16708 18935 16711
rect 18966 16708 18972 16720
rect 18923 16680 18972 16708
rect 18923 16677 18935 16680
rect 18877 16671 18935 16677
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 22112 16708 22140 16736
rect 23753 16711 23811 16717
rect 22112 16680 22784 16708
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16640 11391 16643
rect 11422 16640 11428 16652
rect 11379 16612 11428 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11698 16649 11704 16652
rect 11692 16640 11704 16649
rect 11659 16612 11704 16640
rect 11692 16603 11704 16612
rect 11698 16600 11704 16603
rect 11756 16600 11762 16652
rect 13906 16640 13912 16652
rect 13867 16612 13912 16640
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15620 16612 15669 16640
rect 15620 16600 15626 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 15804 16612 15849 16640
rect 15804 16600 15810 16612
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16724 16612 17233 16640
rect 16724 16600 16730 16612
rect 17221 16609 17233 16612
rect 17267 16609 17279 16643
rect 17221 16603 17279 16609
rect 18138 16600 18144 16652
rect 18196 16640 18202 16652
rect 18785 16643 18843 16649
rect 18785 16640 18797 16643
rect 18196 16612 18797 16640
rect 18196 16600 18202 16612
rect 18785 16609 18797 16612
rect 18831 16609 18843 16643
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 18785 16603 18843 16609
rect 19260 16612 19809 16640
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 17494 16572 17500 16584
rect 17455 16544 17500 16572
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16572 18107 16575
rect 18506 16572 18512 16584
rect 18095 16544 18512 16572
rect 18095 16541 18107 16544
rect 18049 16535 18107 16541
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 19058 16572 19064 16584
rect 19019 16544 19064 16572
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 10873 16507 10931 16513
rect 10873 16473 10885 16507
rect 10919 16504 10931 16507
rect 10919 16476 11468 16504
rect 10919 16473 10931 16476
rect 10873 16467 10931 16473
rect 11440 16448 11468 16476
rect 18414 16464 18420 16516
rect 18472 16504 18478 16516
rect 19260 16504 19288 16612
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 21266 16640 21272 16652
rect 21227 16612 21272 16640
rect 19797 16603 19855 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21361 16643 21419 16649
rect 21361 16609 21373 16643
rect 21407 16640 21419 16643
rect 21634 16640 21640 16652
rect 21407 16612 21640 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 22152 16612 22293 16640
rect 22152 16600 22158 16612
rect 22281 16609 22293 16612
rect 22327 16609 22339 16643
rect 22281 16603 22339 16609
rect 22756 16584 22784 16680
rect 23753 16677 23765 16711
rect 23799 16708 23811 16711
rect 23934 16708 23940 16720
rect 23799 16680 23940 16708
rect 23799 16677 23811 16680
rect 23753 16671 23811 16677
rect 23934 16668 23940 16680
rect 23992 16708 23998 16720
rect 25222 16708 25228 16720
rect 23992 16680 25228 16708
rect 23992 16668 23998 16680
rect 22833 16643 22891 16649
rect 22833 16609 22845 16643
rect 22879 16640 22891 16643
rect 23106 16640 23112 16652
rect 22879 16612 23112 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 24394 16640 24400 16652
rect 24355 16612 24400 16640
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 21450 16572 21456 16584
rect 21411 16544 21456 16572
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 22738 16532 22744 16584
rect 22796 16572 22802 16584
rect 22925 16575 22983 16581
rect 22925 16572 22937 16575
rect 22796 16544 22937 16572
rect 22796 16532 22802 16544
rect 22925 16541 22937 16544
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 23014 16532 23020 16584
rect 23072 16572 23078 16584
rect 24596 16581 24624 16680
rect 25222 16668 25228 16680
rect 25280 16668 25286 16720
rect 25041 16643 25099 16649
rect 25041 16640 25053 16643
rect 24780 16612 25053 16640
rect 24581 16575 24639 16581
rect 23072 16544 23117 16572
rect 23072 16532 23078 16544
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24780 16572 24808 16612
rect 25041 16609 25053 16612
rect 25087 16609 25099 16643
rect 25498 16640 25504 16652
rect 25411 16612 25504 16640
rect 25041 16603 25099 16609
rect 25498 16600 25504 16612
rect 25556 16640 25562 16652
rect 26142 16640 26148 16652
rect 25556 16612 26148 16640
rect 25556 16600 25562 16612
rect 26142 16600 26148 16612
rect 26200 16600 26206 16652
rect 24581 16535 24639 16541
rect 24688 16544 24808 16572
rect 18472 16476 19288 16504
rect 18472 16464 18478 16476
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 24688 16504 24716 16544
rect 24176 16476 24716 16504
rect 24176 16464 24182 16476
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 12710 16436 12716 16448
rect 11480 16408 12716 16436
rect 11480 16396 11486 16408
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 15289 16439 15347 16445
rect 15289 16405 15301 16439
rect 15335 16436 15347 16439
rect 15470 16436 15476 16448
rect 15335 16408 15476 16436
rect 15335 16405 15347 16408
rect 15289 16399 15347 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 18506 16396 18512 16448
rect 18564 16436 18570 16448
rect 19429 16439 19487 16445
rect 19429 16436 19441 16439
rect 18564 16408 19441 16436
rect 18564 16396 18570 16408
rect 19429 16405 19441 16408
rect 19475 16405 19487 16439
rect 20530 16436 20536 16448
rect 20491 16408 20536 16436
rect 19429 16399 19487 16405
rect 20530 16396 20536 16408
rect 20588 16396 20594 16448
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 20901 16439 20959 16445
rect 20901 16436 20913 16439
rect 20772 16408 20913 16436
rect 20772 16396 20778 16408
rect 20901 16405 20913 16408
rect 20947 16405 20959 16439
rect 20901 16399 20959 16405
rect 23566 16396 23572 16448
rect 23624 16436 23630 16448
rect 23842 16436 23848 16448
rect 23624 16408 23848 16436
rect 23624 16396 23630 16408
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11756 16204 11805 16232
rect 11756 16192 11762 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 15378 16232 15384 16244
rect 15339 16204 15384 16232
rect 11793 16195 11851 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 17402 16192 17408 16244
rect 17460 16232 17466 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17460 16204 17509 16232
rect 17460 16192 17466 16204
rect 17497 16201 17509 16204
rect 17543 16232 17555 16235
rect 17586 16232 17592 16244
rect 17543 16204 17592 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 18012 16204 18061 16232
rect 18012 16192 18018 16204
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 19058 16232 19064 16244
rect 19019 16204 19064 16232
rect 18049 16195 18107 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 24026 16232 24032 16244
rect 23523 16204 24032 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 24670 16232 24676 16244
rect 24631 16204 24676 16232
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 25133 16235 25191 16241
rect 25133 16201 25145 16235
rect 25179 16232 25191 16235
rect 25222 16232 25228 16244
rect 25179 16204 25228 16232
rect 25179 16201 25191 16204
rect 25133 16195 25191 16201
rect 25222 16192 25228 16204
rect 25280 16192 25286 16244
rect 12437 16167 12495 16173
rect 12437 16133 12449 16167
rect 12483 16164 12495 16167
rect 13906 16164 13912 16176
rect 12483 16136 13912 16164
rect 12483 16133 12495 16136
rect 12437 16127 12495 16133
rect 13906 16124 13912 16136
rect 13964 16124 13970 16176
rect 20530 16124 20536 16176
rect 20588 16164 20594 16176
rect 21637 16167 21695 16173
rect 21637 16164 21649 16167
rect 20588 16136 21649 16164
rect 20588 16124 20594 16136
rect 21637 16133 21649 16136
rect 21683 16133 21695 16167
rect 21637 16127 21695 16133
rect 23290 16124 23296 16176
rect 23348 16164 23354 16176
rect 23661 16167 23719 16173
rect 23661 16164 23673 16167
rect 23348 16136 23673 16164
rect 23348 16124 23354 16136
rect 23661 16133 23673 16136
rect 23707 16133 23719 16167
rect 23661 16127 23719 16133
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 11422 16096 11428 16108
rect 10367 16068 11284 16096
rect 11383 16068 11428 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 11146 16028 11152 16040
rect 10735 16000 11152 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 11256 16037 11284 16068
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 12986 16096 12992 16108
rect 12947 16068 12992 16096
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 13814 16056 13820 16108
rect 13872 16096 13878 16108
rect 13998 16096 14004 16108
rect 13872 16068 14004 16096
rect 13872 16056 13878 16068
rect 13998 16056 14004 16068
rect 14056 16056 14062 16108
rect 16206 16096 16212 16108
rect 16119 16068 16212 16096
rect 16206 16056 16212 16068
rect 16264 16096 16270 16108
rect 17494 16096 17500 16108
rect 16264 16068 17500 16096
rect 16264 16056 16270 16068
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 18601 16099 18659 16105
rect 18601 16096 18613 16099
rect 17972 16068 18613 16096
rect 11241 16031 11299 16037
rect 11241 15997 11253 16031
rect 11287 16028 11299 16031
rect 12342 16028 12348 16040
rect 11287 16000 12348 16028
rect 11287 15997 11299 16000
rect 11241 15991 11299 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 14274 16037 14280 16040
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 14268 16028 14280 16037
rect 13955 16000 14280 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 14268 15991 14280 16000
rect 14274 15988 14280 15991
rect 14332 15988 14338 16040
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16356 16000 16681 16028
rect 16356 15988 16362 16000
rect 16669 15997 16681 16000
rect 16715 16028 16727 16031
rect 17862 16028 17868 16040
rect 16715 16000 17868 16028
rect 16715 15997 16727 16000
rect 16669 15991 16727 15997
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 16942 15960 16948 15972
rect 10796 15932 12940 15960
rect 16903 15932 16948 15960
rect 9950 15892 9956 15904
rect 9911 15864 9956 15892
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10796 15901 10824 15932
rect 10781 15895 10839 15901
rect 10781 15861 10793 15895
rect 10827 15861 10839 15895
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 10781 15855 10839 15861
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 12032 15864 12173 15892
rect 12032 15852 12038 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 12802 15892 12808 15904
rect 12763 15864 12808 15892
rect 12161 15855 12219 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 12912 15901 12940 15932
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 17972 15960 18000 16068
rect 18601 16065 18613 16068
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16096 20039 16099
rect 20070 16096 20076 16108
rect 20027 16068 20076 16096
rect 20027 16065 20039 16068
rect 19981 16059 20039 16065
rect 20070 16056 20076 16068
rect 20128 16096 20134 16108
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 20128 16068 20637 16096
rect 20128 16056 20134 16068
rect 20625 16065 20637 16068
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 21818 16056 21824 16108
rect 21876 16096 21882 16108
rect 22189 16099 22247 16105
rect 22189 16096 22201 16099
rect 21876 16068 22201 16096
rect 21876 16056 21882 16068
rect 22189 16065 22201 16068
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 23750 16056 23756 16108
rect 23808 16096 23814 16108
rect 24305 16099 24363 16105
rect 24305 16096 24317 16099
rect 23808 16068 24317 16096
rect 23808 16056 23814 16068
rect 24305 16065 24317 16068
rect 24351 16096 24363 16099
rect 24578 16096 24584 16108
rect 24351 16068 24584 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 20441 16031 20499 16037
rect 20441 15997 20453 16031
rect 20487 16028 20499 16031
rect 20530 16028 20536 16040
rect 20487 16000 20536 16028
rect 20487 15997 20499 16000
rect 20441 15991 20499 15997
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 24026 16028 24032 16040
rect 23987 16000 24032 16028
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 25222 16028 25228 16040
rect 25183 16000 25228 16028
rect 25222 15988 25228 16000
rect 25280 16028 25286 16040
rect 25961 16031 26019 16037
rect 25961 16028 25973 16031
rect 25280 16000 25973 16028
rect 25280 15988 25286 16000
rect 25961 15997 25973 16000
rect 26007 15997 26019 16031
rect 25961 15991 26019 15997
rect 17788 15932 18000 15960
rect 19613 15963 19671 15969
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 12943 15864 13461 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 16577 15895 16635 15901
rect 16577 15861 16589 15895
rect 16623 15892 16635 15895
rect 16666 15892 16672 15904
rect 16623 15864 16672 15892
rect 16623 15861 16635 15864
rect 16577 15855 16635 15861
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 17788 15901 17816 15932
rect 19613 15929 19625 15963
rect 19659 15960 19671 15963
rect 21177 15963 21235 15969
rect 19659 15932 20576 15960
rect 19659 15929 19671 15932
rect 19613 15923 19671 15929
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 16816 15864 17785 15892
rect 16816 15852 16822 15864
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 18414 15892 18420 15904
rect 18375 15864 18420 15892
rect 17773 15855 17831 15861
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 18506 15852 18512 15904
rect 18564 15892 18570 15904
rect 20070 15892 20076 15904
rect 18564 15864 18609 15892
rect 20031 15864 20076 15892
rect 18564 15852 18570 15864
rect 20070 15852 20076 15864
rect 20128 15852 20134 15904
rect 20548 15901 20576 15932
rect 21177 15929 21189 15963
rect 21223 15960 21235 15963
rect 21634 15960 21640 15972
rect 21223 15932 21640 15960
rect 21223 15929 21235 15932
rect 21177 15923 21235 15929
rect 21634 15920 21640 15932
rect 21692 15920 21698 15972
rect 21726 15920 21732 15972
rect 21784 15960 21790 15972
rect 22094 15960 22100 15972
rect 21784 15932 22100 15960
rect 21784 15920 21790 15932
rect 22094 15920 22100 15932
rect 22152 15960 22158 15972
rect 25498 15960 25504 15972
rect 22152 15932 22245 15960
rect 25459 15932 25504 15960
rect 22152 15920 22158 15932
rect 25498 15920 25504 15932
rect 25556 15920 25562 15972
rect 20533 15895 20591 15901
rect 20533 15861 20545 15895
rect 20579 15892 20591 15895
rect 20898 15892 20904 15904
rect 20579 15864 20904 15892
rect 20579 15861 20591 15864
rect 20533 15855 20591 15861
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 21266 15852 21272 15904
rect 21324 15892 21330 15904
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 21324 15864 21465 15892
rect 21324 15852 21330 15864
rect 21453 15861 21465 15864
rect 21499 15861 21511 15895
rect 21453 15855 21511 15861
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 21968 15864 22017 15892
rect 21968 15852 21974 15864
rect 22005 15861 22017 15864
rect 22051 15861 22063 15895
rect 22738 15892 22744 15904
rect 22699 15864 22744 15892
rect 22005 15855 22063 15861
rect 22738 15852 22744 15864
rect 22796 15852 22802 15904
rect 23106 15892 23112 15904
rect 23067 15864 23112 15892
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 24118 15892 24124 15904
rect 24079 15864 24124 15892
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11204 15660 11735 15688
rect 11204 15648 11210 15660
rect 11241 15623 11299 15629
rect 11241 15589 11253 15623
rect 11287 15620 11299 15623
rect 11422 15620 11428 15632
rect 11287 15592 11428 15620
rect 11287 15589 11299 15592
rect 11241 15583 11299 15589
rect 11422 15580 11428 15592
rect 11480 15620 11486 15632
rect 11578 15623 11636 15629
rect 11578 15620 11590 15623
rect 11480 15592 11590 15620
rect 11480 15580 11486 15592
rect 11578 15589 11590 15592
rect 11624 15589 11636 15623
rect 11707 15620 11735 15660
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 12032 15660 12725 15688
rect 12032 15648 12038 15660
rect 12713 15657 12725 15660
rect 12759 15688 12771 15691
rect 12986 15688 12992 15700
rect 12759 15660 12992 15688
rect 12759 15657 12771 15660
rect 12713 15651 12771 15657
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 13964 15660 14657 15688
rect 13964 15648 13970 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 15105 15691 15163 15697
rect 15105 15657 15117 15691
rect 15151 15688 15163 15691
rect 15838 15688 15844 15700
rect 15151 15660 15844 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16298 15688 16304 15700
rect 16259 15660 16304 15688
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16574 15648 16580 15700
rect 16632 15688 16638 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 16632 15660 16773 15688
rect 16632 15648 16638 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 16761 15651 16819 15657
rect 17126 15648 17132 15700
rect 17184 15688 17190 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 17184 15660 17233 15688
rect 17184 15648 17190 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 17221 15651 17279 15657
rect 17957 15691 18015 15697
rect 17957 15657 17969 15691
rect 18003 15688 18015 15691
rect 18138 15688 18144 15700
rect 18003 15660 18144 15688
rect 18003 15657 18015 15660
rect 17957 15651 18015 15657
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 18325 15691 18383 15697
rect 18325 15657 18337 15691
rect 18371 15688 18383 15691
rect 18782 15688 18788 15700
rect 18371 15660 18788 15688
rect 18371 15657 18383 15660
rect 18325 15651 18383 15657
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 18966 15688 18972 15700
rect 18927 15660 18972 15688
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 19242 15688 19248 15700
rect 19203 15660 19248 15688
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 20898 15688 20904 15700
rect 20859 15660 20904 15688
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 22465 15691 22523 15697
rect 22465 15657 22477 15691
rect 22511 15688 22523 15691
rect 23014 15688 23020 15700
rect 22511 15660 23020 15688
rect 22511 15657 22523 15660
rect 22465 15651 22523 15657
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 24210 15648 24216 15700
rect 24268 15688 24274 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 24268 15660 24501 15688
rect 24268 15648 24274 15660
rect 24489 15657 24501 15660
rect 24535 15657 24547 15691
rect 24489 15651 24547 15657
rect 24578 15648 24584 15700
rect 24636 15688 24642 15700
rect 24857 15691 24915 15697
rect 24857 15688 24869 15691
rect 24636 15660 24869 15688
rect 24636 15648 24642 15660
rect 24857 15657 24869 15660
rect 24903 15657 24915 15691
rect 24857 15651 24915 15657
rect 13078 15620 13084 15632
rect 11707 15592 13084 15620
rect 11578 15583 11636 15589
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 14182 15620 14188 15632
rect 14143 15592 14188 15620
rect 14182 15580 14188 15592
rect 14240 15580 14246 15632
rect 15654 15580 15660 15632
rect 15712 15620 15718 15632
rect 15749 15623 15807 15629
rect 15749 15620 15761 15623
rect 15712 15592 15761 15620
rect 15712 15580 15718 15592
rect 15749 15589 15761 15592
rect 15795 15589 15807 15623
rect 20717 15623 20775 15629
rect 20717 15620 20729 15623
rect 15749 15583 15807 15589
rect 19904 15592 20729 15620
rect 11330 15552 11336 15564
rect 11291 15524 11336 15552
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 13909 15555 13967 15561
rect 13909 15552 13921 15555
rect 13872 15524 13921 15552
rect 13872 15512 13878 15524
rect 13909 15521 13921 15524
rect 13955 15521 13967 15555
rect 15470 15552 15476 15564
rect 15431 15524 15476 15552
rect 13909 15515 13967 15521
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15552 17187 15555
rect 17218 15552 17224 15564
rect 17175 15524 17224 15552
rect 17175 15521 17187 15524
rect 17129 15515 17187 15521
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 19610 15552 19616 15564
rect 19571 15524 19616 15552
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 19904 15496 19932 15592
rect 20717 15589 20729 15592
rect 20763 15620 20775 15623
rect 21450 15620 21456 15632
rect 20763 15592 21456 15620
rect 20763 15589 20775 15592
rect 20717 15583 20775 15589
rect 21450 15580 21456 15592
rect 21508 15580 21514 15632
rect 24946 15580 24952 15632
rect 25004 15620 25010 15632
rect 25317 15623 25375 15629
rect 25317 15620 25329 15623
rect 25004 15592 25329 15620
rect 25004 15580 25010 15592
rect 25317 15589 25329 15592
rect 25363 15589 25375 15623
rect 25317 15583 25375 15589
rect 20349 15555 20407 15561
rect 20349 15521 20361 15555
rect 20395 15552 20407 15555
rect 20898 15552 20904 15564
rect 20395 15524 20904 15552
rect 20395 15521 20407 15524
rect 20349 15515 20407 15521
rect 20898 15512 20904 15524
rect 20956 15552 20962 15564
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 20956 15524 21281 15552
rect 20956 15512 20962 15524
rect 21269 15521 21281 15524
rect 21315 15521 21327 15555
rect 22554 15552 22560 15564
rect 22515 15524 22560 15552
rect 21269 15515 21327 15521
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 22830 15561 22836 15564
rect 22824 15515 22836 15561
rect 22888 15552 22894 15564
rect 25038 15552 25044 15564
rect 22888 15524 22924 15552
rect 24999 15524 25044 15552
rect 22830 15512 22836 15515
rect 22888 15512 22894 15524
rect 25038 15512 25044 15524
rect 25096 15512 25102 15564
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10962 15484 10968 15496
rect 10367 15456 10968 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 15654 15444 15660 15496
rect 15712 15484 15718 15496
rect 16022 15484 16028 15496
rect 15712 15456 16028 15484
rect 15712 15444 15718 15456
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 17313 15487 17371 15493
rect 17313 15453 17325 15487
rect 17359 15453 17371 15487
rect 19702 15484 19708 15496
rect 19663 15456 19708 15484
rect 17313 15447 17371 15453
rect 10778 15416 10784 15428
rect 10739 15388 10784 15416
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 13817 15419 13875 15425
rect 13817 15385 13829 15419
rect 13863 15416 13875 15419
rect 15562 15416 15568 15428
rect 13863 15388 15568 15416
rect 13863 15385 13875 15388
rect 13817 15379 13875 15385
rect 15562 15376 15568 15388
rect 15620 15376 15626 15428
rect 17328 15416 17356 15447
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 19886 15484 19892 15496
rect 19799 15456 19892 15484
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 20772 15456 21373 15484
rect 20772 15444 20778 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15484 21603 15487
rect 21818 15484 21824 15496
rect 21591 15456 21824 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 16592 15388 17356 15416
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 12802 15348 12808 15360
rect 12492 15320 12808 15348
rect 12492 15308 12498 15320
rect 12802 15308 12808 15320
rect 12860 15348 12866 15360
rect 13265 15351 13323 15357
rect 13265 15348 13277 15351
rect 12860 15320 13277 15348
rect 12860 15308 12866 15320
rect 13265 15317 13277 15320
rect 13311 15317 13323 15351
rect 13265 15311 13323 15317
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 16592 15357 16620 15388
rect 21450 15376 21456 15428
rect 21508 15416 21514 15428
rect 21508 15388 22600 15416
rect 21508 15376 21514 15388
rect 16577 15351 16635 15357
rect 16577 15348 16589 15351
rect 16540 15320 16589 15348
rect 16540 15308 16546 15320
rect 16577 15317 16589 15320
rect 16623 15317 16635 15351
rect 16577 15311 16635 15317
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 17126 15348 17132 15360
rect 16908 15320 17132 15348
rect 16908 15308 16914 15320
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 18690 15348 18696 15360
rect 18651 15320 18696 15348
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 21910 15348 21916 15360
rect 21871 15320 21916 15348
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 22572 15348 22600 15388
rect 23937 15351 23995 15357
rect 23937 15348 23949 15351
rect 22572 15320 23949 15348
rect 23937 15317 23949 15320
rect 23983 15317 23995 15351
rect 23937 15311 23995 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 10870 15144 10876 15156
rect 10827 15116 10876 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11112 15116 11805 15144
rect 11112 15104 11118 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 10321 15079 10379 15085
rect 10321 15045 10333 15079
rect 10367 15076 10379 15079
rect 10367 15048 11376 15076
rect 10367 15045 10379 15048
rect 10321 15039 10379 15045
rect 11348 15020 11376 15048
rect 9950 15008 9956 15020
rect 9863 14980 9956 15008
rect 9950 14968 9956 14980
rect 10008 15008 10014 15020
rect 10778 15008 10784 15020
rect 10008 14980 10784 15008
rect 10008 14968 10014 14980
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 11238 15008 11244 15020
rect 11199 14980 11244 15008
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 11330 14968 11336 15020
rect 11388 15008 11394 15020
rect 11388 14980 11481 15008
rect 11388 14968 11394 14980
rect 11808 14940 11836 15107
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12492 15116 12537 15144
rect 12492 15104 12498 15116
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 14737 15147 14795 15153
rect 14737 15144 14749 15147
rect 13872 15116 14749 15144
rect 13872 15104 13878 15116
rect 14737 15113 14749 15116
rect 14783 15113 14795 15147
rect 14737 15107 14795 15113
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 17276 15116 17325 15144
rect 17276 15104 17282 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17313 15107 17371 15113
rect 18782 15104 18788 15156
rect 18840 15104 18846 15156
rect 21177 15147 21235 15153
rect 21177 15113 21189 15147
rect 21223 15144 21235 15147
rect 21818 15144 21824 15156
rect 21223 15116 21824 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 22370 15144 22376 15156
rect 22331 15116 22376 15144
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 22888 15116 23029 15144
rect 22888 15104 22894 15116
rect 23017 15113 23029 15116
rect 23063 15144 23075 15147
rect 23385 15147 23443 15153
rect 23385 15144 23397 15147
rect 23063 15116 23397 15144
rect 23063 15113 23075 15116
rect 23017 15107 23075 15113
rect 23385 15113 23397 15116
rect 23431 15113 23443 15147
rect 23385 15107 23443 15113
rect 13998 15036 14004 15088
rect 14056 15076 14062 15088
rect 18800 15076 18828 15104
rect 14056 15048 15424 15076
rect 14056 15036 14062 15048
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12768 14980 13001 15008
rect 12768 14968 12774 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 13722 14968 13728 15020
rect 13780 15008 13786 15020
rect 14016 15008 14044 15036
rect 13780 14980 14044 15008
rect 14277 15011 14335 15017
rect 13780 14968 13786 14980
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 14366 15008 14372 15020
rect 14323 14980 14372 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 15396 15017 15424 15048
rect 18616 15048 18828 15076
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 11808 14912 12817 14940
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 13998 14940 14004 14952
rect 13959 14912 14004 14940
rect 12805 14903 12863 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 18616 14949 18644 15048
rect 18690 14968 18696 15020
rect 18748 15008 18754 15020
rect 18785 15011 18843 15017
rect 18785 15008 18797 15011
rect 18748 14980 18797 15008
rect 18748 14968 18754 14980
rect 18785 14977 18797 14980
rect 18831 14977 18843 15011
rect 23400 15008 23428 15107
rect 24854 15104 24860 15156
rect 24912 15144 24918 15156
rect 25409 15147 25467 15153
rect 25409 15144 25421 15147
rect 24912 15116 25421 15144
rect 24912 15104 24918 15116
rect 25409 15113 25421 15116
rect 25455 15113 25467 15147
rect 26234 15144 26240 15156
rect 26195 15116 26240 15144
rect 25409 15107 25467 15113
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 23661 15079 23719 15085
rect 23661 15045 23673 15079
rect 23707 15076 23719 15079
rect 25038 15076 25044 15088
rect 23707 15048 25044 15076
rect 23707 15045 23719 15048
rect 23661 15039 23719 15045
rect 25038 15036 25044 15048
rect 25096 15036 25102 15088
rect 23934 15008 23940 15020
rect 23400 14980 23940 15008
rect 18785 14971 18843 14977
rect 23934 14968 23940 14980
rect 23992 15008 23998 15020
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23992 14980 24225 15008
rect 23992 14968 23998 14980
rect 24213 14977 24225 14980
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 18601 14943 18659 14949
rect 18601 14909 18613 14943
rect 18647 14909 18659 14943
rect 18601 14903 18659 14909
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 19797 14943 19855 14949
rect 19797 14940 19809 14943
rect 19576 14912 19809 14940
rect 19576 14900 19582 14912
rect 19797 14909 19809 14912
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 19886 14900 19892 14952
rect 19944 14940 19950 14952
rect 20053 14943 20111 14949
rect 20053 14940 20065 14943
rect 19944 14912 20065 14940
rect 19944 14900 19950 14912
rect 20053 14909 20065 14912
rect 20099 14909 20111 14943
rect 20053 14903 20111 14909
rect 22370 14900 22376 14952
rect 22428 14940 22434 14952
rect 22465 14943 22523 14949
rect 22465 14940 22477 14943
rect 22428 14912 22477 14940
rect 22428 14900 22434 14912
rect 22465 14909 22477 14912
rect 22511 14909 22523 14943
rect 22465 14903 22523 14909
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 24176 14912 25237 14940
rect 24176 14900 24182 14912
rect 25225 14909 25237 14912
rect 25271 14940 25283 14943
rect 25777 14943 25835 14949
rect 25777 14940 25789 14943
rect 25271 14912 25789 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25777 14909 25789 14912
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 12253 14875 12311 14881
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 12897 14875 12955 14881
rect 12897 14872 12909 14875
rect 12299 14844 12909 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12897 14841 12909 14844
rect 12943 14872 12955 14875
rect 14366 14872 14372 14884
rect 12943 14844 14372 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 15648 14875 15706 14881
rect 15648 14841 15660 14875
rect 15694 14841 15706 14875
rect 15648 14835 15706 14841
rect 17865 14875 17923 14881
rect 17865 14841 17877 14875
rect 17911 14872 17923 14875
rect 18693 14875 18751 14881
rect 18693 14872 18705 14875
rect 17911 14844 18705 14872
rect 17911 14841 17923 14844
rect 17865 14835 17923 14841
rect 18693 14841 18705 14844
rect 18739 14872 18751 14875
rect 18782 14872 18788 14884
rect 18739 14844 18788 14872
rect 18739 14841 18751 14844
rect 18693 14835 18751 14841
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 11146 14804 11152 14816
rect 10735 14776 11152 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11238 14764 11244 14816
rect 11296 14804 11302 14816
rect 12526 14804 12532 14816
rect 11296 14776 12532 14804
rect 11296 14764 11302 14776
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 13906 14804 13912 14816
rect 13771 14776 13912 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15672 14804 15700 14835
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 19337 14875 19395 14881
rect 19337 14841 19349 14875
rect 19383 14872 19395 14875
rect 19610 14872 19616 14884
rect 19383 14844 19616 14872
rect 19383 14841 19395 14844
rect 19337 14835 19395 14841
rect 19610 14832 19616 14844
rect 19668 14832 19674 14884
rect 19702 14832 19708 14884
rect 19760 14872 19766 14884
rect 23014 14872 23020 14884
rect 19760 14844 23020 14872
rect 19760 14832 19766 14844
rect 23014 14832 23020 14844
rect 23072 14832 23078 14884
rect 15746 14804 15752 14816
rect 15335 14776 15752 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15746 14764 15752 14776
rect 15804 14804 15810 14816
rect 16482 14804 16488 14816
rect 15804 14776 16488 14804
rect 15804 14764 15810 14776
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16758 14804 16764 14816
rect 16719 14776 16764 14804
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 18230 14804 18236 14816
rect 18191 14776 18236 14804
rect 18230 14764 18236 14776
rect 18288 14764 18294 14816
rect 22649 14807 22707 14813
rect 22649 14773 22661 14807
rect 22695 14804 22707 14807
rect 23842 14804 23848 14816
rect 22695 14776 23848 14804
rect 22695 14773 22707 14776
rect 22649 14767 22707 14773
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 24026 14804 24032 14816
rect 23987 14776 24032 14804
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 24121 14807 24179 14813
rect 24121 14773 24133 14807
rect 24167 14804 24179 14807
rect 24302 14804 24308 14816
rect 24167 14776 24308 14804
rect 24167 14773 24179 14776
rect 24121 14767 24179 14773
rect 24302 14764 24308 14776
rect 24360 14804 24366 14816
rect 24673 14807 24731 14813
rect 24673 14804 24685 14807
rect 24360 14776 24685 14804
rect 24360 14764 24366 14776
rect 24673 14773 24685 14776
rect 24719 14773 24731 14807
rect 24673 14767 24731 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10778 14600 10784 14612
rect 10643 14572 10784 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10226 14396 10232 14408
rect 10187 14368 10232 14396
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10704 14405 10732 14572
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 12710 14600 12716 14612
rect 12671 14572 12716 14600
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 13998 14600 14004 14612
rect 13679 14572 14004 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 13998 14560 14004 14572
rect 14056 14600 14062 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14056 14572 14657 14600
rect 14056 14560 14062 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 16025 14603 16083 14609
rect 16025 14600 16037 14603
rect 14884 14572 16037 14600
rect 14884 14560 14890 14572
rect 16025 14569 16037 14572
rect 16071 14600 16083 14603
rect 16482 14600 16488 14612
rect 16071 14572 16488 14600
rect 16071 14569 16083 14572
rect 16025 14563 16083 14569
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 18506 14600 18512 14612
rect 18467 14572 18512 14600
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 19889 14603 19947 14609
rect 19889 14569 19901 14603
rect 19935 14600 19947 14603
rect 20438 14600 20444 14612
rect 19935 14572 20444 14600
rect 19935 14569 19947 14572
rect 19889 14563 19947 14569
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 20714 14600 20720 14612
rect 20675 14572 20720 14600
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 20898 14600 20904 14612
rect 20859 14572 20904 14600
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 23934 14600 23940 14612
rect 23895 14572 23940 14600
rect 23934 14560 23940 14572
rect 23992 14560 23998 14612
rect 25225 14603 25283 14609
rect 25225 14569 25237 14603
rect 25271 14600 25283 14603
rect 25314 14600 25320 14612
rect 25271 14572 25320 14600
rect 25271 14569 25283 14572
rect 25225 14563 25283 14569
rect 25314 14560 25320 14572
rect 25372 14560 25378 14612
rect 19337 14535 19395 14541
rect 19337 14501 19349 14535
rect 19383 14532 19395 14535
rect 19978 14532 19984 14544
rect 19383 14504 19984 14532
rect 19383 14501 19395 14504
rect 19337 14495 19395 14501
rect 19978 14492 19984 14504
rect 20036 14532 20042 14544
rect 20257 14535 20315 14541
rect 20257 14532 20269 14535
rect 20036 14504 20269 14532
rect 20036 14492 20042 14504
rect 20257 14501 20269 14504
rect 20303 14501 20315 14535
rect 20257 14495 20315 14501
rect 10778 14424 10784 14476
rect 10836 14464 10842 14476
rect 10945 14467 11003 14473
rect 10945 14464 10957 14467
rect 10836 14436 10957 14464
rect 10836 14424 10842 14436
rect 10945 14433 10957 14436
rect 10991 14464 11003 14467
rect 11974 14464 11980 14476
rect 10991 14436 11980 14464
rect 10991 14433 11003 14436
rect 10945 14427 11003 14433
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 13998 14464 14004 14476
rect 13959 14436 14004 14464
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 15930 14464 15936 14476
rect 15891 14436 15936 14464
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 17385 14467 17443 14473
rect 17385 14464 17397 14467
rect 16776 14436 17397 14464
rect 16776 14408 16804 14436
rect 17385 14433 17397 14436
rect 17431 14464 17443 14467
rect 17954 14464 17960 14476
rect 17431 14436 17960 14464
rect 17431 14433 17443 14436
rect 17385 14427 17443 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19705 14467 19763 14473
rect 19705 14464 19717 14467
rect 19484 14436 19717 14464
rect 19484 14424 19490 14436
rect 19705 14433 19717 14436
rect 19751 14433 19763 14467
rect 21266 14464 21272 14476
rect 21227 14436 21272 14464
rect 19705 14427 19763 14433
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13630 14396 13636 14408
rect 13587 14368 13636 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 13630 14356 13636 14368
rect 13688 14396 13694 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13688 14368 14105 14396
rect 13688 14356 13694 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14274 14396 14280 14408
rect 14235 14368 14280 14396
rect 14093 14359 14151 14365
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 15286 14356 15292 14408
rect 15344 14396 15350 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15344 14368 16129 14396
rect 15344 14356 15350 14368
rect 16117 14365 16129 14368
rect 16163 14396 16175 14399
rect 16758 14396 16764 14408
rect 16163 14368 16764 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 17126 14396 17132 14408
rect 17087 14368 17132 14396
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 19720 14396 19748 14427
rect 21266 14424 21272 14436
rect 21324 14424 21330 14476
rect 22830 14473 22836 14476
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 22824 14464 22836 14473
rect 22143 14436 22836 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 22824 14427 22836 14436
rect 22830 14424 22836 14427
rect 22888 14424 22894 14476
rect 25038 14464 25044 14476
rect 24999 14436 25044 14464
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 20254 14396 20260 14408
rect 19720 14368 20260 14396
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20956 14368 21373 14396
rect 20956 14356 20962 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 22557 14399 22615 14405
rect 21508 14368 21553 14396
rect 21508 14356 21514 14368
rect 22557 14365 22569 14399
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 15562 14328 15568 14340
rect 15523 14300 15568 14328
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 12066 14260 12072 14272
rect 12027 14232 12072 14260
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14240 14232 15025 14260
rect 14240 14220 14246 14232
rect 15013 14229 15025 14232
rect 15059 14260 15071 14263
rect 16482 14260 16488 14272
rect 15059 14232 16488 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 16482 14220 16488 14232
rect 16540 14220 16546 14272
rect 16850 14260 16856 14272
rect 16811 14232 16856 14260
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 22465 14263 22523 14269
rect 22465 14229 22477 14263
rect 22511 14260 22523 14263
rect 22572 14260 22600 14359
rect 23934 14288 23940 14340
rect 23992 14328 23998 14340
rect 23992 14300 24992 14328
rect 23992 14288 23998 14300
rect 23952 14260 23980 14288
rect 22511 14232 23980 14260
rect 22511 14229 22523 14232
rect 22465 14223 22523 14229
rect 24026 14220 24032 14272
rect 24084 14260 24090 14272
rect 24964 14269 24992 14300
rect 24489 14263 24547 14269
rect 24489 14260 24501 14263
rect 24084 14232 24501 14260
rect 24084 14220 24090 14232
rect 24489 14229 24501 14232
rect 24535 14229 24547 14263
rect 24489 14223 24547 14229
rect 24949 14263 25007 14269
rect 24949 14229 24961 14263
rect 24995 14260 25007 14263
rect 26050 14260 26056 14272
rect 24995 14232 26056 14260
rect 24995 14229 25007 14232
rect 24949 14223 25007 14229
rect 26050 14220 26056 14232
rect 26108 14220 26114 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 10321 14059 10379 14065
rect 10321 14025 10333 14059
rect 10367 14056 10379 14059
rect 10778 14056 10784 14068
rect 10367 14028 10784 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11388 14028 12173 14056
rect 11388 14016 11394 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 12805 14059 12863 14065
rect 12805 14025 12817 14059
rect 12851 14056 12863 14059
rect 13446 14056 13452 14068
rect 12851 14028 13452 14056
rect 12851 14025 12863 14028
rect 12805 14019 12863 14025
rect 12176 13988 12204 14019
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13722 14016 13728 14068
rect 13780 14016 13786 14068
rect 13998 14016 14004 14068
rect 14056 14056 14062 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 14056 14028 16129 14056
rect 14056 14016 14062 14028
rect 16117 14025 16129 14028
rect 16163 14025 16175 14059
rect 16117 14019 16175 14025
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17218 14056 17224 14068
rect 17000 14028 17224 14056
rect 17000 14016 17006 14028
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 18506 14016 18512 14068
rect 18564 14056 18570 14068
rect 18601 14059 18659 14065
rect 18601 14056 18613 14059
rect 18564 14028 18613 14056
rect 18564 14016 18570 14028
rect 18601 14025 18613 14028
rect 18647 14025 18659 14059
rect 18601 14019 18659 14025
rect 13740 13988 13768 14016
rect 12176 13960 13400 13988
rect 13740 13960 14412 13988
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 9999 13892 11345 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 11333 13889 11345 13892
rect 11379 13920 11391 13923
rect 12158 13920 12164 13932
rect 11379 13892 12164 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 13372 13929 13400 13960
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13722 13920 13728 13932
rect 13403 13892 13728 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 14384 13929 14412 13960
rect 15396 13960 16804 13988
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 11020 13824 11253 13852
rect 11020 13812 11026 13824
rect 11241 13821 11253 13824
rect 11287 13852 11299 13855
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11287 13824 11805 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 13262 13852 13268 13864
rect 12759 13824 13268 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15396 13852 15424 13960
rect 16482 13880 16488 13932
rect 16540 13920 16546 13932
rect 16776 13929 16804 13960
rect 16577 13923 16635 13929
rect 16577 13920 16589 13923
rect 16540 13892 16589 13920
rect 16540 13880 16546 13892
rect 16577 13889 16589 13892
rect 16623 13889 16635 13923
rect 16577 13883 16635 13889
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 16807 13892 17785 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 17773 13889 17785 13892
rect 17819 13889 17831 13923
rect 18616 13920 18644 14019
rect 18690 14016 18696 14068
rect 18748 14056 18754 14068
rect 19978 14056 19984 14068
rect 18748 14028 19984 14056
rect 18748 14016 18754 14028
rect 19978 14016 19984 14028
rect 20036 14056 20042 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 20036 14028 20177 14056
rect 20036 14016 20042 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 20165 14019 20223 14025
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 22002 14056 22008 14068
rect 21963 14028 22008 14056
rect 22002 14016 22008 14028
rect 22060 14016 22066 14068
rect 24762 14016 24768 14068
rect 24820 14056 24826 14068
rect 25501 14059 25559 14065
rect 25501 14056 25513 14059
rect 24820 14028 25513 14056
rect 24820 14016 24826 14028
rect 25501 14025 25513 14028
rect 25547 14025 25559 14059
rect 26050 14056 26056 14068
rect 26011 14028 26056 14056
rect 25501 14019 25559 14025
rect 26050 14016 26056 14028
rect 26108 14016 26114 14068
rect 18616 13892 18920 13920
rect 17773 13883 17831 13889
rect 15470 13852 15476 13864
rect 15252 13824 15476 13852
rect 15252 13812 15258 13824
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15746 13812 15752 13864
rect 15804 13812 15810 13864
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 16592 13824 17417 13852
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10597 13787 10655 13793
rect 10597 13784 10609 13787
rect 9824 13756 10609 13784
rect 9824 13744 9830 13756
rect 10597 13753 10609 13756
rect 10643 13784 10655 13787
rect 11149 13787 11207 13793
rect 11149 13784 11161 13787
rect 10643 13756 11161 13784
rect 10643 13753 10655 13756
rect 10597 13747 10655 13753
rect 11149 13753 11161 13756
rect 11195 13753 11207 13787
rect 11149 13747 11207 13753
rect 13909 13787 13967 13793
rect 13909 13753 13921 13787
rect 13955 13784 13967 13787
rect 14274 13784 14280 13796
rect 13955 13756 14280 13784
rect 13955 13753 13967 13756
rect 13909 13747 13967 13753
rect 14274 13744 14280 13756
rect 14332 13784 14338 13796
rect 14636 13787 14694 13793
rect 14636 13784 14648 13787
rect 14332 13756 14648 13784
rect 14332 13744 14338 13756
rect 14636 13753 14648 13756
rect 14682 13784 14694 13787
rect 14734 13784 14740 13796
rect 14682 13756 14740 13784
rect 14682 13753 14694 13756
rect 14636 13747 14694 13753
rect 14734 13744 14740 13756
rect 14792 13744 14798 13796
rect 14918 13744 14924 13796
rect 14976 13784 14982 13796
rect 15378 13784 15384 13796
rect 14976 13756 15384 13784
rect 14976 13744 14982 13756
rect 15378 13744 15384 13756
rect 15436 13744 15442 13796
rect 10778 13716 10784 13728
rect 10739 13688 10784 13716
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 15764 13725 15792 13812
rect 16592 13784 16620 13824
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 18414 13812 18420 13864
rect 18472 13852 18478 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 18472 13824 18797 13852
rect 18472 13812 18478 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18892 13852 18920 13892
rect 20806 13880 20812 13932
rect 20864 13920 20870 13932
rect 21818 13920 21824 13932
rect 20864 13892 21824 13920
rect 20864 13880 20870 13892
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 22830 13920 22836 13932
rect 22695 13892 22836 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 22830 13880 22836 13892
rect 22888 13920 22894 13932
rect 24029 13923 24087 13929
rect 22888 13892 23152 13920
rect 22888 13880 22894 13892
rect 19041 13855 19099 13861
rect 19041 13852 19053 13855
rect 18892 13824 19053 13852
rect 18785 13815 18843 13821
rect 19041 13821 19053 13824
rect 19087 13821 19099 13855
rect 19041 13815 19099 13821
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 20438 13852 20444 13864
rect 19392 13824 20444 13852
rect 19392 13812 19398 13824
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 20898 13852 20904 13864
rect 20859 13824 20904 13852
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 22738 13852 22744 13864
rect 21324 13824 22744 13852
rect 21324 13812 21330 13824
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 23124 13861 23152 13892
rect 24029 13889 24041 13923
rect 24075 13920 24087 13923
rect 24075 13892 24256 13920
rect 24075 13889 24087 13892
rect 24029 13883 24087 13889
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 23477 13855 23535 13861
rect 23155 13824 23428 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 16500 13756 16620 13784
rect 16500 13728 16528 13756
rect 16666 13744 16672 13796
rect 16724 13784 16730 13796
rect 16945 13787 17003 13793
rect 16945 13784 16957 13787
rect 16724 13756 16957 13784
rect 16724 13744 16730 13756
rect 16945 13753 16957 13756
rect 16991 13753 17003 13787
rect 16945 13747 17003 13753
rect 21818 13744 21824 13796
rect 21876 13784 21882 13796
rect 22465 13787 22523 13793
rect 22465 13784 22477 13787
rect 21876 13756 22477 13784
rect 21876 13744 21882 13756
rect 22465 13753 22477 13756
rect 22511 13753 22523 13787
rect 23400 13784 23428 13824
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 23934 13852 23940 13864
rect 23523 13824 23940 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 23934 13812 23940 13824
rect 23992 13852 23998 13864
rect 24121 13855 24179 13861
rect 24121 13852 24133 13855
rect 23992 13824 24133 13852
rect 23992 13812 23998 13824
rect 24121 13821 24133 13824
rect 24167 13821 24179 13855
rect 24228 13852 24256 13892
rect 24377 13855 24435 13861
rect 24377 13852 24389 13855
rect 24228 13824 24389 13852
rect 24121 13815 24179 13821
rect 24377 13821 24389 13824
rect 24423 13852 24435 13855
rect 24854 13852 24860 13864
rect 24423 13824 24860 13852
rect 24423 13821 24435 13824
rect 24377 13815 24435 13821
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 24762 13784 24768 13796
rect 23400 13756 24768 13784
rect 22465 13747 22523 13753
rect 24762 13744 24768 13756
rect 24820 13744 24826 13796
rect 13173 13719 13231 13725
rect 13173 13716 13185 13719
rect 12952 13688 13185 13716
rect 12952 13676 12958 13688
rect 13173 13685 13185 13688
rect 13219 13685 13231 13719
rect 13173 13679 13231 13685
rect 15749 13719 15807 13725
rect 15749 13685 15761 13719
rect 15795 13685 15807 13719
rect 16482 13716 16488 13728
rect 16443 13688 16488 13716
rect 15749 13679 15807 13685
rect 16482 13676 16488 13688
rect 16540 13676 16546 13728
rect 18325 13719 18383 13725
rect 18325 13685 18337 13719
rect 18371 13716 18383 13719
rect 18506 13716 18512 13728
rect 18371 13688 18512 13716
rect 18371 13685 18383 13688
rect 18325 13679 18383 13685
rect 18506 13676 18512 13688
rect 18564 13676 18570 13728
rect 21266 13676 21272 13728
rect 21324 13716 21330 13728
rect 21634 13716 21640 13728
rect 21324 13688 21640 13716
rect 21324 13676 21330 13688
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 22370 13716 22376 13728
rect 22331 13688 22376 13716
rect 22370 13676 22376 13688
rect 22428 13676 22434 13728
rect 25130 13676 25136 13728
rect 25188 13716 25194 13728
rect 26050 13716 26056 13728
rect 25188 13688 26056 13716
rect 25188 13676 25194 13688
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 9766 13512 9772 13524
rect 9727 13484 9772 13512
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10321 13515 10379 13521
rect 10321 13512 10333 13515
rect 10008 13484 10333 13512
rect 10008 13472 10014 13484
rect 10321 13481 10333 13484
rect 10367 13512 10379 13515
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10367 13484 10701 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 10689 13481 10701 13484
rect 10735 13512 10747 13515
rect 10870 13512 10876 13524
rect 10735 13484 10876 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 10796 13385 10824 13484
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 13630 13512 13636 13524
rect 13591 13484 13636 13512
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14737 13515 14795 13521
rect 14737 13481 14749 13515
rect 14783 13512 14795 13515
rect 14826 13512 14832 13524
rect 14783 13484 14832 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 15102 13512 15108 13524
rect 15063 13484 15108 13512
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 17865 13515 17923 13521
rect 17865 13481 17877 13515
rect 17911 13512 17923 13515
rect 19518 13512 19524 13524
rect 17911 13484 19524 13512
rect 17911 13481 17923 13484
rect 17865 13475 17923 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 20254 13512 20260 13524
rect 20215 13484 20260 13512
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 20901 13515 20959 13521
rect 20901 13481 20913 13515
rect 20947 13512 20959 13515
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 20947 13484 22845 13512
rect 20947 13481 20959 13484
rect 20901 13475 20959 13481
rect 22833 13481 22845 13484
rect 22879 13512 22891 13515
rect 23477 13515 23535 13521
rect 23477 13512 23489 13515
rect 22879 13484 23489 13512
rect 22879 13481 22891 13484
rect 22833 13475 22891 13481
rect 23477 13481 23489 13484
rect 23523 13481 23535 13515
rect 23477 13475 23535 13481
rect 24029 13515 24087 13521
rect 24029 13481 24041 13515
rect 24075 13512 24087 13515
rect 24302 13512 24308 13524
rect 24075 13484 24308 13512
rect 24075 13481 24087 13484
rect 24029 13475 24087 13481
rect 24302 13472 24308 13484
rect 24360 13472 24366 13524
rect 25038 13512 25044 13524
rect 24999 13484 25044 13512
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 11048 13447 11106 13453
rect 11048 13413 11060 13447
rect 11094 13444 11106 13447
rect 11330 13444 11336 13456
rect 11094 13416 11336 13444
rect 11094 13413 11106 13416
rect 11048 13407 11106 13413
rect 11330 13404 11336 13416
rect 11388 13444 11394 13456
rect 12066 13444 12072 13456
rect 11388 13416 12072 13444
rect 11388 13404 11394 13416
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 16025 13447 16083 13453
rect 16025 13413 16037 13447
rect 16071 13444 16083 13447
rect 16114 13444 16120 13456
rect 16071 13416 16120 13444
rect 16071 13413 16083 13416
rect 16025 13407 16083 13413
rect 16114 13404 16120 13416
rect 16172 13404 16178 13456
rect 18230 13444 18236 13456
rect 18143 13416 18236 13444
rect 18230 13404 18236 13416
rect 18288 13444 18294 13456
rect 19242 13444 19248 13456
rect 18288 13416 19248 13444
rect 18288 13404 18294 13416
rect 19242 13404 19248 13416
rect 19300 13404 19306 13456
rect 20717 13447 20775 13453
rect 20717 13413 20729 13447
rect 20763 13444 20775 13447
rect 21450 13444 21456 13456
rect 20763 13416 21456 13444
rect 20763 13413 20775 13416
rect 20717 13407 20775 13413
rect 21450 13404 21456 13416
rect 21508 13404 21514 13456
rect 22925 13447 22983 13453
rect 22925 13413 22937 13447
rect 22971 13444 22983 13447
rect 23290 13444 23296 13456
rect 22971 13416 23296 13444
rect 22971 13413 22983 13416
rect 22925 13407 22983 13413
rect 23290 13404 23296 13416
rect 23348 13404 23354 13456
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13345 10839 13379
rect 12894 13376 12900 13388
rect 12855 13348 12900 13376
rect 10781 13339 10839 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13998 13376 14004 13388
rect 13959 13348 14004 13376
rect 13998 13336 14004 13348
rect 14056 13376 14062 13388
rect 15378 13376 15384 13388
rect 14056 13348 15384 13376
rect 14056 13336 14062 13348
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 18325 13379 18383 13385
rect 18325 13345 18337 13379
rect 18371 13376 18383 13379
rect 19150 13376 19156 13388
rect 18371 13348 19156 13376
rect 18371 13345 18383 13348
rect 18325 13339 18383 13345
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19610 13376 19616 13388
rect 19571 13348 19616 13376
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 21269 13379 21327 13385
rect 21269 13345 21281 13379
rect 21315 13376 21327 13379
rect 21818 13376 21824 13388
rect 21315 13348 21824 13376
rect 21315 13345 21327 13348
rect 21269 13339 21327 13345
rect 21818 13336 21824 13348
rect 21876 13336 21882 13388
rect 24026 13336 24032 13388
rect 24084 13376 24090 13388
rect 24397 13379 24455 13385
rect 24397 13376 24409 13379
rect 24084 13348 24409 13376
rect 24084 13336 24090 13348
rect 24397 13345 24409 13348
rect 24443 13345 24455 13379
rect 24397 13339 24455 13345
rect 24489 13379 24547 13385
rect 24489 13345 24501 13379
rect 24535 13376 24547 13379
rect 24670 13376 24676 13388
rect 24535 13348 24676 13376
rect 24535 13345 24547 13348
rect 24489 13339 24547 13345
rect 24670 13336 24676 13348
rect 24728 13376 24734 13388
rect 25409 13379 25467 13385
rect 25409 13376 25421 13379
rect 24728 13348 25421 13376
rect 24728 13336 24734 13348
rect 25409 13345 25421 13348
rect 25455 13345 25467 13379
rect 25409 13339 25467 13345
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 14090 13308 14096 13320
rect 13587 13280 14096 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14274 13268 14280 13320
rect 14332 13308 14338 13320
rect 15102 13308 15108 13320
rect 14332 13280 15108 13308
rect 14332 13268 14338 13280
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 18506 13308 18512 13320
rect 18419 13280 18512 13308
rect 18506 13268 18512 13280
rect 18564 13308 18570 13320
rect 18874 13308 18880 13320
rect 18564 13280 18880 13308
rect 18564 13268 18570 13280
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 19518 13268 19524 13320
rect 19576 13308 19582 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19576 13280 19717 13308
rect 19576 13268 19582 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19886 13308 19892 13320
rect 19847 13280 19892 13308
rect 19705 13271 19763 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 21082 13268 21088 13320
rect 21140 13308 21146 13320
rect 21361 13311 21419 13317
rect 21361 13308 21373 13311
rect 21140 13280 21373 13308
rect 21140 13268 21146 13280
rect 21361 13277 21373 13280
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 23106 13308 23112 13320
rect 21591 13280 22968 13308
rect 23067 13280 23112 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 15286 13200 15292 13252
rect 15344 13240 15350 13252
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 15344 13212 15577 13240
rect 15344 13200 15350 13212
rect 15565 13209 15577 13212
rect 15611 13240 15623 13243
rect 15930 13240 15936 13252
rect 15611 13212 15936 13240
rect 15611 13209 15623 13212
rect 15565 13203 15623 13209
rect 15930 13200 15936 13212
rect 15988 13200 15994 13252
rect 17310 13240 17316 13252
rect 17271 13212 17316 13240
rect 17310 13200 17316 13212
rect 17368 13240 17374 13252
rect 17586 13240 17592 13252
rect 17368 13212 17592 13240
rect 17368 13200 17374 13212
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 20530 13200 20536 13252
rect 20588 13240 20594 13252
rect 21560 13240 21588 13271
rect 20588 13212 21588 13240
rect 22097 13243 22155 13249
rect 20588 13200 20594 13212
rect 22097 13209 22109 13243
rect 22143 13240 22155 13243
rect 22370 13240 22376 13252
rect 22143 13212 22376 13240
rect 22143 13209 22155 13212
rect 22097 13203 22155 13209
rect 22370 13200 22376 13212
rect 22428 13200 22434 13252
rect 22940 13240 22968 13280
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13308 23995 13311
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 23983 13280 24593 13308
rect 23983 13277 23995 13280
rect 23937 13271 23995 13277
rect 24581 13277 24593 13280
rect 24627 13308 24639 13311
rect 24762 13308 24768 13320
rect 24627 13280 24768 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 23750 13240 23756 13252
rect 22940 13212 23756 13240
rect 23750 13200 23756 13212
rect 23808 13200 23814 13252
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 16390 13172 16396 13184
rect 11204 13144 16396 13172
rect 11204 13132 11210 13144
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 18877 13175 18935 13181
rect 18877 13172 18889 13175
rect 18012 13144 18889 13172
rect 18012 13132 18018 13144
rect 18877 13141 18889 13144
rect 18923 13141 18935 13175
rect 19242 13172 19248 13184
rect 19203 13144 19248 13172
rect 18877 13135 18935 13141
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 22462 13172 22468 13184
rect 22423 13144 22468 13172
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 9950 12968 9956 12980
rect 9911 12940 9956 12968
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 10962 12968 10968 12980
rect 10827 12940 10968 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 12250 12968 12256 12980
rect 12211 12940 12256 12968
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 14148 12940 16221 12968
rect 14148 12928 14154 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 16209 12931 16267 12937
rect 18233 12971 18291 12977
rect 18233 12937 18245 12971
rect 18279 12968 18291 12971
rect 19610 12968 19616 12980
rect 18279 12940 19616 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 19978 12968 19984 12980
rect 19751 12940 19984 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 21082 12928 21088 12980
rect 21140 12968 21146 12980
rect 21729 12971 21787 12977
rect 21729 12968 21741 12971
rect 21140 12940 21741 12968
rect 21140 12928 21146 12940
rect 21729 12937 21741 12940
rect 21775 12937 21787 12971
rect 21729 12931 21787 12937
rect 24854 12928 24860 12980
rect 24912 12968 24918 12980
rect 25130 12968 25136 12980
rect 24912 12940 25136 12968
rect 24912 12928 24918 12940
rect 25130 12928 25136 12940
rect 25188 12968 25194 12980
rect 25501 12971 25559 12977
rect 25501 12968 25513 12971
rect 25188 12940 25513 12968
rect 25188 12928 25194 12940
rect 25501 12937 25513 12940
rect 25547 12937 25559 12971
rect 25501 12931 25559 12937
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 15105 12903 15163 12909
rect 15105 12900 15117 12903
rect 14792 12872 15117 12900
rect 14792 12860 14798 12872
rect 15105 12869 15117 12872
rect 15151 12869 15163 12903
rect 15105 12863 15163 12869
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12900 15807 12903
rect 16114 12900 16120 12912
rect 15795 12872 16120 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 16114 12860 16120 12872
rect 16172 12860 16178 12912
rect 24026 12900 24032 12912
rect 23987 12872 24032 12900
rect 24026 12860 24032 12872
rect 24084 12860 24090 12912
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 11330 12832 11336 12844
rect 10367 12804 11336 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 16758 12832 16764 12844
rect 13679 12804 13860 12832
rect 16719 12804 16764 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 13832 12776 13860 12804
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 18874 12832 18880 12844
rect 17543 12804 18880 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 22557 12835 22615 12841
rect 22557 12832 22569 12835
rect 22244 12804 22569 12832
rect 22244 12792 22250 12804
rect 22557 12801 22569 12804
rect 22603 12801 22615 12835
rect 24118 12832 24124 12844
rect 24079 12804 24124 12832
rect 22557 12795 22615 12801
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 11974 12764 11980 12776
rect 11287 12736 11980 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 12492 12736 13185 12764
rect 12492 12724 12498 12736
rect 13173 12733 13185 12736
rect 13219 12733 13231 12767
rect 13722 12764 13728 12776
rect 13683 12736 13728 12764
rect 13173 12727 13231 12733
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 13992 12767 14050 12773
rect 13992 12764 14004 12767
rect 13872 12736 14004 12764
rect 13872 12724 13878 12736
rect 13992 12733 14004 12736
rect 14038 12764 14050 12767
rect 14274 12764 14280 12776
rect 14038 12736 14280 12764
rect 14038 12733 14050 12736
rect 13992 12727 14050 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 17862 12764 17868 12776
rect 17775 12736 17868 12764
rect 17862 12724 17868 12736
rect 17920 12764 17926 12776
rect 18690 12764 18696 12776
rect 17920 12736 18696 12764
rect 17920 12724 17926 12736
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 19058 12724 19064 12776
rect 19116 12764 19122 12776
rect 19797 12767 19855 12773
rect 19797 12764 19809 12767
rect 19116 12736 19809 12764
rect 19116 12724 19122 12736
rect 19797 12733 19809 12736
rect 19843 12764 19855 12767
rect 20898 12764 20904 12776
rect 19843 12736 20904 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 22278 12764 22284 12776
rect 22191 12736 22284 12764
rect 22278 12724 22284 12736
rect 22336 12764 22342 12776
rect 22462 12764 22468 12776
rect 22336 12736 22468 12764
rect 22336 12724 22342 12736
rect 22462 12724 22468 12736
rect 22520 12724 22526 12776
rect 10689 12699 10747 12705
rect 10689 12665 10701 12699
rect 10735 12696 10747 12699
rect 11149 12699 11207 12705
rect 11149 12696 11161 12699
rect 10735 12668 11161 12696
rect 10735 12665 10747 12668
rect 10689 12659 10747 12665
rect 11149 12665 11161 12668
rect 11195 12696 11207 12699
rect 12066 12696 12072 12708
rect 11195 12668 12072 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 12713 12699 12771 12705
rect 12713 12665 12725 12699
rect 12759 12696 12771 12699
rect 13630 12696 13636 12708
rect 12759 12668 13636 12696
rect 12759 12665 12771 12668
rect 12713 12659 12771 12665
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 16482 12656 16488 12708
rect 16540 12696 16546 12708
rect 16669 12699 16727 12705
rect 16669 12696 16681 12699
rect 16540 12668 16681 12696
rect 16540 12656 16546 12668
rect 16669 12665 16681 12668
rect 16715 12665 16727 12699
rect 16669 12659 16727 12665
rect 18322 12656 18328 12708
rect 18380 12696 18386 12708
rect 19337 12699 19395 12705
rect 18380 12668 18828 12696
rect 18380 12656 18386 12668
rect 18800 12640 18828 12668
rect 19337 12665 19349 12699
rect 19383 12696 19395 12699
rect 19886 12696 19892 12708
rect 19383 12668 19892 12696
rect 19383 12665 19395 12668
rect 19337 12659 19395 12665
rect 19886 12656 19892 12668
rect 19944 12656 19950 12708
rect 19978 12656 19984 12708
rect 20036 12705 20042 12708
rect 20036 12699 20100 12705
rect 20036 12665 20054 12699
rect 20088 12696 20100 12699
rect 20254 12696 20260 12708
rect 20088 12668 20260 12696
rect 20088 12665 20100 12668
rect 20036 12659 20100 12665
rect 20036 12656 20042 12659
rect 20254 12656 20260 12668
rect 20312 12656 20318 12708
rect 23106 12696 23112 12708
rect 23019 12668 23112 12696
rect 23106 12656 23112 12668
rect 23164 12696 23170 12708
rect 23477 12699 23535 12705
rect 23477 12696 23489 12699
rect 23164 12668 23489 12696
rect 23164 12656 23170 12668
rect 23477 12665 23489 12668
rect 23523 12696 23535 12699
rect 24388 12699 24446 12705
rect 24388 12696 24400 12699
rect 23523 12668 24400 12696
rect 23523 12665 23535 12668
rect 23477 12659 23535 12665
rect 24388 12665 24400 12668
rect 24434 12696 24446 12699
rect 24946 12696 24952 12708
rect 24434 12668 24952 12696
rect 24434 12665 24446 12668
rect 24388 12659 24446 12665
rect 24946 12656 24952 12668
rect 25004 12656 25010 12708
rect 11882 12628 11888 12640
rect 11843 12600 11888 12628
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 16114 12628 16120 12640
rect 16075 12600 16120 12628
rect 16114 12588 16120 12600
rect 16172 12628 16178 12640
rect 16577 12631 16635 12637
rect 16577 12628 16589 12631
rect 16172 12600 16589 12628
rect 16172 12588 16178 12600
rect 16577 12597 16589 12600
rect 16623 12597 16635 12631
rect 16577 12591 16635 12597
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 18601 12631 18659 12637
rect 18601 12628 18613 12631
rect 18564 12600 18613 12628
rect 18564 12588 18570 12600
rect 18601 12597 18613 12600
rect 18647 12597 18659 12631
rect 18601 12591 18659 12597
rect 18782 12588 18788 12640
rect 18840 12588 18846 12640
rect 19904 12628 19932 12656
rect 20530 12628 20536 12640
rect 19904 12600 20536 12628
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 21082 12588 21088 12640
rect 21140 12628 21146 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 21140 12600 21189 12628
rect 21140 12588 21146 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 21177 12591 21235 12597
rect 21818 12588 21824 12640
rect 21876 12628 21882 12640
rect 22189 12631 22247 12637
rect 22189 12628 22201 12631
rect 21876 12600 22201 12628
rect 21876 12588 21882 12600
rect 22189 12597 22201 12600
rect 22235 12628 22247 12631
rect 22922 12628 22928 12640
rect 22235 12600 22928 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11330 12424 11336 12436
rect 11287 12396 11336 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 11974 12424 11980 12436
rect 11532 12396 11980 12424
rect 10873 12359 10931 12365
rect 10873 12325 10885 12359
rect 10919 12356 10931 12359
rect 11532 12356 11560 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 13814 12424 13820 12436
rect 13775 12396 13820 12424
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 14185 12427 14243 12433
rect 14185 12393 14197 12427
rect 14231 12424 14243 12427
rect 15194 12424 15200 12436
rect 14231 12396 15200 12424
rect 14231 12393 14243 12396
rect 14185 12387 14243 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15378 12424 15384 12436
rect 15335 12396 15384 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 15988 12396 16313 12424
rect 15988 12384 15994 12396
rect 16301 12393 16313 12396
rect 16347 12424 16359 12427
rect 16482 12424 16488 12436
rect 16347 12396 16488 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 16758 12424 16764 12436
rect 16719 12396 16764 12424
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 18414 12384 18420 12436
rect 18472 12424 18478 12436
rect 19058 12424 19064 12436
rect 18472 12396 19064 12424
rect 18472 12384 18478 12396
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 20165 12427 20223 12433
rect 20165 12424 20177 12427
rect 19392 12396 20177 12424
rect 19392 12384 19398 12396
rect 20165 12393 20177 12396
rect 20211 12393 20223 12427
rect 20622 12424 20628 12436
rect 20583 12396 20628 12424
rect 20165 12387 20223 12393
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 22830 12424 22836 12436
rect 22791 12396 22836 12424
rect 22830 12384 22836 12396
rect 22888 12384 22894 12436
rect 23290 12424 23296 12436
rect 23251 12396 23296 12424
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 23750 12384 23756 12436
rect 23808 12424 23814 12436
rect 24946 12424 24952 12436
rect 23808 12396 23888 12424
rect 24907 12396 24952 12424
rect 23808 12384 23814 12396
rect 10919 12328 11560 12356
rect 10919 12325 10931 12328
rect 10873 12319 10931 12325
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 11784 12359 11842 12365
rect 11784 12356 11796 12359
rect 11664 12328 11796 12356
rect 11664 12316 11670 12328
rect 11784 12325 11796 12328
rect 11830 12356 11842 12359
rect 12158 12356 12164 12368
rect 11830 12328 12164 12356
rect 11830 12325 11842 12328
rect 11784 12319 11842 12325
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 15657 12359 15715 12365
rect 15657 12325 15669 12359
rect 15703 12356 15715 12359
rect 16206 12356 16212 12368
rect 15703 12328 16212 12356
rect 15703 12325 15715 12328
rect 15657 12319 15715 12325
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 15838 12288 15844 12300
rect 15795 12260 15844 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12189 11575 12223
rect 15102 12220 15108 12232
rect 15063 12192 15108 12220
rect 11517 12183 11575 12189
rect 11532 12084 11560 12183
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 15930 12220 15936 12232
rect 15843 12192 15936 12220
rect 15930 12180 15936 12192
rect 15988 12220 15994 12232
rect 16776 12220 16804 12384
rect 17589 12359 17647 12365
rect 17589 12325 17601 12359
rect 17635 12356 17647 12359
rect 17770 12356 17776 12368
rect 17635 12328 17776 12356
rect 17635 12325 17647 12328
rect 17589 12319 17647 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 18325 12359 18383 12365
rect 18325 12325 18337 12359
rect 18371 12356 18383 12359
rect 18506 12356 18512 12368
rect 18371 12328 18512 12356
rect 18371 12325 18383 12328
rect 18325 12319 18383 12325
rect 18506 12316 18512 12328
rect 18564 12356 18570 12368
rect 19426 12356 19432 12368
rect 18564 12328 19432 12356
rect 18564 12316 18570 12328
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 21082 12316 21088 12368
rect 21140 12365 21146 12368
rect 23860 12365 23888 12396
rect 24946 12384 24952 12396
rect 25004 12384 25010 12436
rect 21140 12359 21204 12365
rect 21140 12325 21158 12359
rect 21192 12325 21204 12359
rect 21140 12319 21204 12325
rect 23836 12359 23894 12365
rect 23836 12325 23848 12359
rect 23882 12325 23894 12359
rect 23836 12319 23894 12325
rect 21140 12316 21146 12319
rect 24118 12316 24124 12368
rect 24176 12356 24182 12368
rect 25314 12356 25320 12368
rect 24176 12328 25320 12356
rect 24176 12316 24182 12328
rect 25314 12316 25320 12328
rect 25372 12356 25378 12368
rect 25501 12359 25559 12365
rect 25501 12356 25513 12359
rect 25372 12328 25513 12356
rect 25372 12316 25378 12328
rect 25501 12325 25513 12328
rect 25547 12325 25559 12359
rect 25501 12319 25559 12325
rect 18874 12288 18880 12300
rect 18524 12260 18880 12288
rect 18524 12232 18552 12260
rect 18874 12248 18880 12260
rect 18932 12288 18938 12300
rect 19153 12291 19211 12297
rect 19153 12288 19165 12291
rect 18932 12260 19165 12288
rect 18932 12248 18938 12260
rect 19153 12257 19165 12260
rect 19199 12257 19211 12291
rect 19153 12251 19211 12257
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 20898 12288 20904 12300
rect 20772 12260 20904 12288
rect 20772 12248 20778 12260
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 22830 12248 22836 12300
rect 22888 12288 22894 12300
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 22888 12260 23581 12288
rect 22888 12248 22894 12260
rect 23569 12257 23581 12260
rect 23615 12288 23627 12291
rect 24136 12288 24164 12316
rect 23615 12260 24164 12288
rect 23615 12257 23627 12260
rect 23569 12251 23627 12257
rect 15988 12192 16804 12220
rect 15988 12180 15994 12192
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 17678 12220 17684 12232
rect 17552 12192 17684 12220
rect 17552 12180 17558 12192
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 16758 12112 16764 12164
rect 16816 12152 16822 12164
rect 17221 12155 17279 12161
rect 17221 12152 17233 12155
rect 16816 12124 17233 12152
rect 16816 12112 16822 12124
rect 17221 12121 17233 12124
rect 17267 12121 17279 12155
rect 17788 12152 17816 12183
rect 18506 12180 18512 12232
rect 18564 12180 18570 12232
rect 19058 12180 19064 12232
rect 19116 12220 19122 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19116 12192 19257 12220
rect 19116 12180 19122 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 19352 12152 19380 12183
rect 17221 12115 17279 12121
rect 17328 12124 17816 12152
rect 18708 12124 19380 12152
rect 17328 12096 17356 12124
rect 18708 12096 18736 12124
rect 11882 12084 11888 12096
rect 11532 12056 11888 12084
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 12897 12087 12955 12093
rect 12897 12053 12909 12087
rect 12943 12084 12955 12087
rect 12986 12084 12992 12096
rect 12943 12056 12992 12084
rect 12943 12053 12955 12056
rect 12897 12047 12955 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 13872 12056 14657 12084
rect 13872 12044 13878 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 17129 12087 17187 12093
rect 17129 12053 17141 12087
rect 17175 12084 17187 12087
rect 17310 12084 17316 12096
rect 17175 12056 17316 12084
rect 17175 12053 17187 12056
rect 17129 12047 17187 12053
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 18690 12084 18696 12096
rect 18651 12056 18696 12084
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 18874 12084 18880 12096
rect 18831 12056 18880 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 19889 12087 19947 12093
rect 19889 12084 19901 12087
rect 19208 12056 19901 12084
rect 19208 12044 19214 12056
rect 19889 12053 19901 12056
rect 19935 12084 19947 12087
rect 20898 12084 20904 12096
rect 19935 12056 20904 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 22244 12056 22293 12084
rect 22244 12044 22250 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22281 12047 22339 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 11606 11880 11612 11892
rect 11567 11852 11612 11880
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 15197 11883 15255 11889
rect 15197 11849 15209 11883
rect 15243 11880 15255 11883
rect 15470 11880 15476 11892
rect 15243 11852 15476 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 16206 11880 16212 11892
rect 16167 11852 16212 11880
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17497 11883 17555 11889
rect 17497 11849 17509 11883
rect 17543 11880 17555 11883
rect 17678 11880 17684 11892
rect 17543 11852 17684 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 18414 11880 18420 11892
rect 18064 11852 18420 11880
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11744 12771 11747
rect 13354 11744 13360 11756
rect 12759 11716 13360 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 16942 11744 16948 11756
rect 16903 11716 16948 11744
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 13173 11679 13231 11685
rect 13173 11676 13185 11679
rect 12492 11648 13185 11676
rect 12492 11636 12498 11648
rect 13173 11645 13185 11648
rect 13219 11645 13231 11679
rect 13814 11676 13820 11688
rect 13775 11648 13820 11676
rect 13173 11639 13231 11645
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 16758 11676 16764 11688
rect 16719 11648 16764 11676
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18064 11685 18092 11852
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 20625 11883 20683 11889
rect 20625 11849 20637 11883
rect 20671 11880 20683 11883
rect 21082 11880 21088 11892
rect 20671 11852 21088 11880
rect 20671 11849 20683 11852
rect 20625 11843 20683 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 23109 11883 23167 11889
rect 23109 11849 23121 11883
rect 23155 11880 23167 11883
rect 23750 11880 23756 11892
rect 23155 11852 23756 11880
rect 23155 11849 23167 11852
rect 23109 11843 23167 11849
rect 23750 11840 23756 11852
rect 23808 11840 23814 11892
rect 25314 11880 25320 11892
rect 25275 11852 25320 11880
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 20530 11772 20536 11824
rect 20588 11812 20594 11824
rect 20809 11815 20867 11821
rect 20809 11812 20821 11815
rect 20588 11784 20821 11812
rect 20588 11772 20594 11784
rect 20809 11781 20821 11784
rect 20855 11812 20867 11815
rect 20901 11815 20959 11821
rect 20901 11812 20913 11815
rect 20855 11784 20913 11812
rect 20855 11781 20867 11784
rect 20809 11775 20867 11781
rect 20901 11781 20913 11784
rect 20947 11781 20959 11815
rect 20901 11775 20959 11781
rect 22465 11815 22523 11821
rect 22465 11781 22477 11815
rect 22511 11812 22523 11815
rect 23014 11812 23020 11824
rect 22511 11784 23020 11812
rect 22511 11781 22523 11784
rect 22465 11775 22523 11781
rect 23014 11772 23020 11784
rect 23072 11772 23078 11824
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 20772 11716 21097 11744
rect 20772 11704 20778 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 24210 11744 24216 11756
rect 24171 11716 24216 11744
rect 21085 11707 21143 11713
rect 24210 11704 24216 11716
rect 24268 11744 24274 11756
rect 24578 11744 24584 11756
rect 24268 11716 24584 11744
rect 24268 11704 24274 11716
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 24946 11744 24952 11756
rect 24907 11716 24952 11744
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 18012 11648 18061 11676
rect 18012 11636 18018 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11676 20867 11679
rect 21341 11679 21399 11685
rect 21341 11676 21353 11679
rect 20855 11648 21353 11676
rect 20855 11645 20867 11648
rect 20809 11639 20867 11645
rect 21341 11645 21353 11648
rect 21387 11676 21399 11679
rect 22186 11676 22192 11688
rect 21387 11648 22192 11676
rect 21387 11645 21399 11648
rect 21341 11639 21399 11645
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 13722 11608 13728 11620
rect 13683 11580 13728 11608
rect 13722 11568 13728 11580
rect 13780 11608 13786 11620
rect 14062 11611 14120 11617
rect 14062 11608 14074 11611
rect 13780 11580 14074 11608
rect 13780 11568 13786 11580
rect 14062 11577 14074 11580
rect 14108 11577 14120 11611
rect 14062 11571 14120 11577
rect 18316 11611 18374 11617
rect 18316 11577 18328 11611
rect 18362 11608 18374 11611
rect 18690 11608 18696 11620
rect 18362 11580 18696 11608
rect 18362 11577 18374 11580
rect 18316 11571 18374 11577
rect 18690 11568 18696 11580
rect 18748 11608 18754 11620
rect 19981 11611 20039 11617
rect 19981 11608 19993 11611
rect 18748 11580 19993 11608
rect 18748 11568 18754 11580
rect 19981 11577 19993 11580
rect 20027 11577 20039 11611
rect 19981 11571 20039 11577
rect 23477 11611 23535 11617
rect 23477 11577 23489 11611
rect 23523 11608 23535 11611
rect 24673 11611 24731 11617
rect 24673 11608 24685 11611
rect 23523 11580 24685 11608
rect 23523 11577 23535 11580
rect 23477 11571 23535 11577
rect 24673 11577 24685 11580
rect 24719 11608 24731 11611
rect 24854 11608 24860 11620
rect 24719 11580 24860 11608
rect 24719 11577 24731 11580
rect 24673 11571 24731 11577
rect 24854 11568 24860 11580
rect 24912 11568 24918 11620
rect 11882 11540 11888 11552
rect 11843 11512 11888 11540
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 15838 11540 15844 11552
rect 15799 11512 15844 11540
rect 15838 11500 15844 11512
rect 15896 11500 15902 11552
rect 16298 11500 16304 11552
rect 16356 11540 16362 11552
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 16356 11512 16405 11540
rect 16356 11500 16362 11512
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 17770 11540 17776 11552
rect 16908 11512 16953 11540
rect 17731 11512 17776 11540
rect 16908 11500 16914 11512
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 19392 11512 19441 11540
rect 19392 11500 19398 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 21726 11500 21732 11552
rect 21784 11540 21790 11552
rect 23658 11540 23664 11552
rect 21784 11512 23664 11540
rect 21784 11500 21790 11512
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 24210 11500 24216 11552
rect 24268 11540 24274 11552
rect 24305 11543 24363 11549
rect 24305 11540 24317 11543
rect 24268 11512 24317 11540
rect 24268 11500 24274 11512
rect 24305 11509 24317 11512
rect 24351 11509 24363 11543
rect 24305 11503 24363 11509
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 24765 11543 24823 11549
rect 24765 11540 24777 11543
rect 24636 11512 24777 11540
rect 24636 11500 24642 11512
rect 24765 11509 24777 11512
rect 24811 11509 24823 11543
rect 24765 11503 24823 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 13817 11339 13875 11345
rect 13817 11336 13829 11339
rect 13780 11308 13829 11336
rect 13780 11296 13786 11308
rect 13817 11305 13829 11308
rect 13863 11336 13875 11339
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 13863 11308 14473 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 14461 11305 14473 11308
rect 14507 11336 14519 11339
rect 14826 11336 14832 11348
rect 14507 11308 14832 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 14826 11296 14832 11308
rect 14884 11336 14890 11348
rect 15105 11339 15163 11345
rect 15105 11336 15117 11339
rect 14884 11308 15117 11336
rect 14884 11296 14890 11308
rect 15105 11305 15117 11308
rect 15151 11336 15163 11339
rect 15930 11336 15936 11348
rect 15151 11308 15936 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 16942 11336 16948 11348
rect 16623 11308 16948 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 16942 11296 16948 11308
rect 17000 11336 17006 11348
rect 18230 11336 18236 11348
rect 17000 11308 18236 11336
rect 17000 11296 17006 11308
rect 18230 11296 18236 11308
rect 18288 11336 18294 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 18288 11308 18429 11336
rect 18288 11296 18294 11308
rect 18417 11305 18429 11308
rect 18463 11305 18475 11339
rect 18417 11299 18475 11305
rect 18785 11339 18843 11345
rect 18785 11305 18797 11339
rect 18831 11336 18843 11339
rect 19058 11336 19064 11348
rect 18831 11308 19064 11336
rect 18831 11305 18843 11308
rect 18785 11299 18843 11305
rect 19058 11296 19064 11308
rect 19116 11336 19122 11348
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 19116 11308 19349 11336
rect 19116 11296 19122 11308
rect 19337 11305 19349 11308
rect 19383 11305 19395 11339
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 19337 11299 19395 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20898 11336 20904 11348
rect 20859 11308 20904 11336
rect 20898 11296 20904 11308
rect 20956 11296 20962 11348
rect 21269 11339 21327 11345
rect 21269 11305 21281 11339
rect 21315 11336 21327 11339
rect 21450 11336 21456 11348
rect 21315 11308 21456 11336
rect 21315 11305 21327 11308
rect 21269 11299 21327 11305
rect 21450 11296 21456 11308
rect 21508 11336 21514 11348
rect 22002 11336 22008 11348
rect 21508 11308 22008 11336
rect 21508 11296 21514 11308
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11336 22799 11339
rect 22830 11336 22836 11348
rect 22787 11308 22836 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23750 11296 23756 11348
rect 23808 11336 23814 11348
rect 24213 11339 24271 11345
rect 24213 11336 24225 11339
rect 23808 11308 24225 11336
rect 23808 11296 23814 11308
rect 24213 11305 24225 11308
rect 24259 11305 24271 11339
rect 24213 11299 24271 11305
rect 24857 11339 24915 11345
rect 24857 11305 24869 11339
rect 24903 11336 24915 11339
rect 24946 11336 24952 11348
rect 24903 11308 24952 11336
rect 24903 11305 24915 11308
rect 24857 11299 24915 11305
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 25682 11336 25688 11348
rect 25547 11308 25688 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 25682 11296 25688 11308
rect 25740 11296 25746 11348
rect 12452 11240 13860 11268
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 12452 11209 12480 11240
rect 13832 11212 13860 11240
rect 15378 11228 15384 11280
rect 15436 11268 15442 11280
rect 16022 11268 16028 11280
rect 15436 11240 16028 11268
rect 15436 11228 15442 11240
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 19797 11271 19855 11277
rect 19797 11237 19809 11271
rect 19843 11268 19855 11271
rect 20162 11268 20168 11280
rect 19843 11240 20168 11268
rect 19843 11237 19855 11240
rect 19797 11231 19855 11237
rect 20162 11228 20168 11240
rect 20220 11228 20226 11280
rect 20272 11268 20300 11296
rect 20272 11240 21404 11268
rect 12710 11209 12716 11212
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 11940 11172 12449 11200
rect 11940 11160 11946 11172
rect 12437 11169 12449 11172
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 12704 11163 12716 11209
rect 12768 11200 12774 11212
rect 12768 11172 12804 11200
rect 12710 11160 12716 11163
rect 12768 11160 12774 11172
rect 13814 11160 13820 11212
rect 13872 11160 13878 11212
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 16482 11200 16488 11212
rect 15887 11172 16488 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 17310 11209 17316 11212
rect 17304 11200 17316 11209
rect 17271 11172 17316 11200
rect 17304 11163 17316 11172
rect 17310 11160 17316 11163
rect 17368 11160 17374 11212
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19392 11172 19533 11200
rect 19392 11160 19398 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 21376 11200 21404 11240
rect 21376 11172 21496 11200
rect 19521 11163 19579 11169
rect 15930 11132 15936 11144
rect 15891 11104 15936 11132
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 16022 11092 16028 11144
rect 16080 11132 16086 11144
rect 16080 11104 16125 11132
rect 16080 11092 16086 11104
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 17000 11104 17049 11132
rect 17000 11092 17006 11104
rect 17037 11101 17049 11104
rect 17083 11101 17095 11135
rect 21358 11132 21364 11144
rect 21319 11104 21364 11132
rect 17037 11095 17095 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 21468 11141 21496 11172
rect 22646 11160 22652 11212
rect 22704 11200 22710 11212
rect 22848 11209 22876 11296
rect 23014 11228 23020 11280
rect 23072 11277 23078 11280
rect 23072 11271 23136 11277
rect 23072 11237 23090 11271
rect 23124 11237 23136 11271
rect 23072 11231 23136 11237
rect 23072 11228 23078 11231
rect 22833 11203 22891 11209
rect 22833 11200 22845 11203
rect 22704 11172 22845 11200
rect 22704 11160 22710 11172
rect 22833 11169 22845 11172
rect 22879 11169 22891 11203
rect 25314 11200 25320 11212
rect 25275 11172 25320 11200
rect 22833 11163 22891 11169
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 21453 11135 21511 11141
rect 21453 11101 21465 11135
rect 21499 11101 21511 11135
rect 21453 11095 21511 11101
rect 10873 11067 10931 11073
rect 10873 11033 10885 11067
rect 10919 11064 10931 11067
rect 10962 11064 10968 11076
rect 10919 11036 10968 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 11698 11024 11704 11076
rect 11756 11064 11762 11076
rect 15473 11067 15531 11073
rect 11756 11036 12480 11064
rect 11756 11024 11762 11036
rect 11882 10996 11888 11008
rect 11843 10968 11888 10996
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 12342 10996 12348 11008
rect 12303 10968 12348 10996
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 12452 10996 12480 11036
rect 15473 11033 15485 11067
rect 15519 11064 15531 11067
rect 16850 11064 16856 11076
rect 15519 11036 16856 11064
rect 15519 11033 15531 11036
rect 15473 11027 15531 11033
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 18506 11024 18512 11076
rect 18564 11064 18570 11076
rect 19061 11067 19119 11073
rect 19061 11064 19073 11067
rect 18564 11036 19073 11064
rect 18564 11024 18570 11036
rect 19061 11033 19073 11036
rect 19107 11064 19119 11067
rect 21913 11067 21971 11073
rect 21913 11064 21925 11067
rect 19107 11036 19380 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 19352 11008 19380 11036
rect 20640 11036 21925 11064
rect 13998 10996 14004 11008
rect 12452 10968 14004 10996
rect 13998 10956 14004 10968
rect 14056 10996 14062 11008
rect 18785 10999 18843 11005
rect 18785 10996 18797 10999
rect 14056 10968 18797 10996
rect 14056 10956 14062 10968
rect 18785 10965 18797 10968
rect 18831 10965 18843 10999
rect 18785 10959 18843 10965
rect 19334 10956 19340 11008
rect 19392 10956 19398 11008
rect 19886 10956 19892 11008
rect 19944 10996 19950 11008
rect 20640 10996 20668 11036
rect 21913 11033 21925 11036
rect 21959 11033 21971 11067
rect 21913 11027 21971 11033
rect 19944 10968 20668 10996
rect 20717 10999 20775 11005
rect 19944 10956 19950 10968
rect 20717 10965 20729 10999
rect 20763 10996 20775 10999
rect 21634 10996 21640 11008
rect 20763 10968 21640 10996
rect 20763 10965 20775 10968
rect 20717 10959 20775 10965
rect 21634 10956 21640 10968
rect 21692 10956 21698 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 14182 10792 14188 10804
rect 14143 10764 14188 10792
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 17037 10795 17095 10801
rect 17037 10792 17049 10795
rect 16080 10764 17049 10792
rect 16080 10752 16086 10764
rect 17037 10761 17049 10764
rect 17083 10792 17095 10795
rect 17310 10792 17316 10804
rect 17083 10764 17316 10792
rect 17083 10761 17095 10764
rect 17037 10755 17095 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17678 10752 17684 10804
rect 17736 10792 17742 10804
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17736 10764 17785 10792
rect 17736 10752 17742 10764
rect 17773 10761 17785 10764
rect 17819 10792 17831 10795
rect 19150 10792 19156 10804
rect 17819 10764 19156 10792
rect 17819 10761 17831 10764
rect 17773 10755 17831 10761
rect 12437 10727 12495 10733
rect 12437 10724 12449 10727
rect 11808 10696 12449 10724
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10656 10747 10659
rect 11422 10656 11428 10668
rect 10735 10628 11428 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 11112 10560 11161 10588
rect 11112 10548 11118 10560
rect 11149 10557 11161 10560
rect 11195 10588 11207 10591
rect 11808 10588 11836 10696
rect 12437 10693 12449 10696
rect 12483 10693 12495 10727
rect 12437 10687 12495 10693
rect 16574 10684 16580 10736
rect 16632 10724 16638 10736
rect 18049 10727 18107 10733
rect 18049 10724 18061 10727
rect 16632 10696 18061 10724
rect 16632 10684 16638 10696
rect 18049 10693 18061 10696
rect 18095 10693 18107 10727
rect 18049 10687 18107 10693
rect 12342 10616 12348 10668
rect 12400 10656 12406 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12400 10628 13001 10656
rect 12400 10616 12406 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 14550 10656 14556 10668
rect 13771 10628 14556 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 12894 10588 12900 10600
rect 11195 10560 11836 10588
rect 12855 10560 12900 10588
rect 11195 10557 11207 10560
rect 11149 10551 11207 10557
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 11808 10492 12817 10520
rect 11808 10464 11836 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11241 10455 11299 10461
rect 11241 10452 11253 10455
rect 10928 10424 11253 10452
rect 10928 10412 10934 10424
rect 11241 10421 11253 10424
rect 11287 10421 11299 10455
rect 11790 10452 11796 10464
rect 11751 10424 11796 10452
rect 11241 10415 11299 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 12158 10452 12164 10464
rect 12071 10424 12164 10452
rect 12158 10412 12164 10424
rect 12216 10452 12222 10464
rect 12912 10452 12940 10548
rect 12216 10424 12940 10452
rect 12216 10412 12222 10424
rect 13446 10412 13452 10464
rect 13504 10452 13510 10464
rect 13740 10452 13768 10619
rect 14550 10616 14556 10628
rect 14608 10656 14614 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14608 10628 14657 10656
rect 14608 10616 14614 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14826 10656 14832 10668
rect 14787 10628 14832 10656
rect 14645 10619 14703 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 16114 10656 16120 10668
rect 15335 10628 16120 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 16114 10616 16120 10628
rect 16172 10656 16178 10668
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 16172 10628 16221 10656
rect 16172 10616 16178 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10656 16451 10659
rect 16666 10656 16672 10668
rect 16439 10628 16672 10656
rect 16439 10625 16451 10628
rect 16393 10619 16451 10625
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 18046 10588 18052 10600
rect 16908 10560 18052 10588
rect 16908 10548 16914 10560
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 18156 10588 18184 10764
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 19518 10792 19524 10804
rect 19479 10764 19524 10792
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 19702 10792 19708 10804
rect 19663 10764 19708 10792
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 23198 10752 23204 10804
rect 23256 10792 23262 10804
rect 23385 10795 23443 10801
rect 23385 10792 23397 10795
rect 23256 10764 23397 10792
rect 23256 10752 23262 10764
rect 23385 10761 23397 10764
rect 23431 10761 23443 10795
rect 23385 10755 23443 10761
rect 21358 10684 21364 10736
rect 21416 10724 21422 10736
rect 21416 10696 21496 10724
rect 21416 10684 21422 10696
rect 18690 10656 18696 10668
rect 18603 10628 18696 10656
rect 18690 10616 18696 10628
rect 18748 10656 18754 10668
rect 18748 10628 19196 10656
rect 18748 10616 18754 10628
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 18156 10560 18429 10588
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 15657 10523 15715 10529
rect 15657 10489 15669 10523
rect 15703 10520 15715 10523
rect 15838 10520 15844 10532
rect 15703 10492 15844 10520
rect 15703 10489 15715 10492
rect 15657 10483 15715 10489
rect 15838 10480 15844 10492
rect 15896 10520 15902 10532
rect 15896 10492 16160 10520
rect 15896 10480 15902 10492
rect 16132 10464 16160 10492
rect 16390 10480 16396 10532
rect 16448 10520 16454 10532
rect 17405 10523 17463 10529
rect 17405 10520 17417 10523
rect 16448 10492 17417 10520
rect 16448 10480 16454 10492
rect 17405 10489 17417 10492
rect 17451 10520 17463 10523
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 17451 10492 18521 10520
rect 17451 10489 17463 10492
rect 17405 10483 17463 10489
rect 18509 10489 18521 10492
rect 18555 10520 18567 10523
rect 18690 10520 18696 10532
rect 18555 10492 18696 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 18690 10480 18696 10492
rect 18748 10480 18754 10532
rect 13504 10424 13768 10452
rect 13504 10412 13510 10424
rect 13998 10412 14004 10464
rect 14056 10452 14062 10464
rect 14093 10455 14151 10461
rect 14093 10452 14105 10455
rect 14056 10424 14105 10452
rect 14056 10412 14062 10424
rect 14093 10421 14105 10424
rect 14139 10452 14151 10455
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 14139 10424 14565 10452
rect 14139 10421 14151 10424
rect 14093 10415 14151 10421
rect 14553 10421 14565 10424
rect 14599 10452 14611 10455
rect 14826 10452 14832 10464
rect 14599 10424 14832 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 15746 10452 15752 10464
rect 15707 10424 15752 10452
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 16114 10452 16120 10464
rect 16075 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 19168 10461 19196 10628
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19981 10659 20039 10665
rect 19981 10656 19993 10659
rect 19484 10628 19993 10656
rect 19484 10616 19490 10628
rect 19981 10625 19993 10628
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 19886 10588 19892 10600
rect 19847 10560 19892 10588
rect 19886 10548 19892 10560
rect 19944 10548 19950 10600
rect 21468 10597 21496 10696
rect 21634 10656 21640 10668
rect 21595 10628 21640 10656
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 22094 10616 22100 10668
rect 22152 10656 22158 10668
rect 22557 10659 22615 10665
rect 22557 10656 22569 10659
rect 22152 10628 22569 10656
rect 22152 10616 22158 10628
rect 22557 10625 22569 10628
rect 22603 10625 22615 10659
rect 23400 10656 23428 10755
rect 23934 10752 23940 10804
rect 23992 10792 23998 10804
rect 25222 10792 25228 10804
rect 23992 10764 25228 10792
rect 23992 10752 23998 10764
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 25314 10752 25320 10804
rect 25372 10792 25378 10804
rect 25777 10795 25835 10801
rect 25777 10792 25789 10795
rect 25372 10764 25789 10792
rect 25372 10752 25378 10764
rect 25777 10761 25789 10764
rect 25823 10761 25835 10795
rect 25777 10755 25835 10761
rect 24302 10656 24308 10668
rect 23400 10628 24308 10656
rect 22557 10619 22615 10625
rect 24302 10616 24308 10628
rect 24360 10616 24366 10668
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 25317 10659 25375 10665
rect 25317 10656 25329 10659
rect 24912 10628 25329 10656
rect 24912 10616 24918 10628
rect 25317 10625 25329 10628
rect 25363 10625 25375 10659
rect 25317 10619 25375 10625
rect 21453 10591 21511 10597
rect 21453 10557 21465 10591
rect 21499 10588 21511 10591
rect 24121 10591 24179 10597
rect 21499 10560 22140 10588
rect 21499 10557 21511 10560
rect 21453 10551 21511 10557
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 19334 10452 19340 10464
rect 19199 10424 19340 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 19904 10452 19932 10548
rect 20533 10523 20591 10529
rect 20533 10489 20545 10523
rect 20579 10520 20591 10523
rect 20901 10523 20959 10529
rect 20901 10520 20913 10523
rect 20579 10492 20913 10520
rect 20579 10489 20591 10492
rect 20533 10483 20591 10489
rect 20901 10489 20913 10492
rect 20947 10520 20959 10523
rect 20947 10492 21404 10520
rect 20947 10489 20959 10492
rect 20901 10483 20959 10489
rect 20438 10452 20444 10464
rect 19904 10424 20444 10452
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 20993 10455 21051 10461
rect 20993 10421 21005 10455
rect 21039 10452 21051 10455
rect 21174 10452 21180 10464
rect 21039 10424 21180 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 21376 10461 21404 10492
rect 21361 10455 21419 10461
rect 21361 10421 21373 10455
rect 21407 10452 21419 10455
rect 21450 10452 21456 10464
rect 21407 10424 21456 10452
rect 21407 10421 21419 10424
rect 21361 10415 21419 10421
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 22112 10461 22140 10560
rect 24121 10557 24133 10591
rect 24167 10588 24179 10591
rect 24210 10588 24216 10600
rect 24167 10560 24216 10588
rect 24167 10557 24179 10560
rect 24121 10551 24179 10557
rect 24210 10548 24216 10560
rect 24268 10588 24274 10600
rect 24765 10591 24823 10597
rect 24765 10588 24777 10591
rect 24268 10560 24777 10588
rect 24268 10548 24274 10560
rect 24765 10557 24777 10560
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 23106 10480 23112 10532
rect 23164 10520 23170 10532
rect 23290 10520 23296 10532
rect 23164 10492 23296 10520
rect 23164 10480 23170 10492
rect 23290 10480 23296 10492
rect 23348 10480 23354 10532
rect 22097 10455 22155 10461
rect 22097 10421 22109 10455
rect 22143 10452 22155 10455
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 22143 10424 22477 10452
rect 22143 10421 22155 10424
rect 22097 10415 22155 10421
rect 22465 10421 22477 10424
rect 22511 10452 22523 10455
rect 22830 10452 22836 10464
rect 22511 10424 22836 10452
rect 22511 10421 22523 10424
rect 22465 10415 22523 10421
rect 22830 10412 22836 10424
rect 22888 10412 22894 10464
rect 23014 10452 23020 10464
rect 22975 10424 23020 10452
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 23658 10412 23664 10464
rect 23716 10452 23722 10464
rect 23753 10455 23811 10461
rect 23753 10452 23765 10455
rect 23716 10424 23765 10452
rect 23716 10412 23722 10424
rect 23753 10421 23765 10424
rect 23799 10421 23811 10455
rect 23753 10415 23811 10421
rect 24210 10412 24216 10464
rect 24268 10452 24274 10464
rect 24268 10424 24313 10452
rect 24268 10412 24274 10424
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 12710 10248 12716 10260
rect 11480 10220 12716 10248
rect 11480 10208 11486 10220
rect 12710 10208 12716 10220
rect 12768 10248 12774 10260
rect 13265 10251 13323 10257
rect 13265 10248 13277 10251
rect 12768 10220 13277 10248
rect 12768 10208 12774 10220
rect 13265 10217 13277 10220
rect 13311 10217 13323 10251
rect 14734 10248 14740 10260
rect 14695 10220 14740 10248
rect 13265 10211 13323 10217
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 16022 10248 16028 10260
rect 15611 10220 16028 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16117 10251 16175 10257
rect 16117 10217 16129 10251
rect 16163 10248 16175 10251
rect 16206 10248 16212 10260
rect 16163 10220 16212 10248
rect 16163 10217 16175 10220
rect 16117 10211 16175 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 16632 10220 16681 10248
rect 16632 10208 16638 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 16669 10211 16727 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18230 10248 18236 10260
rect 18191 10220 18236 10248
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 18966 10208 18972 10260
rect 19024 10248 19030 10260
rect 19245 10251 19303 10257
rect 19245 10248 19257 10251
rect 19024 10220 19257 10248
rect 19024 10208 19030 10220
rect 19245 10217 19257 10220
rect 19291 10217 19303 10251
rect 19245 10211 19303 10217
rect 19613 10251 19671 10257
rect 19613 10217 19625 10251
rect 19659 10248 19671 10251
rect 20162 10248 20168 10260
rect 19659 10220 20168 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 21082 10208 21088 10260
rect 21140 10248 21146 10260
rect 21266 10248 21272 10260
rect 21140 10220 21272 10248
rect 21140 10208 21146 10220
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21361 10251 21419 10257
rect 21361 10217 21373 10251
rect 21407 10248 21419 10251
rect 21542 10248 21548 10260
rect 21407 10220 21548 10248
rect 21407 10217 21419 10220
rect 21361 10211 21419 10217
rect 21542 10208 21548 10220
rect 21600 10208 21606 10260
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22373 10251 22431 10257
rect 22373 10248 22385 10251
rect 22060 10220 22385 10248
rect 22060 10208 22066 10220
rect 22373 10217 22385 10220
rect 22419 10248 22431 10251
rect 22646 10248 22652 10260
rect 22419 10220 22652 10248
rect 22419 10217 22431 10220
rect 22373 10211 22431 10217
rect 22646 10208 22652 10220
rect 22704 10248 22710 10260
rect 22741 10251 22799 10257
rect 22741 10248 22753 10251
rect 22704 10220 22753 10248
rect 22704 10208 22710 10220
rect 22741 10217 22753 10220
rect 22787 10217 22799 10251
rect 22922 10248 22928 10260
rect 22883 10220 22928 10248
rect 22741 10211 22799 10217
rect 11882 10180 11888 10192
rect 11348 10152 11888 10180
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 11348 10053 11376 10152
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 14185 10183 14243 10189
rect 14185 10149 14197 10183
rect 14231 10180 14243 10183
rect 14642 10180 14648 10192
rect 14231 10152 14648 10180
rect 14231 10149 14243 10152
rect 14185 10143 14243 10149
rect 14642 10140 14648 10152
rect 14700 10140 14706 10192
rect 17494 10140 17500 10192
rect 17552 10180 17558 10192
rect 17589 10183 17647 10189
rect 17589 10180 17601 10183
rect 17552 10152 17601 10180
rect 17552 10140 17558 10152
rect 17589 10149 17601 10152
rect 17635 10149 17647 10183
rect 22756 10180 22784 10211
rect 22922 10208 22928 10220
rect 22980 10208 22986 10260
rect 23842 10248 23848 10260
rect 23755 10220 23848 10248
rect 23842 10208 23848 10220
rect 23900 10248 23906 10260
rect 24210 10248 24216 10260
rect 23900 10220 24216 10248
rect 23900 10208 23906 10220
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 24302 10208 24308 10260
rect 24360 10248 24366 10260
rect 25317 10251 25375 10257
rect 25317 10248 25329 10251
rect 24360 10220 25329 10248
rect 24360 10208 24366 10220
rect 25317 10217 25329 10220
rect 25363 10217 25375 10251
rect 25317 10211 25375 10217
rect 23385 10183 23443 10189
rect 23385 10180 23397 10183
rect 22756 10152 23397 10180
rect 17589 10143 17647 10149
rect 23385 10149 23397 10152
rect 23431 10180 23443 10183
rect 23431 10152 23980 10180
rect 23431 10149 23443 10152
rect 23385 10143 23443 10149
rect 11600 10115 11658 10121
rect 11600 10081 11612 10115
rect 11646 10112 11658 10115
rect 12342 10112 12348 10124
rect 11646 10084 12348 10112
rect 11646 10081 11658 10084
rect 11600 10075 11658 10081
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 14090 10112 14096 10124
rect 14051 10084 14096 10112
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 16022 10112 16028 10124
rect 15983 10084 16028 10112
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 19242 10112 19248 10124
rect 18831 10084 19248 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 19705 10115 19763 10121
rect 19705 10081 19717 10115
rect 19751 10112 19763 10115
rect 19978 10112 19984 10124
rect 19751 10084 19984 10112
rect 19751 10081 19763 10084
rect 19705 10075 19763 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 21140 10084 21281 10112
rect 21140 10072 21146 10084
rect 21269 10081 21281 10084
rect 21315 10112 21327 10115
rect 21450 10112 21456 10124
rect 21315 10084 21456 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 23952 10121 23980 10152
rect 23937 10115 23995 10121
rect 23937 10081 23949 10115
rect 23983 10081 23995 10115
rect 23937 10075 23995 10081
rect 24204 10115 24262 10121
rect 24204 10081 24216 10115
rect 24250 10112 24262 10115
rect 24946 10112 24952 10124
rect 24250 10084 24952 10112
rect 24250 10081 24262 10084
rect 24204 10075 24262 10081
rect 24946 10072 24952 10084
rect 25004 10072 25010 10124
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 11296 10016 11345 10044
rect 11296 10004 11302 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10044 16359 10047
rect 16666 10044 16672 10056
rect 16347 10016 16672 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 15105 9979 15163 9985
rect 15105 9945 15117 9979
rect 15151 9976 15163 9979
rect 16316 9976 16344 10007
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17862 10044 17868 10056
rect 17823 10016 17868 10044
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20070 10044 20076 10056
rect 19935 10016 20076 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 15151 9948 16344 9976
rect 15151 9945 15163 9948
rect 15105 9939 15163 9945
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 17221 9979 17279 9985
rect 17221 9976 17233 9979
rect 16632 9948 17233 9976
rect 16632 9936 16638 9948
rect 17221 9945 17233 9948
rect 17267 9945 17279 9979
rect 17221 9939 17279 9945
rect 19153 9979 19211 9985
rect 19153 9945 19165 9979
rect 19199 9976 19211 9979
rect 19904 9976 19932 10007
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21634 10044 21640 10056
rect 21591 10016 21640 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21634 10004 21640 10016
rect 21692 10004 21698 10056
rect 19199 9948 19932 9976
rect 19199 9945 19211 9948
rect 19153 9939 19211 9945
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 13909 9911 13967 9917
rect 13909 9908 13921 9911
rect 13872 9880 13921 9908
rect 13872 9868 13878 9880
rect 13909 9877 13921 9880
rect 13955 9908 13967 9911
rect 14182 9908 14188 9920
rect 13955 9880 14188 9908
rect 13955 9877 13967 9880
rect 13909 9871 13967 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 15657 9911 15715 9917
rect 15657 9877 15669 9911
rect 15703 9908 15715 9911
rect 15838 9908 15844 9920
rect 15703 9880 15844 9908
rect 15703 9877 15715 9880
rect 15657 9871 15715 9877
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 16942 9868 16948 9920
rect 17000 9908 17006 9920
rect 17129 9911 17187 9917
rect 17129 9908 17141 9911
rect 17000 9880 17141 9908
rect 17000 9868 17006 9880
rect 17129 9877 17141 9880
rect 17175 9908 17187 9911
rect 17678 9908 17684 9920
rect 17175 9880 17684 9908
rect 17175 9877 17187 9880
rect 17129 9871 17187 9877
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 20622 9908 20628 9920
rect 20583 9880 20628 9908
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 20901 9911 20959 9917
rect 20901 9877 20913 9911
rect 20947 9908 20959 9911
rect 20990 9908 20996 9920
rect 20947 9880 20996 9908
rect 20947 9877 20959 9880
rect 20901 9871 20959 9877
rect 20990 9868 20996 9880
rect 21048 9908 21054 9920
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 21048 9880 21925 9908
rect 21048 9868 21054 9880
rect 21913 9877 21925 9880
rect 21959 9877 21971 9911
rect 21913 9871 21971 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 10870 9664 10876 9716
rect 10928 9704 10934 9716
rect 10928 9676 12388 9704
rect 10928 9664 10934 9676
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11790 9568 11796 9580
rect 11379 9540 11796 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10594 9432 10600 9444
rect 10192 9404 10600 9432
rect 10192 9392 10198 9404
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 12360 9432 12388 9676
rect 13078 9664 13084 9716
rect 13136 9664 13142 9716
rect 16206 9704 16212 9716
rect 15120 9676 16212 9704
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12860 9540 13001 9568
rect 12860 9528 12866 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13096 9500 13124 9664
rect 13170 9596 13176 9648
rect 13228 9596 13234 9648
rect 15120 9645 15148 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 17310 9664 17316 9716
rect 17368 9704 17374 9716
rect 17773 9707 17831 9713
rect 17773 9704 17785 9707
rect 17368 9676 17785 9704
rect 17368 9664 17374 9676
rect 17773 9673 17785 9676
rect 17819 9673 17831 9707
rect 17773 9667 17831 9673
rect 20073 9707 20131 9713
rect 20073 9673 20085 9707
rect 20119 9704 20131 9707
rect 20162 9704 20168 9716
rect 20119 9676 20168 9704
rect 20119 9673 20131 9676
rect 20073 9667 20131 9673
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 21542 9704 21548 9716
rect 20640 9676 21548 9704
rect 15105 9639 15163 9645
rect 15105 9605 15117 9639
rect 15151 9605 15163 9639
rect 19426 9636 19432 9648
rect 19387 9608 19432 9636
rect 15105 9599 15163 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 20441 9639 20499 9645
rect 20441 9605 20453 9639
rect 20487 9636 20499 9639
rect 20640 9636 20668 9676
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 21634 9664 21640 9716
rect 21692 9704 21698 9716
rect 21913 9707 21971 9713
rect 21913 9704 21925 9707
rect 21692 9676 21925 9704
rect 21692 9664 21698 9676
rect 21913 9673 21925 9676
rect 21959 9673 21971 9707
rect 22646 9704 22652 9716
rect 22607 9676 22652 9704
rect 21913 9667 21971 9673
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 22830 9664 22836 9716
rect 22888 9704 22894 9716
rect 23842 9704 23848 9716
rect 22888 9676 23428 9704
rect 23803 9676 23848 9704
rect 22888 9664 22894 9676
rect 20487 9608 20668 9636
rect 20487 9605 20499 9608
rect 20441 9599 20499 9605
rect 13188 9568 13216 9596
rect 13262 9568 13268 9580
rect 13188 9540 13268 9568
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 14734 9568 14740 9580
rect 14647 9540 14740 9568
rect 14734 9528 14740 9540
rect 14792 9568 14798 9580
rect 15841 9571 15899 9577
rect 15841 9568 15853 9571
rect 14792 9540 15853 9568
rect 14792 9528 14798 9540
rect 15841 9537 15853 9540
rect 15887 9568 15899 9571
rect 16390 9568 16396 9580
rect 15887 9540 16396 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 16574 9568 16580 9580
rect 16500 9540 16580 9568
rect 13170 9500 13176 9512
rect 13096 9472 13176 9500
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 14415 9472 15669 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 15657 9469 15669 9472
rect 15703 9500 15715 9503
rect 16500 9500 16528 9540
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9568 17003 9571
rect 17770 9568 17776 9580
rect 16991 9540 17776 9568
rect 16991 9537 17003 9540
rect 16945 9531 17003 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 20990 9568 20996 9580
rect 20951 9540 20996 9568
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 21140 9540 21185 9568
rect 21140 9528 21146 9540
rect 21450 9528 21456 9580
rect 21508 9568 21514 9580
rect 21545 9571 21603 9577
rect 21545 9568 21557 9571
rect 21508 9540 21557 9568
rect 21508 9528 21514 9540
rect 21545 9537 21557 9540
rect 21591 9537 21603 9571
rect 21545 9531 21603 9537
rect 23400 9512 23428 9676
rect 23842 9664 23848 9676
rect 23900 9664 23906 9716
rect 24946 9704 24952 9716
rect 24907 9676 24952 9704
rect 24946 9664 24952 9676
rect 25004 9704 25010 9716
rect 25225 9707 25283 9713
rect 25225 9704 25237 9707
rect 25004 9676 25237 9704
rect 25004 9664 25010 9676
rect 25225 9673 25237 9676
rect 25271 9673 25283 9707
rect 25225 9667 25283 9673
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9568 24547 9571
rect 24946 9568 24952 9580
rect 24535 9540 24952 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 25406 9568 25412 9580
rect 25367 9540 25412 9568
rect 25406 9528 25412 9540
rect 25464 9528 25470 9580
rect 16666 9500 16672 9512
rect 15703 9472 16528 9500
rect 16579 9472 16672 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 16666 9460 16672 9472
rect 16724 9500 16730 9512
rect 17862 9500 17868 9512
rect 16724 9472 17868 9500
rect 16724 9460 16730 9472
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 18012 9472 18061 9500
rect 18012 9460 18018 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 20622 9460 20628 9512
rect 20680 9500 20686 9512
rect 20901 9503 20959 9509
rect 20901 9500 20913 9503
rect 20680 9472 20913 9500
rect 20680 9460 20686 9472
rect 20901 9469 20913 9472
rect 20947 9500 20959 9503
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 20947 9472 22109 9500
rect 20947 9469 20959 9472
rect 20901 9463 20959 9469
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 23382 9460 23388 9512
rect 23440 9460 23446 9512
rect 12360 9404 12480 9432
rect 11238 9364 11244 9376
rect 11199 9336 11244 9364
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11885 9367 11943 9373
rect 11885 9333 11897 9367
rect 11931 9364 11943 9367
rect 12253 9367 12311 9373
rect 12253 9364 12265 9367
rect 11931 9336 12265 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12253 9333 12265 9336
rect 12299 9364 12311 9367
rect 12342 9364 12348 9376
rect 12299 9336 12348 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 12452 9373 12480 9404
rect 12526 9392 12532 9444
rect 12584 9432 12590 9444
rect 12805 9435 12863 9441
rect 12805 9432 12817 9435
rect 12584 9404 12817 9432
rect 12584 9392 12590 9404
rect 12805 9401 12817 9404
rect 12851 9432 12863 9435
rect 13817 9435 13875 9441
rect 13817 9432 13829 9435
rect 12851 9404 13829 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 13817 9401 13829 9404
rect 13863 9401 13875 9435
rect 13817 9395 13875 9401
rect 15565 9435 15623 9441
rect 15565 9401 15577 9435
rect 15611 9432 15623 9435
rect 15746 9432 15752 9444
rect 15611 9404 15752 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 18230 9392 18236 9444
rect 18288 9441 18294 9444
rect 18288 9435 18352 9441
rect 18288 9401 18306 9435
rect 18340 9401 18352 9435
rect 23014 9432 23020 9444
rect 22975 9404 23020 9432
rect 18288 9395 18352 9401
rect 18288 9392 18294 9395
rect 23014 9392 23020 9404
rect 23072 9432 23078 9444
rect 24305 9435 24363 9441
rect 24305 9432 24317 9435
rect 23072 9404 24317 9432
rect 23072 9392 23078 9404
rect 24305 9401 24317 9404
rect 24351 9401 24363 9435
rect 24305 9395 24363 9401
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 12952 9336 13461 9364
rect 12952 9324 12958 9336
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15286 9364 15292 9376
rect 15243 9336 15292 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 16080 9336 16221 9364
rect 16080 9324 16086 9336
rect 16209 9333 16221 9336
rect 16255 9333 16267 9367
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 16209 9327 16267 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 20533 9367 20591 9373
rect 20533 9333 20545 9367
rect 20579 9364 20591 9367
rect 20622 9364 20628 9376
rect 20579 9336 20628 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 23474 9364 23480 9376
rect 23387 9336 23480 9364
rect 23474 9324 23480 9336
rect 23532 9364 23538 9376
rect 24210 9364 24216 9376
rect 23532 9336 24216 9364
rect 23532 9324 23538 9336
rect 24210 9324 24216 9336
rect 24268 9324 24274 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12802 9160 12808 9172
rect 12400 9132 12808 9160
rect 12400 9120 12406 9132
rect 12802 9120 12808 9132
rect 12860 9160 12866 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12860 9132 12909 9160
rect 12860 9120 12866 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 14001 9163 14059 9169
rect 14001 9129 14013 9163
rect 14047 9160 14059 9163
rect 14090 9160 14096 9172
rect 14047 9132 14096 9160
rect 14047 9129 14059 9132
rect 14001 9123 14059 9129
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 14829 9163 14887 9169
rect 14829 9129 14841 9163
rect 14875 9160 14887 9163
rect 15746 9160 15752 9172
rect 14875 9132 15752 9160
rect 14875 9129 14887 9132
rect 14829 9123 14887 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 17862 9160 17868 9172
rect 17635 9132 17868 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19429 9163 19487 9169
rect 19429 9160 19441 9163
rect 19392 9132 19441 9160
rect 19392 9120 19398 9132
rect 19429 9129 19441 9132
rect 19475 9129 19487 9163
rect 20070 9160 20076 9172
rect 20031 9132 20076 9160
rect 19429 9123 19487 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 20162 9120 20168 9172
rect 20220 9160 20226 9172
rect 20438 9160 20444 9172
rect 20220 9132 20444 9160
rect 20220 9120 20226 9132
rect 20438 9120 20444 9132
rect 20496 9160 20502 9172
rect 20533 9163 20591 9169
rect 20533 9160 20545 9163
rect 20496 9132 20545 9160
rect 20496 9120 20502 9132
rect 20533 9129 20545 9132
rect 20579 9129 20591 9163
rect 20533 9123 20591 9129
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 21818 9160 21824 9172
rect 21232 9132 21824 9160
rect 21232 9120 21238 9132
rect 21818 9120 21824 9132
rect 21876 9160 21882 9172
rect 22833 9163 22891 9169
rect 22833 9160 22845 9163
rect 21876 9132 22845 9160
rect 21876 9120 21882 9132
rect 22833 9129 22845 9132
rect 22879 9129 22891 9163
rect 22833 9123 22891 9129
rect 24026 9120 24032 9172
rect 24084 9160 24090 9172
rect 24305 9163 24363 9169
rect 24305 9160 24317 9163
rect 24084 9132 24317 9160
rect 24084 9120 24090 9132
rect 24305 9129 24317 9132
rect 24351 9129 24363 9163
rect 24305 9123 24363 9129
rect 15832 9095 15890 9101
rect 15832 9061 15844 9095
rect 15878 9092 15890 9095
rect 16114 9092 16120 9104
rect 15878 9064 16120 9092
rect 15878 9061 15890 9064
rect 15832 9055 15890 9061
rect 16114 9052 16120 9064
rect 16172 9092 16178 9104
rect 16666 9092 16672 9104
rect 16172 9064 16672 9092
rect 16172 9052 16178 9064
rect 16666 9052 16672 9064
rect 16724 9052 16730 9104
rect 22002 9092 22008 9104
rect 20916 9064 22008 9092
rect 20916 9036 20944 9064
rect 22002 9052 22008 9064
rect 22060 9052 22066 9104
rect 11422 8984 11428 9036
rect 11480 9024 11486 9036
rect 11773 9027 11831 9033
rect 11773 9024 11785 9027
rect 11480 8996 11785 9024
rect 11480 8984 11486 8996
rect 11773 8993 11785 8996
rect 11819 8993 11831 9027
rect 11773 8987 11831 8993
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 16206 9024 16212 9036
rect 15151 8996 16212 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 18322 9033 18328 9036
rect 18316 8987 18328 9033
rect 18380 9024 18386 9036
rect 20714 9024 20720 9036
rect 18380 8996 18416 9024
rect 20675 8996 20720 9024
rect 18322 8984 18328 8987
rect 18380 8984 18386 8996
rect 20714 8984 20720 8996
rect 20772 8984 20778 9036
rect 20898 9024 20904 9036
rect 20859 8996 20904 9024
rect 20898 8984 20904 8996
rect 20956 8984 20962 9036
rect 20990 8984 20996 9036
rect 21048 9024 21054 9036
rect 21157 9027 21215 9033
rect 21157 9024 21169 9027
rect 21048 8996 21169 9024
rect 21048 8984 21054 8996
rect 21157 8993 21169 8996
rect 21203 9024 21215 9027
rect 21634 9024 21640 9036
rect 21203 8996 21640 9024
rect 21203 8993 21215 8996
rect 21157 8987 21215 8993
rect 21634 8984 21640 8996
rect 21692 8984 21698 9036
rect 23106 8984 23112 9036
rect 23164 9024 23170 9036
rect 24213 9027 24271 9033
rect 24213 9024 24225 9027
rect 23164 8996 24225 9024
rect 23164 8984 23170 8996
rect 24213 8993 24225 8996
rect 24259 9024 24271 9027
rect 24762 9024 24768 9036
rect 24259 8996 24768 9024
rect 24259 8993 24271 8996
rect 24213 8987 24271 8993
rect 24762 8984 24768 8996
rect 24820 8984 24826 9036
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 11238 8956 11244 8968
rect 10376 8928 11244 8956
rect 10376 8916 10382 8928
rect 11238 8916 11244 8928
rect 11296 8956 11302 8968
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 11296 8928 11529 8956
rect 11296 8916 11302 8928
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 14240 8928 14381 8956
rect 14240 8916 14246 8928
rect 14369 8925 14381 8928
rect 14415 8956 14427 8959
rect 15562 8956 15568 8968
rect 14415 8928 15568 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 17678 8916 17684 8968
rect 17736 8956 17742 8968
rect 18046 8956 18052 8968
rect 17736 8928 18052 8956
rect 17736 8916 17742 8928
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 20070 8916 20076 8968
rect 20128 8956 20134 8968
rect 20254 8956 20260 8968
rect 20128 8928 20260 8956
rect 20128 8916 20134 8928
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 24397 8959 24455 8965
rect 24397 8925 24409 8959
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 14090 8848 14096 8900
rect 14148 8888 14154 8900
rect 14550 8888 14556 8900
rect 14148 8860 14556 8888
rect 14148 8848 14154 8860
rect 14550 8848 14556 8860
rect 14608 8888 14614 8900
rect 14921 8891 14979 8897
rect 14921 8888 14933 8891
rect 14608 8860 14933 8888
rect 14608 8848 14614 8860
rect 14921 8857 14933 8860
rect 14967 8857 14979 8891
rect 14921 8851 14979 8857
rect 23753 8891 23811 8897
rect 23753 8857 23765 8891
rect 23799 8888 23811 8891
rect 23934 8888 23940 8900
rect 23799 8860 23940 8888
rect 23799 8857 23811 8860
rect 23753 8851 23811 8857
rect 23934 8848 23940 8860
rect 23992 8888 23998 8900
rect 24412 8888 24440 8919
rect 23992 8860 24440 8888
rect 23992 8848 23998 8860
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 11422 8820 11428 8832
rect 10919 8792 11428 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 15746 8820 15752 8832
rect 15528 8792 15752 8820
rect 15528 8780 15534 8792
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16482 8780 16488 8832
rect 16540 8820 16546 8832
rect 16945 8823 17003 8829
rect 16945 8820 16957 8823
rect 16540 8792 16957 8820
rect 16540 8780 16546 8792
rect 16945 8789 16957 8792
rect 16991 8789 17003 8823
rect 17954 8820 17960 8832
rect 17915 8792 17960 8820
rect 16945 8783 17003 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 20254 8780 20260 8832
rect 20312 8820 20318 8832
rect 20349 8823 20407 8829
rect 20349 8820 20361 8823
rect 20312 8792 20361 8820
rect 20312 8780 20318 8792
rect 20349 8789 20361 8792
rect 20395 8789 20407 8823
rect 22278 8820 22284 8832
rect 22239 8792 22284 8820
rect 20349 8783 20407 8789
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 23382 8820 23388 8832
rect 23343 8792 23388 8820
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 23842 8820 23848 8832
rect 23803 8792 23848 8820
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 10318 8616 10324 8628
rect 10279 8588 10324 8616
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10778 8616 10784 8628
rect 10739 8588 10784 8616
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 12526 8616 12532 8628
rect 12487 8588 12532 8616
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 13262 8616 13268 8628
rect 13136 8588 13268 8616
rect 13136 8576 13142 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 16114 8616 16120 8628
rect 16075 8588 16120 8616
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 16485 8619 16543 8625
rect 16485 8616 16497 8619
rect 16264 8588 16497 8616
rect 16264 8576 16270 8588
rect 16485 8585 16497 8588
rect 16531 8616 16543 8619
rect 17586 8616 17592 8628
rect 16531 8588 17592 8616
rect 16531 8585 16543 8588
rect 16485 8579 16543 8585
rect 17586 8576 17592 8588
rect 17644 8616 17650 8628
rect 17862 8616 17868 8628
rect 17644 8588 17868 8616
rect 17644 8576 17650 8588
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 18322 8576 18328 8588
rect 18380 8616 18386 8628
rect 20349 8619 20407 8625
rect 20349 8616 20361 8619
rect 18380 8588 20361 8616
rect 18380 8576 18386 8588
rect 20349 8585 20361 8588
rect 20395 8616 20407 8619
rect 20806 8616 20812 8628
rect 20395 8588 20812 8616
rect 20395 8585 20407 8588
rect 20349 8579 20407 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 23106 8616 23112 8628
rect 23067 8588 23112 8616
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 24026 8616 24032 8628
rect 23523 8588 24032 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 24026 8576 24032 8588
rect 24084 8576 24090 8628
rect 24946 8576 24952 8628
rect 25004 8616 25010 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25004 8588 25237 8616
rect 25004 8576 25010 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 25225 8579 25283 8585
rect 11977 8551 12035 8557
rect 11977 8517 11989 8551
rect 12023 8548 12035 8551
rect 12894 8548 12900 8560
rect 12023 8520 12900 8548
rect 12023 8517 12035 8520
rect 11977 8511 12035 8517
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 15473 8551 15531 8557
rect 15473 8517 15485 8551
rect 15519 8548 15531 8551
rect 15930 8548 15936 8560
rect 15519 8520 15936 8548
rect 15519 8517 15531 8520
rect 15473 8511 15531 8517
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 11422 8480 11428 8492
rect 11335 8452 11428 8480
rect 11422 8440 11428 8452
rect 11480 8480 11486 8492
rect 12526 8480 12532 8492
rect 11480 8452 12532 8480
rect 11480 8440 11486 8452
rect 12526 8440 12532 8452
rect 12584 8480 12590 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 12584 8452 13185 8480
rect 12584 8440 12590 8452
rect 13173 8449 13185 8452
rect 13219 8480 13231 8483
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 13219 8452 13553 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8480 14059 8483
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 14047 8452 14228 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 11330 8372 11336 8424
rect 11388 8412 11394 8424
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11388 8384 11805 8412
rect 11388 8372 11394 8384
rect 11793 8381 11805 8384
rect 11839 8412 11851 8415
rect 11977 8415 12035 8421
rect 11977 8412 11989 8415
rect 11839 8384 11989 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 11977 8381 11989 8384
rect 12023 8381 12035 8415
rect 11977 8375 12035 8381
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12299 8384 13001 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12989 8381 13001 8384
rect 13035 8412 13047 8415
rect 13262 8412 13268 8424
rect 13035 8384 13268 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 14090 8412 14096 8424
rect 14051 8384 14096 8412
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14200 8412 14228 8452
rect 21284 8452 22017 8480
rect 14360 8415 14418 8421
rect 14360 8412 14372 8415
rect 14200 8384 14372 8412
rect 14360 8381 14372 8384
rect 14406 8412 14418 8415
rect 14734 8412 14740 8424
rect 14406 8384 14740 8412
rect 14406 8381 14418 8384
rect 14360 8375 14418 8381
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 18969 8415 19027 8421
rect 18969 8412 18981 8415
rect 17420 8384 18981 8412
rect 10689 8347 10747 8353
rect 10689 8313 10701 8347
rect 10735 8344 10747 8347
rect 11241 8347 11299 8353
rect 11241 8344 11253 8347
rect 10735 8316 11253 8344
rect 10735 8313 10747 8316
rect 10689 8307 10747 8313
rect 11241 8313 11253 8316
rect 11287 8344 11299 8347
rect 12618 8344 12624 8356
rect 11287 8316 12624 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 12618 8304 12624 8316
rect 12676 8304 12682 8356
rect 12894 8344 12900 8356
rect 12855 8316 12900 8344
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 16577 8347 16635 8353
rect 16577 8344 16589 8347
rect 16540 8316 16589 8344
rect 16540 8304 16546 8316
rect 16577 8313 16589 8316
rect 16623 8313 16635 8347
rect 16577 8307 16635 8313
rect 17420 8288 17448 8384
rect 18969 8381 18981 8384
rect 19015 8381 19027 8415
rect 21082 8412 21088 8424
rect 18969 8375 19027 8381
rect 20272 8384 21088 8412
rect 20272 8356 20300 8384
rect 21082 8372 21088 8384
rect 21140 8412 21146 8424
rect 21284 8421 21312 8452
rect 22005 8449 22017 8452
rect 22051 8480 22063 8483
rect 22278 8480 22284 8492
rect 22051 8452 22284 8480
rect 22051 8449 22063 8452
rect 22005 8443 22063 8449
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 21269 8415 21327 8421
rect 21269 8412 21281 8415
rect 21140 8384 21281 8412
rect 21140 8372 21146 8384
rect 21269 8381 21281 8384
rect 21315 8381 21327 8415
rect 21818 8412 21824 8424
rect 21779 8384 21824 8412
rect 21269 8375 21327 8381
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 22554 8372 22560 8424
rect 22612 8412 22618 8424
rect 23382 8412 23388 8424
rect 22612 8384 23388 8412
rect 22612 8372 22618 8384
rect 23382 8372 23388 8384
rect 23440 8412 23446 8424
rect 23845 8415 23903 8421
rect 23845 8412 23857 8415
rect 23440 8384 23857 8412
rect 23440 8372 23446 8384
rect 23845 8381 23857 8384
rect 23891 8381 23903 8415
rect 23845 8375 23903 8381
rect 18877 8347 18935 8353
rect 18877 8313 18889 8347
rect 18923 8344 18935 8347
rect 19214 8347 19272 8353
rect 19214 8344 19226 8347
rect 18923 8316 19226 8344
rect 18923 8313 18935 8316
rect 18877 8307 18935 8313
rect 19214 8313 19226 8316
rect 19260 8344 19272 8347
rect 20254 8344 20260 8356
rect 19260 8316 20260 8344
rect 19260 8313 19272 8316
rect 19214 8307 19272 8313
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 24118 8353 24124 8356
rect 21913 8347 21971 8353
rect 21913 8344 21925 8347
rect 20640 8316 21925 8344
rect 10870 8236 10876 8288
rect 10928 8276 10934 8288
rect 11149 8279 11207 8285
rect 11149 8276 11161 8279
rect 10928 8248 11161 8276
rect 10928 8236 10934 8248
rect 11149 8245 11161 8248
rect 11195 8245 11207 8279
rect 11149 8239 11207 8245
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 17034 8276 17040 8288
rect 12032 8248 17040 8276
rect 12032 8236 12038 8248
rect 17034 8236 17040 8248
rect 17092 8236 17098 8288
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 20438 8236 20444 8288
rect 20496 8276 20502 8288
rect 20640 8276 20668 8316
rect 21913 8313 21925 8316
rect 21959 8344 21971 8347
rect 22465 8347 22523 8353
rect 22465 8344 22477 8347
rect 21959 8316 22477 8344
rect 21959 8313 21971 8316
rect 21913 8307 21971 8313
rect 22465 8313 22477 8316
rect 22511 8313 22523 8347
rect 24112 8344 24124 8353
rect 24079 8316 24124 8344
rect 22465 8307 22523 8313
rect 24112 8307 24124 8316
rect 24118 8304 24124 8307
rect 24176 8304 24182 8356
rect 20990 8276 20996 8288
rect 20496 8248 20668 8276
rect 20951 8248 20996 8276
rect 20496 8236 20502 8248
rect 20990 8236 20996 8248
rect 21048 8236 21054 8288
rect 21450 8276 21456 8288
rect 21411 8248 21456 8276
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 14001 8075 14059 8081
rect 14001 8041 14013 8075
rect 14047 8072 14059 8075
rect 14274 8072 14280 8084
rect 14047 8044 14280 8072
rect 14047 8041 14059 8044
rect 14001 8035 14059 8041
rect 14274 8032 14280 8044
rect 14332 8072 14338 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 14332 8044 15301 8072
rect 14332 8032 14338 8044
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 15289 8035 15347 8041
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 16114 8072 16120 8084
rect 15703 8044 16120 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16114 8032 16120 8044
rect 16172 8072 16178 8084
rect 16482 8072 16488 8084
rect 16172 8044 16488 8072
rect 16172 8032 16178 8044
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 17773 8075 17831 8081
rect 17773 8041 17785 8075
rect 17819 8072 17831 8075
rect 17862 8072 17868 8084
rect 17819 8044 17868 8072
rect 17819 8041 17831 8044
rect 17773 8035 17831 8041
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 18046 8072 18052 8084
rect 18007 8044 18052 8072
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18693 8075 18751 8081
rect 18693 8041 18705 8075
rect 18739 8072 18751 8075
rect 18782 8072 18788 8084
rect 18739 8044 18788 8072
rect 18739 8041 18751 8044
rect 18693 8035 18751 8041
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 20772 8044 21281 8072
rect 20772 8032 20778 8044
rect 21269 8041 21281 8044
rect 21315 8072 21327 8075
rect 22186 8072 22192 8084
rect 21315 8044 22192 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 22186 8032 22192 8044
rect 22244 8032 22250 8084
rect 23934 8072 23940 8084
rect 23895 8044 23940 8072
rect 23934 8032 23940 8044
rect 23992 8032 23998 8084
rect 24854 8032 24860 8084
rect 24912 8072 24918 8084
rect 25041 8075 25099 8081
rect 25041 8072 25053 8075
rect 24912 8044 25053 8072
rect 24912 8032 24918 8044
rect 25041 8041 25053 8044
rect 25087 8041 25099 8075
rect 25041 8035 25099 8041
rect 10137 8007 10195 8013
rect 10137 7973 10149 8007
rect 10183 8004 10195 8007
rect 11146 8004 11152 8016
rect 10183 7976 11152 8004
rect 10183 7973 10195 7976
rect 10137 7967 10195 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 14090 8004 14096 8016
rect 14003 7976 14096 8004
rect 14090 7964 14096 7976
rect 14148 8004 14154 8016
rect 15102 8004 15108 8016
rect 14148 7976 15108 8004
rect 14148 7964 14154 7976
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 15749 8007 15807 8013
rect 15749 7973 15761 8007
rect 15795 8004 15807 8007
rect 15838 8004 15844 8016
rect 15795 7976 15844 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 17221 8007 17279 8013
rect 17221 7973 17233 8007
rect 17267 8004 17279 8007
rect 19242 8004 19248 8016
rect 17267 7976 19248 8004
rect 17267 7973 17279 7976
rect 17221 7967 17279 7973
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 19705 8007 19763 8013
rect 19705 7973 19717 8007
rect 19751 8004 19763 8007
rect 21361 8007 21419 8013
rect 21361 8004 21373 8007
rect 19751 7976 21373 8004
rect 19751 7973 19763 7976
rect 19705 7967 19763 7973
rect 21361 7973 21373 7976
rect 21407 8004 21419 8007
rect 21450 8004 21456 8016
rect 21407 7976 21456 8004
rect 21407 7973 21419 7976
rect 21361 7967 21419 7973
rect 21450 7964 21456 7976
rect 21508 7964 21514 8016
rect 9858 7936 9864 7948
rect 9819 7908 9864 7936
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11405 7939 11463 7945
rect 11405 7936 11417 7939
rect 11296 7908 11417 7936
rect 11296 7896 11302 7908
rect 11405 7905 11417 7908
rect 11451 7905 11463 7939
rect 11405 7899 11463 7905
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 15620 7908 16313 7936
rect 15620 7896 15626 7908
rect 16301 7905 16313 7908
rect 16347 7936 16359 7939
rect 18046 7936 18052 7948
rect 16347 7908 18052 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18598 7936 18604 7948
rect 18559 7908 18604 7936
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 22462 7896 22468 7948
rect 22520 7936 22526 7948
rect 22813 7939 22871 7945
rect 22813 7936 22825 7939
rect 22520 7908 22825 7936
rect 22520 7896 22526 7908
rect 22813 7905 22825 7908
rect 22859 7905 22871 7939
rect 22813 7899 22871 7905
rect 11146 7868 11152 7880
rect 11107 7840 11152 7868
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14366 7868 14372 7880
rect 14323 7840 14372 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14366 7828 14372 7840
rect 14424 7828 14430 7880
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7868 15991 7871
rect 16390 7868 16396 7880
rect 15979 7840 16396 7868
rect 15979 7837 15991 7840
rect 15933 7831 15991 7837
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 18322 7760 18328 7812
rect 18380 7800 18386 7812
rect 18800 7800 18828 7831
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 19797 7871 19855 7877
rect 19797 7868 19809 7871
rect 19484 7840 19809 7868
rect 19484 7828 19490 7840
rect 19797 7837 19809 7840
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 21450 7868 21456 7880
rect 20864 7840 21456 7868
rect 20864 7828 20870 7840
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 22554 7868 22560 7880
rect 22515 7840 22560 7868
rect 22554 7828 22560 7840
rect 22612 7828 22618 7880
rect 18380 7772 18828 7800
rect 18380 7760 18386 7772
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 22152 7772 22600 7800
rect 22152 7760 22158 7772
rect 10870 7732 10876 7744
rect 10831 7704 10876 7732
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 13081 7735 13139 7741
rect 13081 7732 13093 7735
rect 12952 7704 13093 7732
rect 12952 7692 12958 7704
rect 13081 7701 13093 7704
rect 13127 7701 13139 7735
rect 13630 7732 13636 7744
rect 13591 7704 13636 7732
rect 13081 7695 13139 7701
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 15105 7735 15163 7741
rect 15105 7732 15117 7735
rect 14056 7704 15117 7732
rect 14056 7692 14062 7704
rect 15105 7701 15117 7704
rect 15151 7732 15163 7735
rect 15746 7732 15752 7744
rect 15151 7704 15752 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 18233 7735 18291 7741
rect 18233 7701 18245 7735
rect 18279 7732 18291 7735
rect 18506 7732 18512 7744
rect 18279 7704 18512 7732
rect 18279 7701 18291 7704
rect 18233 7695 18291 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 20533 7735 20591 7741
rect 20533 7701 20545 7735
rect 20579 7732 20591 7735
rect 20622 7732 20628 7744
rect 20579 7704 20628 7732
rect 20579 7701 20591 7704
rect 20533 7695 20591 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 20898 7732 20904 7744
rect 20859 7704 20904 7732
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 22462 7732 22468 7744
rect 22423 7704 22468 7732
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 22572 7732 22600 7772
rect 22738 7732 22744 7744
rect 22572 7704 22744 7732
rect 22738 7692 22744 7704
rect 22796 7692 22802 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24489 7735 24547 7741
rect 24489 7732 24501 7735
rect 24176 7704 24501 7732
rect 24176 7692 24182 7704
rect 24489 7701 24501 7704
rect 24535 7701 24547 7735
rect 24489 7695 24547 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 9858 7528 9864 7540
rect 9447 7500 9864 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 11238 7528 11244 7540
rect 11199 7500 11244 7528
rect 11238 7488 11244 7500
rect 11296 7528 11302 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11296 7500 11805 7528
rect 11296 7488 11302 7500
rect 11793 7497 11805 7500
rect 11839 7528 11851 7531
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11839 7500 12173 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 12176 7392 12204 7491
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 14090 7528 14096 7540
rect 12492 7500 12537 7528
rect 14051 7500 14096 7528
rect 12492 7488 12498 7500
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 16114 7528 16120 7540
rect 16075 7500 16120 7528
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 16390 7528 16396 7540
rect 16351 7500 16396 7528
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 17862 7528 17868 7540
rect 17775 7500 17868 7528
rect 17862 7488 17868 7500
rect 17920 7528 17926 7540
rect 18598 7528 18604 7540
rect 17920 7500 18604 7528
rect 17920 7488 17926 7500
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 20438 7528 20444 7540
rect 20399 7500 20444 7528
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 21450 7528 21456 7540
rect 21411 7500 21456 7528
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 21818 7528 21824 7540
rect 21779 7500 21824 7528
rect 21818 7488 21824 7500
rect 21876 7528 21882 7540
rect 22002 7528 22008 7540
rect 21876 7500 22008 7528
rect 21876 7488 21882 7500
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 13725 7463 13783 7469
rect 13725 7429 13737 7463
rect 13771 7460 13783 7463
rect 14366 7460 14372 7472
rect 13771 7432 14372 7460
rect 13771 7429 13783 7432
rect 13725 7423 13783 7429
rect 14366 7420 14372 7432
rect 14424 7420 14430 7472
rect 15838 7420 15844 7472
rect 15896 7460 15902 7472
rect 16761 7463 16819 7469
rect 16761 7460 16773 7463
rect 15896 7432 16773 7460
rect 15896 7420 15902 7432
rect 16761 7429 16773 7432
rect 16807 7429 16819 7463
rect 20346 7460 20352 7472
rect 20307 7432 20352 7460
rect 16761 7423 16819 7429
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12176 7364 13001 7392
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 15470 7392 15476 7404
rect 15431 7364 15476 7392
rect 12989 7355 13047 7361
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7392 15715 7395
rect 15746 7392 15752 7404
rect 15703 7364 15752 7392
rect 15703 7361 15715 7364
rect 15657 7355 15715 7361
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7392 19487 7395
rect 19475 7364 19509 7392
rect 19475 7361 19487 7364
rect 19429 7355 19487 7361
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8352 7296 9045 7324
rect 8352 7284 8358 7296
rect 9033 7293 9045 7296
rect 9079 7324 9091 7327
rect 9858 7324 9864 7336
rect 9079 7296 9864 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 10652 7296 11192 7324
rect 10652 7284 10658 7296
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7256 9827 7259
rect 10106 7259 10164 7265
rect 10106 7256 10118 7259
rect 9815 7228 10118 7256
rect 9815 7225 9827 7228
rect 9769 7219 9827 7225
rect 10106 7225 10118 7228
rect 10152 7256 10164 7259
rect 11054 7256 11060 7268
rect 10152 7228 11060 7256
rect 10152 7225 10164 7228
rect 10106 7219 10164 7225
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11164 7256 11192 7296
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 12066 7324 12072 7336
rect 11296 7296 12072 7324
rect 11296 7284 11302 7296
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12894 7324 12900 7336
rect 12492 7296 12900 7324
rect 12492 7284 12498 7296
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 14550 7324 14556 7336
rect 14511 7296 14556 7324
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18012 7296 18705 7324
rect 18012 7284 18018 7296
rect 18693 7293 18705 7296
rect 18739 7324 18751 7327
rect 19242 7324 19248 7336
rect 18739 7296 19012 7324
rect 19203 7296 19248 7324
rect 18739 7293 18751 7296
rect 18693 7287 18751 7293
rect 14829 7259 14887 7265
rect 14829 7256 14841 7259
rect 11164 7228 14841 7256
rect 14829 7225 14841 7228
rect 14875 7256 14887 7259
rect 15381 7259 15439 7265
rect 15381 7256 15393 7259
rect 14875 7228 15393 7256
rect 14875 7225 14887 7228
rect 14829 7219 14887 7225
rect 15381 7225 15393 7228
rect 15427 7256 15439 7259
rect 16022 7256 16028 7268
rect 15427 7228 16028 7256
rect 15427 7225 15439 7228
rect 15381 7219 15439 7225
rect 16022 7216 16028 7228
rect 16080 7216 16086 7268
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12124 7160 12817 7188
rect 12124 7148 12130 7160
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 14366 7188 14372 7200
rect 14327 7160 14372 7188
rect 12805 7151 12863 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 15013 7191 15071 7197
rect 15013 7157 15025 7191
rect 15059 7188 15071 7191
rect 15286 7188 15292 7200
rect 15059 7160 15292 7188
rect 15059 7157 15071 7160
rect 15013 7151 15071 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 16942 7188 16948 7200
rect 16903 7160 16948 7188
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 17494 7188 17500 7200
rect 17455 7160 17500 7188
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 18325 7191 18383 7197
rect 18325 7157 18337 7191
rect 18371 7188 18383 7191
rect 18690 7188 18696 7200
rect 18371 7160 18696 7188
rect 18371 7157 18383 7160
rect 18325 7151 18383 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 18874 7188 18880 7200
rect 18835 7160 18880 7188
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 18984 7188 19012 7296
rect 19242 7284 19248 7296
rect 19300 7284 19306 7336
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19444 7324 19472 7355
rect 19889 7327 19947 7333
rect 19889 7324 19901 7327
rect 19392 7296 19901 7324
rect 19392 7284 19398 7296
rect 19889 7293 19901 7296
rect 19935 7293 19947 7327
rect 20364 7324 20392 7420
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 20990 7392 20996 7404
rect 20680 7364 20996 7392
rect 20680 7352 20686 7364
rect 20990 7352 20996 7364
rect 21048 7392 21054 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 21048 7364 21097 7392
rect 21048 7352 21054 7364
rect 21085 7361 21097 7364
rect 21131 7392 21143 7395
rect 21450 7392 21456 7404
rect 21131 7364 21456 7392
rect 21131 7361 21143 7364
rect 21085 7355 21143 7361
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 22462 7352 22468 7404
rect 22520 7392 22526 7404
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22520 7364 22661 7392
rect 22520 7352 22526 7364
rect 22649 7361 22661 7364
rect 22695 7392 22707 7395
rect 23477 7395 23535 7401
rect 22695 7364 23152 7392
rect 22695 7361 22707 7364
rect 22649 7355 22707 7361
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 20364 7296 20821 7324
rect 19889 7287 19947 7293
rect 20809 7293 20821 7296
rect 20855 7324 20867 7327
rect 21910 7324 21916 7336
rect 20855 7296 21916 7324
rect 20855 7293 20867 7296
rect 20809 7287 20867 7293
rect 21910 7284 21916 7296
rect 21968 7284 21974 7336
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22060 7296 22416 7324
rect 22060 7284 22066 7296
rect 20714 7216 20720 7268
rect 20772 7256 20778 7268
rect 20901 7259 20959 7265
rect 20901 7256 20913 7259
rect 20772 7228 20913 7256
rect 20772 7216 20778 7228
rect 20901 7225 20913 7228
rect 20947 7256 20959 7259
rect 21358 7256 21364 7268
rect 20947 7228 21364 7256
rect 20947 7225 20959 7228
rect 20901 7219 20959 7225
rect 21358 7216 21364 7228
rect 21416 7216 21422 7268
rect 22388 7200 22416 7296
rect 19337 7191 19395 7197
rect 19337 7188 19349 7191
rect 18984 7160 19349 7188
rect 19337 7157 19349 7160
rect 19383 7188 19395 7191
rect 20070 7188 20076 7200
rect 19383 7160 20076 7188
rect 19383 7157 19395 7160
rect 19337 7151 19395 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 22002 7188 22008 7200
rect 21963 7160 22008 7188
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 22370 7188 22376 7200
rect 22331 7160 22376 7188
rect 22370 7148 22376 7160
rect 22428 7148 22434 7200
rect 22465 7191 22523 7197
rect 22465 7157 22477 7191
rect 22511 7188 22523 7191
rect 22738 7188 22744 7200
rect 22511 7160 22744 7188
rect 22511 7157 22523 7160
rect 22465 7151 22523 7157
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 23124 7197 23152 7364
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 23523 7364 23796 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7293 23719 7327
rect 23768 7324 23796 7364
rect 23934 7333 23940 7336
rect 23928 7324 23940 7333
rect 23768 7296 23940 7324
rect 23661 7287 23719 7293
rect 23928 7287 23940 7296
rect 23676 7256 23704 7287
rect 23934 7284 23940 7287
rect 23992 7284 23998 7336
rect 23676 7228 23980 7256
rect 23952 7200 23980 7228
rect 23109 7191 23167 7197
rect 23109 7157 23121 7191
rect 23155 7188 23167 7191
rect 23198 7188 23204 7200
rect 23155 7160 23204 7188
rect 23155 7157 23167 7160
rect 23109 7151 23167 7157
rect 23198 7148 23204 7160
rect 23256 7148 23262 7200
rect 23934 7148 23940 7200
rect 23992 7148 23998 7200
rect 24118 7148 24124 7200
rect 24176 7188 24182 7200
rect 25041 7191 25099 7197
rect 25041 7188 25053 7191
rect 24176 7160 25053 7188
rect 24176 7148 24182 7160
rect 25041 7157 25053 7160
rect 25087 7157 25099 7191
rect 25041 7151 25099 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 11054 6984 11060 6996
rect 11015 6956 11060 6984
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 12066 6984 12072 6996
rect 12027 6956 12072 6984
rect 12066 6944 12072 6956
rect 12124 6984 12130 6996
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 12124 6956 12173 6984
rect 12124 6944 12130 6956
rect 12161 6953 12173 6956
rect 12207 6953 12219 6987
rect 12161 6947 12219 6953
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12529 6987 12587 6993
rect 12529 6984 12541 6987
rect 12308 6956 12541 6984
rect 12308 6944 12314 6956
rect 12529 6953 12541 6956
rect 12575 6984 12587 6987
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 12575 6956 13737 6984
rect 12575 6953 12587 6956
rect 12529 6947 12587 6953
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 14274 6984 14280 6996
rect 14235 6956 14280 6984
rect 13725 6947 13783 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 14550 6984 14556 6996
rect 14511 6956 14556 6984
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15470 6984 15476 6996
rect 15151 6956 15476 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 16669 6987 16727 6993
rect 16669 6984 16681 6987
rect 15804 6956 16681 6984
rect 15804 6944 15810 6956
rect 16669 6953 16681 6956
rect 16715 6953 16727 6987
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 16669 6947 16727 6953
rect 17402 6944 17408 6956
rect 17460 6984 17466 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 17460 6956 17969 6984
rect 17460 6944 17466 6956
rect 11882 6876 11888 6928
rect 11940 6916 11946 6928
rect 12621 6919 12679 6925
rect 12621 6916 12633 6919
rect 11940 6888 12633 6916
rect 11940 6876 11946 6888
rect 12621 6885 12633 6888
rect 12667 6885 12679 6919
rect 13998 6916 14004 6928
rect 12621 6879 12679 6885
rect 13832 6888 14004 6916
rect 9950 6857 9956 6860
rect 9944 6848 9956 6857
rect 9911 6820 9956 6848
rect 9944 6811 9956 6820
rect 9950 6808 9956 6811
rect 10008 6808 10014 6860
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 12710 6780 12716 6792
rect 12671 6752 12716 6780
rect 9677 6743 9735 6749
rect 9692 6644 9720 6743
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13832 6780 13860 6888
rect 13998 6876 14004 6888
rect 14056 6876 14062 6928
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 14424 6888 15148 6916
rect 14424 6876 14430 6888
rect 15120 6848 15148 6888
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 15120 6820 15301 6848
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 15378 6848 15384 6860
rect 15335 6820 15384 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15556 6851 15614 6857
rect 15556 6817 15568 6851
rect 15602 6848 15614 6851
rect 15930 6848 15936 6860
rect 15602 6820 15936 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 13495 6752 13860 6780
rect 17788 6780 17816 6956
rect 17957 6953 17969 6956
rect 18003 6953 18015 6987
rect 17957 6947 18015 6953
rect 22373 6987 22431 6993
rect 22373 6953 22385 6987
rect 22419 6984 22431 6987
rect 23198 6984 23204 6996
rect 22419 6956 23204 6984
rect 22419 6953 22431 6956
rect 22373 6947 22431 6953
rect 23198 6944 23204 6956
rect 23256 6944 23262 6996
rect 18874 6916 18880 6928
rect 18064 6888 18880 6916
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6848 17923 6851
rect 18064 6848 18092 6888
rect 18874 6876 18880 6888
rect 18932 6876 18938 6928
rect 20714 6916 20720 6928
rect 20640 6888 20720 6916
rect 17911 6820 18092 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 18196 6820 18241 6848
rect 18196 6808 18202 6820
rect 18322 6808 18328 6860
rect 18380 6848 18386 6860
rect 18489 6851 18547 6857
rect 18489 6848 18501 6851
rect 18380 6820 18501 6848
rect 18380 6808 18386 6820
rect 18489 6817 18501 6820
rect 18535 6817 18547 6851
rect 18489 6811 18547 6817
rect 20533 6851 20591 6857
rect 20533 6817 20545 6851
rect 20579 6848 20591 6851
rect 20640 6848 20668 6888
rect 20714 6876 20720 6888
rect 20772 6876 20778 6928
rect 20579 6820 20668 6848
rect 20579 6817 20591 6820
rect 20533 6811 20591 6817
rect 21082 6808 21088 6860
rect 21140 6848 21146 6860
rect 21249 6851 21307 6857
rect 21249 6848 21261 6851
rect 21140 6820 21261 6848
rect 21140 6808 21146 6820
rect 21249 6817 21261 6820
rect 21295 6817 21307 6851
rect 21249 6811 21307 6817
rect 22094 6808 22100 6860
rect 22152 6808 22158 6860
rect 23385 6851 23443 6857
rect 23385 6817 23397 6851
rect 23431 6848 23443 6851
rect 23842 6848 23848 6860
rect 23431 6820 23848 6848
rect 23431 6817 23443 6820
rect 23385 6811 23443 6817
rect 23842 6808 23848 6820
rect 23900 6808 23906 6860
rect 18230 6780 18236 6792
rect 17788 6752 18236 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20312 6752 21005 6780
rect 20312 6740 20318 6752
rect 20993 6749 21005 6752
rect 21039 6749 21051 6783
rect 22112 6780 22140 6808
rect 23290 6780 23296 6792
rect 22112 6752 23296 6780
rect 20993 6743 21051 6749
rect 23290 6740 23296 6752
rect 23348 6780 23354 6792
rect 23937 6783 23995 6789
rect 23937 6780 23949 6783
rect 23348 6752 23949 6780
rect 23348 6740 23354 6752
rect 23937 6749 23949 6752
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 24026 6740 24032 6792
rect 24084 6780 24090 6792
rect 25038 6780 25044 6792
rect 24084 6752 24129 6780
rect 24999 6752 25044 6780
rect 24084 6740 24090 6752
rect 25038 6740 25044 6752
rect 25096 6740 25102 6792
rect 22554 6672 22560 6724
rect 22612 6712 22618 6724
rect 23017 6715 23075 6721
rect 23017 6712 23029 6715
rect 22612 6684 23029 6712
rect 22612 6672 22618 6684
rect 23017 6681 23029 6684
rect 23063 6712 23075 6715
rect 23063 6684 23980 6712
rect 23063 6681 23075 6684
rect 23017 6675 23075 6681
rect 23952 6656 23980 6684
rect 9858 6644 9864 6656
rect 9692 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6644 9922 6656
rect 11146 6644 11152 6656
rect 9916 6616 11152 6644
rect 9916 6604 9922 6616
rect 11146 6604 11152 6616
rect 11204 6644 11210 6656
rect 11698 6644 11704 6656
rect 11204 6616 11704 6644
rect 11204 6604 11210 6616
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 19392 6616 19625 6644
rect 19392 6604 19398 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 23477 6647 23535 6653
rect 23477 6613 23489 6647
rect 23523 6644 23535 6647
rect 23566 6644 23572 6656
rect 23523 6616 23572 6644
rect 23523 6613 23535 6616
rect 23477 6607 23535 6613
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 23934 6604 23940 6656
rect 23992 6644 23998 6656
rect 24489 6647 24547 6653
rect 24489 6644 24501 6647
rect 23992 6616 24501 6644
rect 23992 6604 23998 6616
rect 24489 6613 24501 6616
rect 24535 6613 24547 6647
rect 24489 6607 24547 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 566 6400 572 6452
rect 624 6440 630 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 624 6412 7849 6440
rect 624 6400 630 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 10781 6443 10839 6449
rect 10781 6409 10793 6443
rect 10827 6440 10839 6443
rect 11882 6440 11888 6452
rect 10827 6412 11888 6440
rect 10827 6409 10839 6412
rect 10781 6403 10839 6409
rect 7852 6304 7880 6403
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12250 6440 12256 6452
rect 12211 6412 12256 6440
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 15930 6440 15936 6452
rect 15891 6412 15936 6440
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 17494 6440 17500 6452
rect 17455 6412 17500 6440
rect 17494 6400 17500 6412
rect 17552 6440 17558 6452
rect 18322 6440 18328 6452
rect 17552 6412 18328 6440
rect 17552 6400 17558 6412
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 21082 6440 21088 6452
rect 18708 6412 21088 6440
rect 9401 6375 9459 6381
rect 9401 6341 9413 6375
rect 9447 6341 9459 6375
rect 9401 6335 9459 6341
rect 9416 6304 9444 6335
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 12710 6372 12716 6384
rect 11112 6344 12716 6372
rect 11112 6332 11118 6344
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 9950 6304 9956 6316
rect 7852 6276 8156 6304
rect 9416 6276 9956 6304
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8128 6236 8156 6276
rect 9950 6264 9956 6276
rect 10008 6304 10014 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 10008 6276 10333 6304
rect 10008 6264 10014 6276
rect 10321 6273 10333 6276
rect 10367 6304 10379 6307
rect 11422 6304 11428 6316
rect 10367 6276 11428 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 13817 6307 13875 6313
rect 13817 6304 13829 6307
rect 12676 6276 13829 6304
rect 12676 6264 12682 6276
rect 13280 6248 13308 6276
rect 13817 6273 13829 6276
rect 13863 6273 13875 6307
rect 13998 6304 14004 6316
rect 13959 6276 14004 6304
rect 13817 6267 13875 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 15286 6264 15292 6316
rect 15344 6304 15350 6316
rect 15381 6307 15439 6313
rect 15381 6304 15393 6307
rect 15344 6276 15393 6304
rect 15344 6264 15350 6276
rect 15381 6273 15393 6276
rect 15427 6273 15439 6307
rect 15562 6304 15568 6316
rect 15523 6276 15568 6304
rect 15381 6267 15439 6273
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 18708 6313 18736 6412
rect 21082 6400 21088 6412
rect 21140 6440 21146 6452
rect 21637 6443 21695 6449
rect 21637 6440 21649 6443
rect 21140 6412 21649 6440
rect 21140 6400 21146 6412
rect 21637 6409 21649 6412
rect 21683 6409 21695 6443
rect 21637 6403 21695 6409
rect 22097 6443 22155 6449
rect 22097 6409 22109 6443
rect 22143 6440 22155 6443
rect 22186 6440 22192 6452
rect 22143 6412 22192 6440
rect 22143 6409 22155 6412
rect 22097 6403 22155 6409
rect 22186 6400 22192 6412
rect 22244 6400 22250 6452
rect 23842 6400 23848 6452
rect 23900 6440 23906 6452
rect 24397 6443 24455 6449
rect 24397 6440 24409 6443
rect 23900 6412 24409 6440
rect 23900 6400 23906 6412
rect 24397 6409 24409 6412
rect 24443 6409 24455 6443
rect 24397 6403 24455 6409
rect 23477 6375 23535 6381
rect 23477 6341 23489 6375
rect 23523 6372 23535 6375
rect 24026 6372 24032 6384
rect 23523 6344 24032 6372
rect 23523 6341 23535 6344
rect 23477 6335 23535 6341
rect 24026 6332 24032 6344
rect 24084 6332 24090 6384
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 17911 6276 18705 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18693 6273 18705 6276
rect 18739 6273 18751 6307
rect 18693 6267 18751 6273
rect 23198 6264 23204 6316
rect 23256 6304 23262 6316
rect 24578 6304 24584 6316
rect 23256 6276 24584 6304
rect 23256 6264 23262 6276
rect 24578 6264 24584 6276
rect 24636 6304 24642 6316
rect 24949 6307 25007 6313
rect 24949 6304 24961 6307
rect 24636 6276 24961 6304
rect 24636 6264 24642 6276
rect 24949 6273 24961 6276
rect 24995 6273 25007 6307
rect 24949 6267 25007 6273
rect 8277 6239 8335 6245
rect 8277 6236 8289 6239
rect 8128 6208 8289 6236
rect 8021 6199 8079 6205
rect 8277 6205 8289 6208
rect 8323 6205 8335 6239
rect 8277 6199 8335 6205
rect 8036 6100 8064 6199
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 9732 6208 10701 6236
rect 9732 6196 9738 6208
rect 10689 6205 10701 6208
rect 10735 6236 10747 6239
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 10735 6208 11161 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 11149 6205 11161 6208
rect 11195 6236 11207 6239
rect 11606 6236 11612 6248
rect 11195 6208 11612 6236
rect 11195 6205 11207 6208
rect 11149 6199 11207 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 13262 6236 13268 6248
rect 13223 6208 13268 6236
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 13722 6236 13728 6248
rect 13683 6208 13728 6236
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 18509 6239 18567 6245
rect 16899 6208 16933 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 18509 6205 18521 6239
rect 18555 6236 18567 6239
rect 18874 6236 18880 6248
rect 18555 6208 18880 6236
rect 18555 6205 18567 6208
rect 18509 6199 18567 6205
rect 10778 6128 10784 6180
rect 10836 6168 10842 6180
rect 11241 6171 11299 6177
rect 11241 6168 11253 6171
rect 10836 6140 11253 6168
rect 10836 6128 10842 6140
rect 11241 6137 11253 6140
rect 11287 6168 11299 6171
rect 11330 6168 11336 6180
rect 11287 6140 11336 6168
rect 11287 6137 11299 6140
rect 11241 6131 11299 6137
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 15289 6171 15347 6177
rect 15289 6168 15301 6171
rect 13372 6140 14044 6168
rect 8202 6100 8208 6112
rect 8036 6072 8208 6100
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 13372 6109 13400 6140
rect 14016 6112 14044 6140
rect 14752 6140 15301 6168
rect 14752 6112 14780 6140
rect 15289 6137 15301 6140
rect 15335 6137 15347 6171
rect 15289 6131 15347 6137
rect 16761 6171 16819 6177
rect 16761 6137 16773 6171
rect 16807 6168 16819 6171
rect 16868 6168 16896 6199
rect 18874 6196 18880 6208
rect 18932 6196 18938 6248
rect 19705 6239 19763 6245
rect 19705 6236 19717 6239
rect 19444 6208 19717 6236
rect 17862 6168 17868 6180
rect 16807 6140 17868 6168
rect 16807 6137 16819 6140
rect 16761 6131 16819 6137
rect 17862 6128 17868 6140
rect 17920 6128 17926 6180
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 19444 6168 19472 6208
rect 19705 6205 19717 6208
rect 19751 6236 19763 6239
rect 20254 6236 20260 6248
rect 19751 6208 20260 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22189 6239 22247 6245
rect 22189 6236 22201 6239
rect 22152 6208 22201 6236
rect 22152 6196 22158 6208
rect 22189 6205 22201 6208
rect 22235 6236 22247 6239
rect 22741 6239 22799 6245
rect 22741 6236 22753 6239
rect 22235 6208 22753 6236
rect 22235 6205 22247 6208
rect 22189 6199 22247 6205
rect 22741 6205 22753 6208
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 24305 6239 24363 6245
rect 24305 6205 24317 6239
rect 24351 6236 24363 6239
rect 24762 6236 24768 6248
rect 24351 6208 24768 6236
rect 24351 6205 24363 6208
rect 24305 6199 24363 6205
rect 24762 6196 24768 6208
rect 24820 6236 24826 6248
rect 24857 6239 24915 6245
rect 24857 6236 24869 6239
rect 24820 6208 24869 6236
rect 24820 6196 24826 6208
rect 24857 6205 24869 6208
rect 24903 6205 24915 6239
rect 24857 6199 24915 6205
rect 19950 6171 20008 6177
rect 19950 6168 19962 6171
rect 18288 6140 19472 6168
rect 19536 6140 19962 6168
rect 18288 6128 18294 6140
rect 13357 6103 13415 6109
rect 13357 6069 13369 6103
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 14056 6072 14381 6100
rect 14056 6060 14062 6072
rect 14369 6069 14381 6072
rect 14415 6069 14427 6103
rect 14734 6100 14740 6112
rect 14695 6072 14740 6100
rect 14369 6063 14427 6069
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 15378 6100 15384 6112
rect 14967 6072 15384 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15746 6100 15752 6112
rect 15528 6072 15752 6100
rect 15528 6060 15534 6072
rect 15746 6060 15752 6072
rect 15804 6100 15810 6112
rect 16301 6103 16359 6109
rect 16301 6100 16313 6103
rect 15804 6072 16313 6100
rect 15804 6060 15810 6072
rect 16301 6069 16313 6072
rect 16347 6069 16359 6103
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 16301 6063 16359 6069
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 18138 6100 18144 6112
rect 18099 6072 18144 6100
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 18598 6060 18604 6072
rect 18656 6100 18662 6112
rect 19153 6103 19211 6109
rect 19153 6100 19165 6103
rect 18656 6072 19165 6100
rect 18656 6060 18662 6072
rect 19153 6069 19165 6072
rect 19199 6069 19211 6103
rect 19153 6063 19211 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19536 6109 19564 6140
rect 19950 6137 19962 6140
rect 19996 6137 20008 6171
rect 19950 6131 20008 6137
rect 19521 6103 19579 6109
rect 19521 6100 19533 6103
rect 19392 6072 19533 6100
rect 19392 6060 19398 6072
rect 19521 6069 19533 6072
rect 19567 6069 19579 6103
rect 19521 6063 19579 6069
rect 22373 6103 22431 6109
rect 22373 6069 22385 6103
rect 22419 6100 22431 6103
rect 23382 6100 23388 6112
rect 22419 6072 23388 6100
rect 22419 6069 22431 6072
rect 22373 6063 22431 6069
rect 23382 6060 23388 6072
rect 23440 6060 23446 6112
rect 23937 6103 23995 6109
rect 23937 6069 23949 6103
rect 23983 6100 23995 6103
rect 24765 6103 24823 6109
rect 24765 6100 24777 6103
rect 23983 6072 24777 6100
rect 23983 6069 23995 6072
rect 23937 6063 23995 6069
rect 24765 6069 24777 6072
rect 24811 6100 24823 6103
rect 24854 6100 24860 6112
rect 24811 6072 24860 6100
rect 24811 6069 24823 6072
rect 24765 6063 24823 6069
rect 24854 6060 24860 6072
rect 24912 6060 24918 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 8113 5899 8171 5905
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 8202 5896 8208 5908
rect 8159 5868 8208 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 9950 5896 9956 5908
rect 9911 5868 9956 5896
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 11701 5899 11759 5905
rect 11701 5865 11713 5899
rect 11747 5896 11759 5899
rect 12342 5896 12348 5908
rect 11747 5868 12348 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13449 5899 13507 5905
rect 13449 5865 13461 5899
rect 13495 5896 13507 5899
rect 13722 5896 13728 5908
rect 13495 5868 13728 5896
rect 13495 5865 13507 5868
rect 13449 5859 13507 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 13998 5896 14004 5908
rect 13959 5868 14004 5896
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 15286 5856 15292 5908
rect 15344 5896 15350 5908
rect 15473 5899 15531 5905
rect 15473 5896 15485 5899
rect 15344 5868 15485 5896
rect 15344 5856 15350 5868
rect 15473 5865 15485 5868
rect 15519 5865 15531 5899
rect 15473 5859 15531 5865
rect 17129 5899 17187 5905
rect 17129 5865 17141 5899
rect 17175 5865 17187 5899
rect 17129 5859 17187 5865
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 18046 5896 18052 5908
rect 17819 5868 18052 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 16482 5788 16488 5840
rect 16540 5828 16546 5840
rect 17144 5828 17172 5859
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18322 5896 18328 5908
rect 18187 5868 18328 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18322 5856 18328 5868
rect 18380 5896 18386 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 18380 5868 19625 5896
rect 18380 5856 18386 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 20254 5896 20260 5908
rect 20215 5868 20260 5896
rect 19613 5859 19671 5865
rect 20254 5856 20260 5868
rect 20312 5896 20318 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 20312 5868 20637 5896
rect 20312 5856 20318 5868
rect 20625 5865 20637 5868
rect 20671 5865 20683 5899
rect 20625 5859 20683 5865
rect 18414 5828 18420 5840
rect 16540 5800 18420 5828
rect 16540 5788 16546 5800
rect 18414 5788 18420 5800
rect 18472 5837 18478 5840
rect 18472 5831 18536 5837
rect 18472 5797 18490 5831
rect 18524 5797 18536 5831
rect 18472 5791 18536 5797
rect 18472 5788 18478 5791
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 11698 5760 11704 5772
rect 10367 5732 11704 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 12066 5760 12072 5772
rect 12027 5732 12072 5760
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 16005 5763 16063 5769
rect 16005 5760 16017 5763
rect 15580 5732 16017 5760
rect 10778 5692 10784 5704
rect 10739 5664 10784 5692
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 12158 5692 12164 5704
rect 12119 5664 12164 5692
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5692 12403 5695
rect 12710 5692 12716 5704
rect 12391 5664 12716 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 14090 5692 14096 5704
rect 14051 5664 14096 5692
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14185 5695 14243 5701
rect 14185 5661 14197 5695
rect 14231 5661 14243 5695
rect 14185 5655 14243 5661
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 14200 5624 14228 5655
rect 15580 5636 15608 5732
rect 16005 5729 16017 5732
rect 16051 5729 16063 5763
rect 18230 5760 18236 5772
rect 18191 5732 18236 5760
rect 16005 5723 16063 5729
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 20640 5760 20668 5859
rect 21450 5856 21456 5908
rect 21508 5896 21514 5908
rect 22373 5899 22431 5905
rect 22373 5896 22385 5899
rect 21508 5868 22385 5896
rect 21508 5856 21514 5868
rect 22373 5865 22385 5868
rect 22419 5865 22431 5899
rect 22373 5859 22431 5865
rect 23017 5899 23075 5905
rect 23017 5865 23029 5899
rect 23063 5896 23075 5899
rect 23750 5896 23756 5908
rect 23063 5868 23756 5896
rect 23063 5865 23075 5868
rect 23017 5859 23075 5865
rect 23750 5856 23756 5868
rect 23808 5896 23814 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 23808 5868 23857 5896
rect 23808 5856 23814 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 24578 5896 24584 5908
rect 24539 5868 24584 5896
rect 23845 5859 23903 5865
rect 24578 5856 24584 5868
rect 24636 5856 24642 5908
rect 21174 5788 21180 5840
rect 21232 5837 21238 5840
rect 21232 5831 21296 5837
rect 21232 5797 21250 5831
rect 21284 5797 21296 5831
rect 23290 5828 23296 5840
rect 23251 5800 23296 5828
rect 21232 5791 21296 5797
rect 21232 5788 21238 5791
rect 23290 5788 23296 5800
rect 23348 5788 23354 5840
rect 23474 5788 23480 5840
rect 23532 5828 23538 5840
rect 23934 5828 23940 5840
rect 23532 5800 23940 5828
rect 23532 5788 23538 5800
rect 23934 5788 23940 5800
rect 23992 5788 23998 5840
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20640 5732 21005 5760
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 25041 5763 25099 5769
rect 25041 5729 25053 5763
rect 25087 5760 25099 5763
rect 25590 5760 25596 5772
rect 25087 5732 25596 5760
rect 25087 5729 25099 5732
rect 25041 5723 25099 5729
rect 25590 5720 25596 5732
rect 25648 5720 25654 5772
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 23566 5652 23572 5704
rect 23624 5692 23630 5704
rect 23937 5695 23995 5701
rect 23937 5692 23949 5695
rect 23624 5664 23949 5692
rect 23624 5652 23630 5664
rect 23937 5661 23949 5664
rect 23983 5661 23995 5695
rect 23937 5655 23995 5661
rect 24026 5652 24032 5704
rect 24084 5692 24090 5704
rect 24084 5664 24129 5692
rect 24084 5652 24090 5664
rect 14921 5627 14979 5633
rect 14921 5624 14933 5627
rect 13872 5596 14933 5624
rect 13872 5584 13878 5596
rect 14921 5593 14933 5596
rect 14967 5624 14979 5627
rect 15562 5624 15568 5636
rect 14967 5596 15568 5624
rect 14967 5593 14979 5596
rect 14921 5587 14979 5593
rect 15562 5584 15568 5596
rect 15620 5584 15626 5636
rect 13633 5559 13691 5565
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 13906 5556 13912 5568
rect 13679 5528 13912 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 23474 5556 23480 5568
rect 23435 5528 23480 5556
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 23842 5516 23848 5568
rect 23900 5556 23906 5568
rect 24857 5559 24915 5565
rect 24857 5556 24869 5559
rect 23900 5528 24869 5556
rect 23900 5516 23906 5528
rect 24857 5525 24869 5528
rect 24903 5525 24915 5559
rect 24857 5519 24915 5525
rect 25225 5559 25283 5565
rect 25225 5525 25237 5559
rect 25271 5556 25283 5559
rect 26142 5556 26148 5568
rect 25271 5528 26148 5556
rect 25271 5525 25283 5528
rect 25225 5519 25283 5525
rect 26142 5516 26148 5528
rect 26200 5516 26206 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 11241 5355 11299 5361
rect 11241 5321 11253 5355
rect 11287 5352 11299 5355
rect 12158 5352 12164 5364
rect 11287 5324 12164 5352
rect 11287 5321 11299 5324
rect 11241 5315 11299 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 13722 5352 13728 5364
rect 13683 5324 13728 5352
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 13998 5352 14004 5364
rect 13959 5324 14004 5352
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 15562 5352 15568 5364
rect 15523 5324 15568 5352
rect 15562 5312 15568 5324
rect 15620 5352 15626 5364
rect 16117 5355 16175 5361
rect 16117 5352 16129 5355
rect 15620 5324 16129 5352
rect 15620 5312 15626 5324
rect 16117 5321 16129 5324
rect 16163 5321 16175 5355
rect 16117 5315 16175 5321
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23566 5352 23572 5364
rect 23155 5324 23572 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23566 5312 23572 5324
rect 23624 5312 23630 5364
rect 24026 5352 24032 5364
rect 23860 5324 24032 5352
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12621 5287 12679 5293
rect 12621 5284 12633 5287
rect 12124 5256 12633 5284
rect 12124 5244 12130 5256
rect 12621 5253 12633 5256
rect 12667 5253 12679 5287
rect 12621 5247 12679 5253
rect 11330 5216 11336 5228
rect 11291 5188 11336 5216
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 12802 5176 12808 5228
rect 12860 5216 12866 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 12860 5188 13093 5216
rect 12860 5176 12866 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5216 13323 5219
rect 13354 5216 13360 5228
rect 13311 5188 13360 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12529 5151 12587 5157
rect 12529 5148 12541 5151
rect 12299 5120 12541 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12529 5117 12541 5120
rect 12575 5117 12587 5151
rect 12529 5111 12587 5117
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 11885 5083 11943 5089
rect 11885 5080 11897 5083
rect 11480 5052 11897 5080
rect 11480 5040 11486 5052
rect 11885 5049 11897 5052
rect 11931 5080 11943 5083
rect 13280 5080 13308 5179
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14016 5216 14044 5312
rect 23477 5287 23535 5293
rect 23477 5253 23489 5287
rect 23523 5284 23535 5287
rect 23860 5284 23888 5324
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 25590 5312 25596 5364
rect 25648 5352 25654 5364
rect 25777 5355 25835 5361
rect 25777 5352 25789 5355
rect 25648 5324 25789 5352
rect 25648 5312 25654 5324
rect 25777 5321 25789 5324
rect 25823 5321 25835 5355
rect 25777 5315 25835 5321
rect 23523 5256 23888 5284
rect 23523 5253 23535 5256
rect 23477 5247 23535 5253
rect 14016 5188 14320 5216
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5117 14243 5151
rect 14292 5148 14320 5188
rect 18322 5176 18328 5228
rect 18380 5216 18386 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18380 5188 18797 5216
rect 18380 5176 18386 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 19610 5216 19616 5228
rect 19571 5188 19616 5216
rect 18785 5179 18843 5185
rect 19610 5176 19616 5188
rect 19668 5216 19674 5228
rect 20346 5216 20352 5228
rect 19668 5188 20208 5216
rect 20307 5188 20352 5216
rect 19668 5176 19674 5188
rect 14441 5151 14499 5157
rect 14441 5148 14453 5151
rect 14292 5120 14453 5148
rect 14185 5111 14243 5117
rect 14441 5117 14453 5120
rect 14487 5148 14499 5151
rect 14826 5148 14832 5160
rect 14487 5120 14832 5148
rect 14487 5117 14499 5120
rect 14441 5111 14499 5117
rect 11931 5052 13308 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12529 5015 12587 5021
rect 12529 4981 12541 5015
rect 12575 5012 12587 5015
rect 12989 5015 13047 5021
rect 12989 5012 13001 5015
rect 12575 4984 13001 5012
rect 12575 4981 12587 4984
rect 12529 4975 12587 4981
rect 12989 4981 13001 4984
rect 13035 5012 13047 5015
rect 13262 5012 13268 5024
rect 13035 4984 13268 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 14200 5012 14228 5111
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 16850 5108 16856 5120
rect 16908 5148 16914 5160
rect 20180 5157 20208 5188
rect 20346 5176 20352 5188
rect 20404 5176 20410 5228
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21174 5216 21180 5228
rect 21131 5188 21180 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 21174 5176 21180 5188
rect 21232 5216 21238 5228
rect 23566 5216 23572 5228
rect 21232 5188 23572 5216
rect 21232 5176 21238 5188
rect 23566 5176 23572 5188
rect 23624 5176 23630 5228
rect 17405 5151 17463 5157
rect 17405 5148 17417 5151
rect 16908 5120 17417 5148
rect 16908 5108 16914 5120
rect 17405 5117 17417 5120
rect 17451 5117 17463 5151
rect 17405 5111 17463 5117
rect 20165 5151 20223 5157
rect 20165 5117 20177 5151
rect 20211 5117 20223 5151
rect 21358 5148 21364 5160
rect 21271 5120 21364 5148
rect 20165 5111 20223 5117
rect 21358 5108 21364 5120
rect 21416 5148 21422 5160
rect 21913 5151 21971 5157
rect 21913 5148 21925 5151
rect 21416 5120 21925 5148
rect 21416 5108 21422 5120
rect 21913 5117 21925 5120
rect 21959 5117 21971 5151
rect 21913 5111 21971 5117
rect 22465 5151 22523 5157
rect 22465 5117 22477 5151
rect 22511 5148 22523 5151
rect 23842 5148 23848 5160
rect 22511 5120 22545 5148
rect 23803 5120 23848 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 17865 5083 17923 5089
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 18601 5083 18659 5089
rect 18601 5080 18613 5083
rect 17911 5052 18613 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18601 5049 18613 5052
rect 18647 5080 18659 5083
rect 18782 5080 18788 5092
rect 18647 5052 18788 5080
rect 18647 5049 18659 5052
rect 18601 5043 18659 5049
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 22373 5083 22431 5089
rect 22373 5049 22385 5083
rect 22419 5080 22431 5083
rect 22480 5080 22508 5111
rect 23842 5108 23848 5120
rect 23900 5108 23906 5160
rect 23198 5080 23204 5092
rect 22419 5052 23204 5080
rect 22419 5049 22431 5052
rect 22373 5043 22431 5049
rect 23198 5040 23204 5052
rect 23256 5040 23262 5092
rect 24118 5089 24124 5092
rect 24112 5080 24124 5089
rect 24079 5052 24124 5080
rect 24112 5043 24124 5052
rect 24118 5040 24124 5043
rect 24176 5040 24182 5092
rect 15746 5012 15752 5024
rect 14200 4984 15752 5012
rect 15746 4972 15752 4984
rect 15804 5012 15810 5024
rect 16577 5015 16635 5021
rect 16577 5012 16589 5015
rect 15804 4984 16589 5012
rect 15804 4972 15810 4984
rect 16577 4981 16589 4984
rect 16623 5012 16635 5015
rect 16758 5012 16764 5024
rect 16623 4984 16764 5012
rect 16623 4981 16635 4984
rect 16577 4975 16635 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 17034 5012 17040 5024
rect 16995 4984 17040 5012
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 18690 5012 18696 5024
rect 18651 4984 18696 5012
rect 18690 4972 18696 4984
rect 18748 5012 18754 5024
rect 19245 5015 19303 5021
rect 19245 5012 19257 5015
rect 18748 4984 19257 5012
rect 18748 4972 18754 4984
rect 19245 4981 19257 4984
rect 19291 4981 19303 5015
rect 19245 4975 19303 4981
rect 19797 5015 19855 5021
rect 19797 4981 19809 5015
rect 19843 5012 19855 5015
rect 19978 5012 19984 5024
rect 19843 4984 19984 5012
rect 19843 4981 19855 4984
rect 19797 4975 19855 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20254 5012 20260 5024
rect 20215 4984 20260 5012
rect 20254 4972 20260 4984
rect 20312 4972 20318 5024
rect 21542 5012 21548 5024
rect 21503 4984 21548 5012
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 22646 5012 22652 5024
rect 22607 4984 22652 5012
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 24854 4972 24860 5024
rect 24912 5012 24918 5024
rect 25225 5015 25283 5021
rect 25225 5012 25237 5015
rect 24912 4984 25237 5012
rect 24912 4972 24918 4984
rect 25225 4981 25237 4984
rect 25271 4981 25283 5015
rect 25225 4975 25283 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 12066 4808 12072 4820
rect 12027 4780 12072 4808
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 12437 4811 12495 4817
rect 12437 4808 12449 4811
rect 12216 4780 12449 4808
rect 12216 4768 12222 4780
rect 12437 4777 12449 4780
rect 12483 4777 12495 4811
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 12437 4771 12495 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 14090 4808 14096 4820
rect 14047 4780 14096 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 14826 4808 14832 4820
rect 14787 4780 14832 4808
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15436 4780 15669 4808
rect 15436 4768 15442 4780
rect 15657 4777 15669 4780
rect 15703 4808 15715 4811
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 15703 4780 16313 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 16301 4771 16359 4777
rect 18325 4811 18383 4817
rect 18325 4777 18337 4811
rect 18371 4808 18383 4811
rect 18598 4808 18604 4820
rect 18371 4780 18604 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 19889 4811 19947 4817
rect 19889 4777 19901 4811
rect 19935 4808 19947 4811
rect 20254 4808 20260 4820
rect 19935 4780 20260 4808
rect 19935 4777 19947 4780
rect 19889 4771 19947 4777
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 23017 4811 23075 4817
rect 23017 4777 23029 4811
rect 23063 4808 23075 4811
rect 23106 4808 23112 4820
rect 23063 4780 23112 4808
rect 23063 4777 23075 4780
rect 23017 4771 23075 4777
rect 23106 4768 23112 4780
rect 23164 4768 23170 4820
rect 23290 4768 23296 4820
rect 23348 4808 23354 4820
rect 23385 4811 23443 4817
rect 23385 4808 23397 4811
rect 23348 4780 23397 4808
rect 23348 4768 23354 4780
rect 23385 4777 23397 4780
rect 23431 4777 23443 4811
rect 23385 4771 23443 4777
rect 24581 4811 24639 4817
rect 24581 4777 24593 4811
rect 24627 4808 24639 4811
rect 24670 4808 24676 4820
rect 24627 4780 24676 4808
rect 24627 4777 24639 4780
rect 24581 4771 24639 4777
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 24762 4768 24768 4820
rect 24820 4808 24826 4820
rect 25038 4808 25044 4820
rect 24820 4780 25044 4808
rect 24820 4768 24826 4780
rect 25038 4768 25044 4780
rect 25096 4768 25102 4820
rect 11793 4743 11851 4749
rect 11793 4709 11805 4743
rect 11839 4740 11851 4743
rect 12710 4740 12716 4752
rect 11839 4712 12716 4740
rect 11839 4709 11851 4712
rect 11793 4703 11851 4709
rect 12710 4700 12716 4712
rect 12768 4700 12774 4752
rect 12802 4700 12808 4752
rect 12860 4740 12866 4752
rect 16390 4740 16396 4752
rect 12860 4712 16396 4740
rect 12860 4700 12866 4712
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 18233 4743 18291 4749
rect 18233 4709 18245 4743
rect 18279 4740 18291 4743
rect 18414 4740 18420 4752
rect 18279 4712 18420 4740
rect 18279 4709 18291 4712
rect 18233 4703 18291 4709
rect 18414 4700 18420 4712
rect 18472 4700 18478 4752
rect 18506 4700 18512 4752
rect 18564 4740 18570 4752
rect 18693 4743 18751 4749
rect 18693 4740 18705 4743
rect 18564 4712 18705 4740
rect 18564 4700 18570 4712
rect 18693 4709 18705 4712
rect 18739 4709 18751 4743
rect 18693 4703 18751 4709
rect 19429 4743 19487 4749
rect 19429 4709 19441 4743
rect 19475 4740 19487 4743
rect 20162 4740 20168 4752
rect 19475 4712 20168 4740
rect 19475 4709 19487 4712
rect 19429 4703 19487 4709
rect 20162 4700 20168 4712
rect 20220 4740 20226 4752
rect 20533 4743 20591 4749
rect 20533 4740 20545 4743
rect 20220 4712 20545 4740
rect 20220 4700 20226 4712
rect 20533 4709 20545 4712
rect 20579 4740 20591 4743
rect 21361 4743 21419 4749
rect 21361 4740 21373 4743
rect 20579 4712 21373 4740
rect 20579 4709 20591 4712
rect 20533 4703 20591 4709
rect 21361 4709 21373 4712
rect 21407 4740 21419 4743
rect 23842 4740 23848 4752
rect 21407 4712 23848 4740
rect 21407 4709 21419 4712
rect 21361 4703 21419 4709
rect 23842 4700 23848 4712
rect 23900 4740 23906 4752
rect 24397 4743 24455 4749
rect 24397 4740 24409 4743
rect 23900 4712 24409 4740
rect 23900 4700 23906 4712
rect 24397 4709 24409 4712
rect 24443 4709 24455 4743
rect 24946 4740 24952 4752
rect 24907 4712 24952 4740
rect 24397 4703 24455 4709
rect 24946 4700 24952 4712
rect 25004 4700 25010 4752
rect 14093 4675 14151 4681
rect 14093 4641 14105 4675
rect 14139 4672 14151 4675
rect 14458 4672 14464 4684
rect 14139 4644 14464 4672
rect 14139 4641 14151 4644
rect 14093 4635 14151 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 15286 4632 15292 4684
rect 15344 4672 15350 4684
rect 15749 4675 15807 4681
rect 15749 4672 15761 4675
rect 15344 4644 15761 4672
rect 15344 4632 15350 4644
rect 15749 4641 15761 4644
rect 15795 4641 15807 4675
rect 15749 4635 15807 4641
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 21913 4675 21971 4681
rect 21913 4641 21925 4675
rect 21959 4672 21971 4675
rect 22002 4672 22008 4684
rect 21959 4644 22008 4672
rect 21959 4641 21971 4644
rect 21913 4635 21971 4641
rect 12894 4604 12900 4616
rect 12855 4576 12900 4604
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13354 4604 13360 4616
rect 13127 4576 13360 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 15930 4604 15936 4616
rect 15843 4576 15936 4604
rect 15930 4564 15936 4576
rect 15988 4604 15994 4616
rect 16482 4604 16488 4616
rect 15988 4576 16488 4604
rect 15988 4564 15994 4576
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 14274 4536 14280 4548
rect 14235 4508 14280 4536
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 15289 4539 15347 4545
rect 15289 4505 15301 4539
rect 15335 4536 15347 4539
rect 16868 4536 16896 4635
rect 22002 4632 22008 4644
rect 22060 4632 22066 4684
rect 17034 4604 17040 4616
rect 16995 4576 17040 4604
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 18230 4564 18236 4616
rect 18288 4604 18294 4616
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 18288 4576 18797 4604
rect 18288 4564 18294 4576
rect 18785 4573 18797 4576
rect 18831 4573 18843 4607
rect 18966 4604 18972 4616
rect 18927 4576 18972 4604
rect 18785 4567 18843 4573
rect 18966 4564 18972 4576
rect 19024 4604 19030 4616
rect 19242 4604 19248 4616
rect 19024 4576 19248 4604
rect 19024 4564 19030 4576
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 20901 4607 20959 4613
rect 20901 4573 20913 4607
rect 20947 4604 20959 4607
rect 21450 4604 21456 4616
rect 20947 4576 21456 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 21450 4564 21456 4576
rect 21508 4564 21514 4616
rect 23106 4564 23112 4616
rect 23164 4604 23170 4616
rect 23477 4607 23535 4613
rect 23477 4604 23489 4607
rect 23164 4576 23489 4604
rect 23164 4564 23170 4576
rect 23477 4573 23489 4576
rect 23523 4573 23535 4607
rect 23477 4567 23535 4573
rect 23566 4564 23572 4616
rect 23624 4604 23630 4616
rect 23661 4607 23719 4613
rect 23661 4604 23673 4607
rect 23624 4576 23673 4604
rect 23624 4564 23630 4576
rect 23661 4573 23673 4576
rect 23707 4604 23719 4607
rect 24854 4604 24860 4616
rect 23707 4576 24860 4604
rect 23707 4573 23719 4576
rect 23661 4567 23719 4573
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 25130 4564 25136 4616
rect 25188 4604 25194 4616
rect 25188 4576 25233 4604
rect 25188 4564 25194 4576
rect 17589 4539 17647 4545
rect 17589 4536 17601 4539
rect 15335 4508 17601 4536
rect 15335 4505 15347 4508
rect 15289 4499 15347 4505
rect 17589 4505 17601 4508
rect 17635 4505 17647 4539
rect 17589 4499 17647 4505
rect 16758 4468 16764 4480
rect 16719 4440 16764 4468
rect 16758 4428 16764 4440
rect 16816 4428 16822 4480
rect 19518 4428 19524 4480
rect 19576 4468 19582 4480
rect 20165 4471 20223 4477
rect 20165 4468 20177 4471
rect 19576 4440 20177 4468
rect 19576 4428 19582 4440
rect 20165 4437 20177 4440
rect 20211 4468 20223 4471
rect 20346 4468 20352 4480
rect 20211 4440 20352 4468
rect 20211 4437 20223 4440
rect 20165 4431 20223 4437
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22554 4468 22560 4480
rect 22152 4440 22197 4468
rect 22515 4440 22560 4468
rect 22152 4428 22158 4440
rect 22554 4428 22560 4440
rect 22612 4428 22618 4480
rect 22830 4468 22836 4480
rect 22791 4440 22836 4468
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 24118 4468 24124 4480
rect 24079 4440 24124 4468
rect 24118 4428 24124 4440
rect 24176 4428 24182 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 12989 4267 13047 4273
rect 12989 4264 13001 4267
rect 12860 4236 13001 4264
rect 12860 4224 12866 4236
rect 12989 4233 13001 4236
rect 13035 4233 13047 4267
rect 13354 4264 13360 4276
rect 13315 4236 13360 4264
rect 12989 4227 13047 4233
rect 13354 4224 13360 4236
rect 13412 4224 13418 4276
rect 14090 4224 14096 4276
rect 14148 4264 14154 4276
rect 14829 4267 14887 4273
rect 14829 4264 14841 4267
rect 14148 4236 14841 4264
rect 14148 4224 14154 4236
rect 14829 4233 14841 4236
rect 14875 4233 14887 4267
rect 15930 4264 15936 4276
rect 15891 4236 15936 4264
rect 14829 4227 14887 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 17865 4267 17923 4273
rect 17865 4233 17877 4267
rect 17911 4264 17923 4267
rect 18230 4264 18236 4276
rect 17911 4236 18236 4264
rect 17911 4233 17923 4236
rect 17865 4227 17923 4233
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 18966 4264 18972 4276
rect 18927 4236 18972 4264
rect 18966 4224 18972 4236
rect 19024 4224 19030 4276
rect 21450 4264 21456 4276
rect 21411 4236 21456 4264
rect 21450 4224 21456 4236
rect 21508 4224 21514 4276
rect 21913 4267 21971 4273
rect 21913 4233 21925 4267
rect 21959 4264 21971 4267
rect 22002 4264 22008 4276
rect 21959 4236 22008 4264
rect 21959 4233 21971 4236
rect 21913 4227 21971 4233
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 23109 4267 23167 4273
rect 23109 4233 23121 4267
rect 23155 4264 23167 4267
rect 23290 4264 23296 4276
rect 23155 4236 23296 4264
rect 23155 4233 23167 4236
rect 23109 4227 23167 4233
rect 23290 4224 23296 4236
rect 23348 4224 23354 4276
rect 24946 4224 24952 4276
rect 25004 4264 25010 4276
rect 25593 4267 25651 4273
rect 25593 4264 25605 4267
rect 25004 4236 25605 4264
rect 25004 4224 25010 4236
rect 25593 4233 25605 4236
rect 25639 4233 25651 4267
rect 25593 4227 25651 4233
rect 934 4156 940 4208
rect 992 4196 998 4208
rect 9582 4196 9588 4208
rect 992 4168 9588 4196
rect 992 4156 998 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 11885 4199 11943 4205
rect 11885 4165 11897 4199
rect 11931 4196 11943 4199
rect 12894 4196 12900 4208
rect 11931 4168 12900 4196
rect 11931 4165 11943 4168
rect 11885 4159 11943 4165
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 14369 4199 14427 4205
rect 14369 4165 14381 4199
rect 14415 4196 14427 4199
rect 14458 4196 14464 4208
rect 14415 4168 14464 4196
rect 14415 4165 14427 4168
rect 14369 4159 14427 4165
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 14918 4156 14924 4208
rect 14976 4196 14982 4208
rect 14976 4168 15424 4196
rect 14976 4156 14982 4168
rect 14476 4128 14504 4156
rect 15396 4137 15424 4168
rect 15289 4131 15347 4137
rect 15289 4128 15301 4131
rect 14476 4100 15301 4128
rect 15289 4097 15301 4100
rect 15335 4097 15347 4131
rect 15289 4091 15347 4097
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4097 15439 4131
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 15381 4091 15439 4097
rect 16298 4088 16304 4100
rect 16356 4128 16362 4140
rect 16356 4100 16436 4128
rect 16356 4088 16362 4100
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 9582 4060 9588 4072
rect 9180 4032 9588 4060
rect 9180 4020 9186 4032
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 11164 4032 11253 4060
rect 11164 3936 11192 4032
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11388 4032 12173 4060
rect 11388 4020 11394 4032
rect 12161 4029 12173 4032
rect 12207 4060 12219 4063
rect 12434 4060 12440 4072
rect 12207 4032 12440 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 12434 4020 12440 4032
rect 12492 4060 12498 4072
rect 13541 4063 13599 4069
rect 12492 4032 12537 4060
rect 12492 4020 12498 4032
rect 13541 4029 13553 4063
rect 13587 4060 13599 4063
rect 13630 4060 13636 4072
rect 13587 4032 13636 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 16408 4069 16436 4100
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17920 4100 18337 4128
rect 17920 4088 17926 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 22554 4128 22560 4140
rect 22515 4100 22560 4128
rect 18325 4091 18383 4097
rect 22554 4088 22560 4100
rect 22612 4088 22618 4140
rect 23477 4131 23535 4137
rect 23477 4097 23489 4131
rect 23523 4128 23535 4131
rect 23566 4128 23572 4140
rect 23523 4100 23572 4128
rect 23523 4097 23535 4100
rect 23477 4091 23535 4097
rect 23566 4088 23572 4100
rect 23624 4088 23630 4140
rect 16393 4063 16451 4069
rect 16393 4029 16405 4063
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4060 17555 4063
rect 18138 4060 18144 4072
rect 17543 4032 18144 4060
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 19429 4063 19487 4069
rect 19429 4029 19441 4063
rect 19475 4060 19487 4063
rect 20162 4060 20168 4072
rect 19475 4032 20168 4060
rect 19475 4029 19487 4032
rect 19429 4023 19487 4029
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 21450 4020 21456 4072
rect 21508 4060 21514 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 21508 4032 22385 4060
rect 21508 4020 21514 4032
rect 22373 4029 22385 4032
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22830 4060 22836 4072
rect 22511 4032 22836 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 13814 3992 13820 4004
rect 13775 3964 13820 3992
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 16666 3992 16672 4004
rect 16627 3964 16672 3992
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 19674 3995 19732 4001
rect 19674 3992 19686 3995
rect 19536 3964 19686 3992
rect 19536 3936 19564 3964
rect 19674 3961 19686 3964
rect 19720 3961 19732 3995
rect 19674 3955 19732 3961
rect 22094 3952 22100 4004
rect 22152 3992 22158 4004
rect 22480 3992 22508 4023
rect 22830 4020 22836 4032
rect 22888 4020 22894 4072
rect 23661 4063 23719 4069
rect 23661 4029 23673 4063
rect 23707 4060 23719 4063
rect 23750 4060 23756 4072
rect 23707 4032 23756 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 22152 3964 22508 3992
rect 22152 3952 22158 3964
rect 23842 3952 23848 4004
rect 23900 4001 23906 4004
rect 23900 3995 23964 4001
rect 23900 3961 23918 3995
rect 23952 3961 23964 3995
rect 23900 3955 23964 3961
rect 23900 3952 23906 3955
rect 11146 3924 11152 3936
rect 11107 3896 11152 3924
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12618 3924 12624 3936
rect 12579 3896 12624 3924
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 15194 3924 15200 3936
rect 14783 3896 15200 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 19337 3927 19395 3933
rect 19337 3893 19349 3927
rect 19383 3924 19395 3927
rect 19518 3924 19524 3936
rect 19383 3896 19524 3924
rect 19383 3893 19395 3896
rect 19337 3887 19395 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 20809 3927 20867 3933
rect 20809 3924 20821 3927
rect 20772 3896 20821 3924
rect 20772 3884 20778 3896
rect 20809 3893 20821 3896
rect 20855 3893 20867 3927
rect 20809 3887 20867 3893
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22005 3927 22063 3933
rect 22005 3924 22017 3927
rect 21968 3896 22017 3924
rect 21968 3884 21974 3896
rect 22005 3893 22017 3896
rect 22051 3893 22063 3927
rect 22005 3887 22063 3893
rect 22922 3884 22928 3936
rect 22980 3924 22986 3936
rect 23750 3924 23756 3936
rect 22980 3896 23756 3924
rect 22980 3884 22986 3896
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 25038 3924 25044 3936
rect 24999 3896 25044 3924
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 11514 3720 11520 3732
rect 11379 3692 11520 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13357 3723 13415 3729
rect 13357 3689 13369 3723
rect 13403 3720 13415 3723
rect 13538 3720 13544 3732
rect 13403 3692 13544 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14461 3723 14519 3729
rect 14461 3720 14473 3723
rect 13964 3692 14473 3720
rect 13964 3680 13970 3692
rect 14461 3689 14473 3692
rect 14507 3720 14519 3723
rect 15102 3720 15108 3732
rect 14507 3692 15108 3720
rect 14507 3689 14519 3692
rect 14461 3683 14519 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 16114 3720 16120 3732
rect 16075 3692 16120 3720
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 18693 3723 18751 3729
rect 18693 3720 18705 3723
rect 18564 3692 18705 3720
rect 18564 3680 18570 3692
rect 18693 3689 18705 3692
rect 18739 3689 18751 3723
rect 19242 3720 19248 3732
rect 19203 3692 19248 3720
rect 18693 3683 18751 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19613 3723 19671 3729
rect 19613 3720 19625 3723
rect 19484 3692 19625 3720
rect 19484 3680 19490 3692
rect 19613 3689 19625 3692
rect 19659 3689 19671 3723
rect 19613 3683 19671 3689
rect 19705 3723 19763 3729
rect 19705 3689 19717 3723
rect 19751 3720 19763 3723
rect 19978 3720 19984 3732
rect 19751 3692 19984 3720
rect 19751 3689 19763 3692
rect 19705 3683 19763 3689
rect 19978 3680 19984 3692
rect 20036 3720 20042 3732
rect 20257 3723 20315 3729
rect 20257 3720 20269 3723
rect 20036 3692 20269 3720
rect 20036 3680 20042 3692
rect 20257 3689 20269 3692
rect 20303 3689 20315 3723
rect 20257 3683 20315 3689
rect 22554 3680 22560 3732
rect 22612 3720 22618 3732
rect 22925 3723 22983 3729
rect 22925 3720 22937 3723
rect 22612 3692 22937 3720
rect 22612 3680 22618 3692
rect 22925 3689 22937 3692
rect 22971 3720 22983 3723
rect 23661 3723 23719 3729
rect 23661 3720 23673 3723
rect 22971 3692 23673 3720
rect 22971 3689 22983 3692
rect 22925 3683 22983 3689
rect 23661 3689 23673 3692
rect 23707 3720 23719 3723
rect 23842 3720 23848 3732
rect 23707 3692 23848 3720
rect 23707 3689 23719 3692
rect 23661 3683 23719 3689
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 24394 3720 24400 3732
rect 24355 3692 24400 3720
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 24946 3680 24952 3732
rect 25004 3720 25010 3732
rect 25041 3723 25099 3729
rect 25041 3720 25053 3723
rect 25004 3692 25053 3720
rect 25004 3680 25010 3692
rect 25041 3689 25053 3692
rect 25087 3689 25099 3723
rect 25041 3683 25099 3689
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 25409 3723 25467 3729
rect 25409 3720 25421 3723
rect 25188 3692 25421 3720
rect 25188 3680 25194 3692
rect 25409 3689 25421 3692
rect 25455 3689 25467 3723
rect 25409 3683 25467 3689
rect 10137 3655 10195 3661
rect 10137 3621 10149 3655
rect 10183 3652 10195 3655
rect 15562 3652 15568 3664
rect 10183 3624 13768 3652
rect 15523 3624 15568 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 13740 3596 13768 3624
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 11146 3584 11152 3596
rect 11107 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 12253 3587 12311 3593
rect 12253 3553 12265 3587
rect 12299 3584 12311 3587
rect 12526 3584 12532 3596
rect 12299 3556 12532 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 13722 3584 13728 3596
rect 13683 3556 13728 3584
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 14829 3587 14887 3593
rect 14829 3584 14841 3587
rect 14516 3556 14841 3584
rect 14516 3544 14522 3556
rect 14829 3553 14841 3556
rect 14875 3553 14887 3587
rect 14829 3547 14887 3553
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 16132 3584 16160 3680
rect 20162 3612 20168 3664
rect 20220 3652 20226 3664
rect 20625 3655 20683 3661
rect 20625 3652 20637 3655
rect 20220 3624 20637 3652
rect 20220 3612 20226 3624
rect 20625 3621 20637 3624
rect 20671 3652 20683 3655
rect 21361 3655 21419 3661
rect 21361 3652 21373 3655
rect 20671 3624 21373 3652
rect 20671 3621 20683 3624
rect 20625 3615 20683 3621
rect 21361 3621 21373 3624
rect 21407 3652 21419 3655
rect 22278 3652 22284 3664
rect 21407 3624 22284 3652
rect 21407 3621 21419 3624
rect 21361 3615 21419 3621
rect 15335 3556 16160 3584
rect 17028 3587 17086 3593
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 17028 3553 17040 3587
rect 17074 3584 17086 3587
rect 17310 3584 17316 3596
rect 17074 3556 17316 3584
rect 17074 3553 17086 3556
rect 17028 3547 17086 3553
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 21560 3593 21588 3624
rect 22278 3612 22284 3624
rect 22336 3612 22342 3664
rect 23934 3612 23940 3664
rect 23992 3652 23998 3664
rect 24489 3655 24547 3661
rect 24489 3652 24501 3655
rect 23992 3624 24501 3652
rect 23992 3612 23998 3624
rect 24489 3621 24501 3624
rect 24535 3652 24547 3655
rect 24670 3652 24676 3664
rect 24535 3624 24676 3652
rect 24535 3621 24547 3624
rect 24489 3615 24547 3621
rect 24670 3612 24676 3624
rect 24728 3612 24734 3664
rect 21818 3593 21824 3596
rect 21545 3587 21603 3593
rect 21545 3553 21557 3587
rect 21591 3553 21603 3587
rect 21545 3547 21603 3553
rect 21812 3547 21824 3593
rect 21876 3584 21882 3596
rect 21876 3556 21912 3584
rect 21818 3544 21824 3547
rect 21876 3544 21882 3556
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 13817 3519 13875 3525
rect 13817 3516 13829 3519
rect 12400 3488 13829 3516
rect 12400 3476 12406 3488
rect 13817 3485 13829 3488
rect 13863 3485 13875 3519
rect 13998 3516 14004 3528
rect 13959 3488 14004 3516
rect 13817 3479 13875 3485
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 16758 3516 16764 3528
rect 16592 3488 16764 3516
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12158 3380 12164 3392
rect 11756 3352 12164 3380
rect 11756 3340 11762 3352
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 13630 3380 13636 3392
rect 12483 3352 13636 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 15378 3340 15384 3392
rect 15436 3380 15442 3392
rect 16592 3389 16620 3488
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 19889 3519 19947 3525
rect 19889 3485 19901 3519
rect 19935 3516 19947 3519
rect 20714 3516 20720 3528
rect 19935 3488 20720 3516
rect 19935 3485 19947 3488
rect 19889 3479 19947 3485
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 25038 3516 25044 3528
rect 24627 3488 25044 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 24118 3408 24124 3460
rect 24176 3448 24182 3460
rect 24596 3448 24624 3479
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 24176 3420 24624 3448
rect 24176 3408 24182 3420
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 15436 3352 16589 3380
rect 15436 3340 15442 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 18138 3380 18144 3392
rect 18099 3352 18144 3380
rect 16577 3343 16635 3349
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 19061 3383 19119 3389
rect 19061 3380 19073 3383
rect 18564 3352 19073 3380
rect 18564 3340 18570 3352
rect 19061 3349 19073 3352
rect 19107 3349 19119 3383
rect 19061 3343 19119 3349
rect 23106 3340 23112 3392
rect 23164 3380 23170 3392
rect 24029 3383 24087 3389
rect 24029 3380 24041 3383
rect 23164 3352 24041 3380
rect 23164 3340 23170 3352
rect 24029 3349 24041 3352
rect 24075 3349 24087 3383
rect 24029 3343 24087 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 10778 3176 10784 3188
rect 10739 3148 10784 3176
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12342 3176 12348 3188
rect 12299 3148 12348 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 12621 3179 12679 3185
rect 12621 3176 12633 3179
rect 12584 3148 12633 3176
rect 12584 3136 12590 3148
rect 12621 3145 12633 3148
rect 12667 3145 12679 3179
rect 12621 3139 12679 3145
rect 13998 3136 14004 3188
rect 14056 3176 14062 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 14056 3148 14289 3176
rect 14056 3136 14062 3148
rect 14277 3145 14289 3148
rect 14323 3176 14335 3179
rect 14829 3179 14887 3185
rect 14829 3176 14841 3179
rect 14323 3148 14841 3176
rect 14323 3145 14335 3148
rect 14277 3139 14335 3145
rect 14829 3145 14841 3148
rect 14875 3176 14887 3179
rect 15197 3179 15255 3185
rect 15197 3176 15209 3179
rect 14875 3148 15209 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 15197 3145 15209 3148
rect 15243 3145 15255 3179
rect 15197 3139 15255 3145
rect 10321 3111 10379 3117
rect 10321 3077 10333 3111
rect 10367 3108 10379 3111
rect 10870 3108 10876 3120
rect 10367 3080 10876 3108
rect 10367 3077 10379 3080
rect 10321 3071 10379 3077
rect 10870 3068 10876 3080
rect 10928 3068 10934 3120
rect 11422 3108 11428 3120
rect 11383 3080 11428 3108
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 15212 3040 15240 3139
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17000 3148 17785 3176
rect 17000 3136 17006 3148
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 17773 3139 17831 3145
rect 15212 3012 15516 3040
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10778 2972 10784 2984
rect 10183 2944 10784 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11790 2972 11796 2984
rect 11287 2944 11796 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12216 2944 12909 2972
rect 12216 2932 12222 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 12912 2836 12940 2935
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13153 2975 13211 2981
rect 13153 2972 13165 2975
rect 13044 2944 13165 2972
rect 13044 2932 13050 2944
rect 13153 2941 13165 2944
rect 13199 2972 13211 2975
rect 15381 2975 15439 2981
rect 13199 2944 13308 2972
rect 13199 2941 13211 2944
rect 13153 2935 13211 2941
rect 13280 2916 13308 2944
rect 15381 2941 15393 2975
rect 15427 2941 15439 2975
rect 15488 2972 15516 3012
rect 15637 2975 15695 2981
rect 15637 2972 15649 2975
rect 15488 2944 15649 2972
rect 15381 2935 15439 2941
rect 15637 2941 15649 2944
rect 15683 2941 15695 2975
rect 17788 2972 17816 3139
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 19337 3179 19395 3185
rect 19337 3145 19349 3179
rect 19383 3176 19395 3179
rect 19426 3176 19432 3188
rect 19383 3148 19432 3176
rect 19383 3145 19395 3148
rect 19337 3139 19395 3145
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 21818 3176 21824 3188
rect 21779 3148 21824 3176
rect 21818 3136 21824 3148
rect 21876 3176 21882 3188
rect 22186 3176 22192 3188
rect 21876 3148 22192 3176
rect 21876 3136 21882 3148
rect 22186 3136 22192 3148
rect 22244 3176 22250 3188
rect 22373 3179 22431 3185
rect 22373 3176 22385 3179
rect 22244 3148 22385 3176
rect 22244 3136 22250 3148
rect 22373 3145 22385 3148
rect 22419 3145 22431 3179
rect 23106 3176 23112 3188
rect 23067 3148 23112 3176
rect 22373 3139 22431 3145
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 24118 3176 24124 3188
rect 23523 3148 24124 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 24118 3136 24124 3148
rect 24176 3136 24182 3188
rect 24210 3136 24216 3188
rect 24268 3176 24274 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 24268 3148 24409 3176
rect 24268 3136 24274 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 24397 3139 24455 3145
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 24765 3179 24823 3185
rect 24765 3176 24777 3179
rect 24728 3148 24777 3176
rect 24728 3136 24734 3148
rect 24765 3145 24777 3148
rect 24811 3145 24823 3179
rect 24765 3139 24823 3145
rect 25406 3136 25412 3188
rect 25464 3176 25470 3188
rect 25501 3179 25559 3185
rect 25501 3176 25513 3179
rect 25464 3148 25513 3176
rect 25464 3136 25470 3148
rect 25501 3145 25513 3148
rect 25547 3145 25559 3179
rect 25501 3139 25559 3145
rect 25133 3111 25191 3117
rect 25133 3077 25145 3111
rect 25179 3108 25191 3111
rect 26878 3108 26884 3120
rect 25179 3080 26884 3108
rect 25179 3077 25191 3080
rect 25133 3071 25191 3077
rect 26878 3068 26884 3080
rect 26936 3068 26942 3120
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 18196 3012 18613 3040
rect 18196 3000 18202 3012
rect 18601 3009 18613 3012
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 19751 3012 20361 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 20349 3009 20361 3012
rect 20395 3040 20407 3043
rect 20395 3012 20576 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17788 2944 18429 2972
rect 15637 2935 15695 2941
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 13262 2864 13268 2916
rect 13320 2864 13326 2916
rect 15396 2848 15424 2935
rect 18874 2932 18880 2984
rect 18932 2972 18938 2984
rect 20162 2972 20168 2984
rect 18932 2944 20168 2972
rect 18932 2932 18938 2944
rect 20162 2932 20168 2944
rect 20220 2972 20226 2984
rect 20441 2975 20499 2981
rect 20441 2972 20453 2975
rect 20220 2944 20453 2972
rect 20220 2932 20226 2944
rect 20441 2941 20453 2944
rect 20487 2941 20499 2975
rect 20548 2972 20576 3012
rect 20714 2981 20720 2984
rect 20708 2972 20720 2981
rect 20548 2944 20720 2972
rect 20441 2935 20499 2941
rect 20708 2935 20720 2944
rect 20714 2932 20720 2935
rect 20772 2932 20778 2984
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23532 2944 23673 2972
rect 23532 2932 23538 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 24949 2975 25007 2981
rect 24949 2941 24961 2975
rect 24995 2972 25007 2975
rect 25406 2972 25412 2984
rect 24995 2944 25412 2972
rect 24995 2941 25007 2944
rect 24949 2935 25007 2941
rect 25406 2932 25412 2944
rect 25464 2932 25470 2984
rect 23934 2904 23940 2916
rect 23895 2876 23940 2904
rect 23934 2864 23940 2876
rect 23992 2864 23998 2916
rect 15378 2836 15384 2848
rect 12912 2808 15384 2836
rect 15378 2796 15384 2808
rect 15436 2796 15442 2848
rect 16761 2839 16819 2845
rect 16761 2805 16773 2839
rect 16807 2836 16819 2839
rect 17310 2836 17316 2848
rect 16807 2808 17316 2836
rect 16807 2805 16819 2808
rect 16761 2799 16819 2805
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 18506 2796 18512 2848
rect 18564 2836 18570 2848
rect 18564 2808 18609 2836
rect 18564 2796 18570 2808
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12492 2604 12633 2632
rect 12492 2592 12498 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 13722 2592 13728 2644
rect 13780 2632 13786 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 13780 2604 14013 2632
rect 13780 2592 13786 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 14001 2595 14059 2601
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15378 2632 15384 2644
rect 15335 2604 15384 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 16298 2632 16304 2644
rect 16259 2604 16304 2632
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 17310 2632 17316 2644
rect 17271 2604 17316 2632
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 18138 2632 18144 2644
rect 17819 2604 18144 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 19576 2604 19717 2632
rect 19576 2592 19582 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 21177 2635 21235 2641
rect 21177 2601 21189 2635
rect 21223 2632 21235 2635
rect 22002 2632 22008 2644
rect 21223 2604 22008 2632
rect 21223 2601 21235 2604
rect 21177 2595 21235 2601
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22186 2632 22192 2644
rect 22147 2604 22192 2632
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 22557 2635 22615 2641
rect 22557 2632 22569 2635
rect 22336 2604 22569 2632
rect 22336 2592 22342 2604
rect 22557 2601 22569 2604
rect 22603 2601 22615 2635
rect 22557 2595 22615 2601
rect 23474 2592 23480 2644
rect 23532 2632 23538 2644
rect 23661 2635 23719 2641
rect 23661 2632 23673 2635
rect 23532 2604 23673 2632
rect 23532 2592 23538 2604
rect 23661 2601 23673 2604
rect 23707 2601 23719 2635
rect 23661 2595 23719 2601
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10888 2496 10916 2592
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 13262 2564 13268 2576
rect 11379 2536 13268 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 18874 2564 18880 2576
rect 18340 2536 18880 2564
rect 10367 2468 10916 2496
rect 11425 2499 11483 2505
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11514 2496 11520 2508
rect 11471 2468 11520 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11514 2456 11520 2468
rect 11572 2496 11578 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11572 2468 11989 2496
rect 11572 2456 11578 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 12526 2496 12532 2508
rect 12483 2468 12532 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 12526 2456 12532 2468
rect 12584 2496 12590 2508
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12584 2468 13001 2496
rect 12584 2456 12590 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14826 2496 14832 2508
rect 14323 2468 14832 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 18340 2505 18368 2536
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 23198 2524 23204 2576
rect 23256 2564 23262 2576
rect 24305 2567 24363 2573
rect 24305 2564 24317 2567
rect 23256 2536 24317 2564
rect 23256 2524 23262 2536
rect 24305 2533 24317 2536
rect 24351 2533 24363 2567
rect 24305 2527 24363 2533
rect 16669 2499 16727 2505
rect 16669 2496 16681 2499
rect 16172 2468 16681 2496
rect 16172 2456 16178 2468
rect 16669 2465 16681 2468
rect 16715 2465 16727 2499
rect 16669 2459 16727 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2465 18383 2499
rect 18581 2499 18639 2505
rect 18581 2496 18593 2499
rect 18325 2459 18383 2465
rect 18432 2468 18593 2496
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13262 2428 13268 2440
rect 13223 2400 13268 2428
rect 13081 2391 13139 2397
rect 13096 2360 13124 2391
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 15712 2400 15853 2428
rect 15712 2388 15718 2400
rect 15841 2397 15853 2400
rect 15887 2428 15899 2431
rect 16758 2428 16764 2440
rect 15887 2400 16764 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17310 2428 17316 2440
rect 16991 2400 17316 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18432 2428 18460 2468
rect 18581 2465 18593 2468
rect 18627 2465 18639 2499
rect 20898 2496 20904 2508
rect 20859 2468 20904 2496
rect 18581 2459 18639 2465
rect 20898 2456 20904 2468
rect 20956 2496 20962 2508
rect 21545 2499 21603 2505
rect 21545 2496 21557 2499
rect 20956 2468 21557 2496
rect 20956 2456 20962 2468
rect 21545 2465 21557 2468
rect 21591 2465 21603 2499
rect 22738 2496 22744 2508
rect 22699 2468 22744 2496
rect 21545 2459 21603 2465
rect 22738 2456 22744 2468
rect 22796 2496 22802 2508
rect 23293 2499 23351 2505
rect 23293 2496 23305 2499
rect 22796 2468 23305 2496
rect 22796 2456 22802 2468
rect 23293 2465 23305 2468
rect 23339 2465 23351 2499
rect 23293 2459 23351 2465
rect 23658 2456 23664 2508
rect 23716 2496 23722 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23716 2468 24041 2496
rect 23716 2456 23722 2468
rect 24029 2465 24041 2468
rect 24075 2496 24087 2499
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24075 2468 24777 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 25314 2496 25320 2508
rect 25275 2468 25320 2496
rect 24765 2459 24823 2465
rect 25314 2456 25320 2468
rect 25372 2496 25378 2508
rect 25869 2499 25927 2505
rect 25869 2496 25881 2499
rect 25372 2468 25881 2496
rect 25372 2456 25378 2468
rect 25869 2465 25881 2468
rect 25915 2465 25927 2499
rect 25869 2459 25927 2465
rect 18196 2400 18460 2428
rect 18196 2388 18202 2400
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20588 2400 20637 2428
rect 20588 2388 20594 2400
rect 20625 2397 20637 2400
rect 20671 2428 20683 2431
rect 21634 2428 21640 2440
rect 20671 2400 21640 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 21634 2388 21640 2400
rect 21692 2388 21698 2440
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2428 21879 2431
rect 22186 2428 22192 2440
rect 21867 2400 22192 2428
rect 21867 2397 21879 2400
rect 21821 2391 21879 2397
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 13722 2360 13728 2372
rect 13096 2332 13728 2360
rect 13722 2320 13728 2332
rect 13780 2320 13786 2372
rect 21358 2320 21364 2372
rect 21416 2360 21422 2372
rect 22925 2363 22983 2369
rect 22925 2360 22937 2363
rect 21416 2332 22937 2360
rect 21416 2320 21422 2332
rect 22925 2329 22937 2332
rect 22971 2329 22983 2363
rect 22925 2323 22983 2329
rect 25501 2363 25559 2369
rect 25501 2329 25513 2363
rect 25547 2360 25559 2363
rect 27522 2360 27528 2372
rect 25547 2332 27528 2360
rect 25547 2329 25559 2332
rect 25501 2323 25559 2329
rect 27522 2320 27528 2332
rect 27580 2320 27586 2372
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 10778 2292 10784 2304
rect 10551 2264 10784 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 13078 2292 13084 2304
rect 12584 2264 13084 2292
rect 12584 2252 12590 2264
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 14458 2292 14464 2304
rect 14419 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14826 2292 14832 2304
rect 14787 2264 14832 2292
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 16114 2292 16120 2304
rect 16075 2264 16120 2292
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 21542 552 21548 604
rect 21600 592 21606 604
rect 24118 592 24124 604
rect 21600 564 24124 592
rect 21600 552 21606 564
rect 24118 552 24124 564
rect 24176 552 24182 604
<< via1 >>
rect 21640 26664 21692 26716
rect 24768 26664 24820 26716
rect 16120 26392 16172 26444
rect 24584 26392 24636 26444
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 18696 25440 18748 25492
rect 24676 25440 24728 25492
rect 26884 25372 26936 25424
rect 16396 25304 16448 25356
rect 18880 25347 18932 25356
rect 18880 25313 18889 25347
rect 18889 25313 18923 25347
rect 18923 25313 18932 25347
rect 18880 25304 18932 25313
rect 20260 25304 20312 25356
rect 21824 25304 21876 25356
rect 22836 25347 22888 25356
rect 22836 25313 22845 25347
rect 22845 25313 22879 25347
rect 22879 25313 22888 25347
rect 22836 25304 22888 25313
rect 24032 25304 24084 25356
rect 26148 25236 26200 25288
rect 24124 25168 24176 25220
rect 24768 25143 24820 25152
rect 24768 25109 24777 25143
rect 24777 25109 24811 25143
rect 24811 25109 24820 25143
rect 24768 25100 24820 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 17868 24760 17920 24812
rect 13176 24692 13228 24744
rect 14372 24692 14424 24744
rect 16304 24692 16356 24744
rect 12716 24599 12768 24608
rect 12716 24565 12725 24599
rect 12725 24565 12759 24599
rect 12759 24565 12768 24599
rect 12716 24556 12768 24565
rect 12900 24556 12952 24608
rect 15108 24624 15160 24676
rect 14924 24599 14976 24608
rect 14924 24565 14933 24599
rect 14933 24565 14967 24599
rect 14967 24565 14976 24599
rect 14924 24556 14976 24565
rect 16488 24624 16540 24676
rect 16304 24556 16356 24608
rect 16580 24556 16632 24608
rect 17224 24556 17276 24608
rect 18696 24692 18748 24744
rect 21732 24692 21784 24744
rect 22192 24692 22244 24744
rect 24584 24735 24636 24744
rect 24584 24701 24593 24735
rect 24593 24701 24627 24735
rect 24627 24701 24636 24735
rect 24584 24692 24636 24701
rect 19248 24624 19300 24676
rect 18420 24556 18472 24608
rect 18880 24599 18932 24608
rect 18880 24565 18889 24599
rect 18889 24565 18923 24599
rect 18923 24565 18932 24599
rect 18880 24556 18932 24565
rect 20628 24624 20680 24676
rect 21824 24667 21876 24676
rect 21824 24633 21833 24667
rect 21833 24633 21867 24667
rect 21867 24633 21876 24667
rect 21824 24624 21876 24633
rect 20260 24556 20312 24608
rect 20720 24556 20772 24608
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 22744 24624 22796 24676
rect 22836 24599 22888 24608
rect 22836 24565 22845 24599
rect 22845 24565 22879 24599
rect 22879 24565 22888 24599
rect 22836 24556 22888 24565
rect 24032 24556 24084 24608
rect 24676 24556 24728 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 15844 24395 15896 24404
rect 15844 24361 15853 24395
rect 15853 24361 15887 24395
rect 15887 24361 15896 24395
rect 15844 24352 15896 24361
rect 17316 24352 17368 24404
rect 17960 24352 18012 24404
rect 20076 24352 20128 24404
rect 22008 24352 22060 24404
rect 23388 24352 23440 24404
rect 23664 24395 23716 24404
rect 23664 24361 23673 24395
rect 23673 24361 23707 24395
rect 23707 24361 23716 24395
rect 23664 24352 23716 24361
rect 12716 24216 12768 24268
rect 14740 24216 14792 24268
rect 16948 24259 17000 24268
rect 16948 24225 16957 24259
rect 16957 24225 16991 24259
rect 16991 24225 17000 24259
rect 16948 24216 17000 24225
rect 17592 24216 17644 24268
rect 20168 24216 20220 24268
rect 20996 24259 21048 24268
rect 20996 24225 21005 24259
rect 21005 24225 21039 24259
rect 21039 24225 21048 24259
rect 20996 24216 21048 24225
rect 22376 24259 22428 24268
rect 22376 24225 22385 24259
rect 22385 24225 22419 24259
rect 22419 24225 22428 24259
rect 22376 24216 22428 24225
rect 23480 24259 23532 24268
rect 23480 24225 23489 24259
rect 23489 24225 23523 24259
rect 23523 24225 23532 24259
rect 23480 24216 23532 24225
rect 24768 24216 24820 24268
rect 13268 24191 13320 24200
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 16028 24191 16080 24200
rect 13360 24148 13412 24157
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 11336 24012 11388 24064
rect 12532 24012 12584 24064
rect 12808 24055 12860 24064
rect 12808 24021 12817 24055
rect 12817 24021 12851 24055
rect 12851 24021 12860 24055
rect 12808 24012 12860 24021
rect 14832 24012 14884 24064
rect 16488 24012 16540 24064
rect 22192 24012 22244 24064
rect 24124 24012 24176 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10784 23851 10836 23860
rect 10784 23817 10793 23851
rect 10793 23817 10827 23851
rect 10827 23817 10836 23851
rect 10784 23808 10836 23817
rect 13912 23808 13964 23860
rect 14740 23851 14792 23860
rect 14740 23817 14749 23851
rect 14749 23817 14783 23851
rect 14783 23817 14792 23851
rect 14740 23808 14792 23817
rect 16028 23808 16080 23860
rect 21640 23808 21692 23860
rect 23296 23808 23348 23860
rect 23480 23851 23532 23860
rect 23480 23817 23489 23851
rect 23489 23817 23523 23851
rect 23523 23817 23532 23851
rect 23480 23808 23532 23817
rect 11336 23715 11388 23724
rect 11336 23681 11345 23715
rect 11345 23681 11379 23715
rect 11379 23681 11388 23715
rect 11336 23672 11388 23681
rect 14832 23672 14884 23724
rect 22376 23715 22428 23724
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 23388 23672 23440 23724
rect 11152 23647 11204 23656
rect 11152 23613 11161 23647
rect 11161 23613 11195 23647
rect 11195 23613 11204 23647
rect 11152 23604 11204 23613
rect 13084 23604 13136 23656
rect 16672 23604 16724 23656
rect 18788 23604 18840 23656
rect 21456 23604 21508 23656
rect 15200 23579 15252 23588
rect 15200 23545 15234 23579
rect 15234 23545 15252 23579
rect 15200 23536 15252 23545
rect 18236 23536 18288 23588
rect 20996 23536 21048 23588
rect 21640 23536 21692 23588
rect 23572 23604 23624 23656
rect 25044 23647 25096 23656
rect 25044 23613 25053 23647
rect 25053 23613 25087 23647
rect 25087 23613 25096 23647
rect 25044 23604 25096 23613
rect 10692 23511 10744 23520
rect 10692 23477 10701 23511
rect 10701 23477 10735 23511
rect 10735 23477 10744 23511
rect 11244 23511 11296 23520
rect 10692 23468 10744 23477
rect 11244 23477 11253 23511
rect 11253 23477 11287 23511
rect 11287 23477 11296 23511
rect 11244 23468 11296 23477
rect 12624 23468 12676 23520
rect 12716 23468 12768 23520
rect 13360 23468 13412 23520
rect 16948 23511 17000 23520
rect 16948 23477 16957 23511
rect 16957 23477 16991 23511
rect 16991 23477 17000 23511
rect 16948 23468 17000 23477
rect 17592 23468 17644 23520
rect 19248 23468 19300 23520
rect 20168 23468 20220 23520
rect 23112 23511 23164 23520
rect 23112 23477 23121 23511
rect 23121 23477 23155 23511
rect 23155 23477 23164 23511
rect 23112 23468 23164 23477
rect 24768 23468 24820 23520
rect 25228 23511 25280 23520
rect 25228 23477 25237 23511
rect 25237 23477 25271 23511
rect 25271 23477 25280 23511
rect 25228 23468 25280 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 10968 23264 11020 23316
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 13084 23264 13136 23316
rect 13268 23264 13320 23316
rect 15844 23264 15896 23316
rect 16028 23264 16080 23316
rect 17960 23264 18012 23316
rect 21364 23264 21416 23316
rect 11152 23196 11204 23248
rect 12808 23196 12860 23248
rect 23112 23239 23164 23248
rect 23112 23205 23121 23239
rect 23121 23205 23155 23239
rect 23155 23205 23164 23239
rect 23112 23196 23164 23205
rect 23480 23196 23532 23248
rect 13820 23128 13872 23180
rect 15384 23128 15436 23180
rect 16672 23128 16724 23180
rect 20996 23128 21048 23180
rect 23296 23128 23348 23180
rect 23940 23128 23992 23180
rect 11060 23060 11112 23112
rect 13268 23060 13320 23112
rect 14740 23060 14792 23112
rect 15200 23060 15252 23112
rect 18512 23060 18564 23112
rect 25412 23103 25464 23112
rect 25412 23069 25421 23103
rect 25421 23069 25455 23103
rect 25455 23069 25464 23103
rect 25412 23060 25464 23069
rect 13360 22924 13412 22976
rect 13636 22967 13688 22976
rect 13636 22933 13645 22967
rect 13645 22933 13679 22967
rect 13679 22933 13688 22967
rect 13636 22924 13688 22933
rect 17500 22967 17552 22976
rect 17500 22933 17509 22967
rect 17509 22933 17543 22967
rect 17543 22933 17552 22967
rect 17500 22924 17552 22933
rect 18236 22924 18288 22976
rect 18604 22967 18656 22976
rect 18604 22933 18613 22967
rect 18613 22933 18647 22967
rect 18647 22933 18656 22967
rect 18604 22924 18656 22933
rect 18788 22924 18840 22976
rect 20536 22924 20588 22976
rect 23572 22924 23624 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 12808 22763 12860 22772
rect 12808 22729 12817 22763
rect 12817 22729 12851 22763
rect 12851 22729 12860 22763
rect 12808 22720 12860 22729
rect 13268 22763 13320 22772
rect 13268 22729 13277 22763
rect 13277 22729 13311 22763
rect 13311 22729 13320 22763
rect 13268 22720 13320 22729
rect 14740 22763 14792 22772
rect 14740 22729 14749 22763
rect 14749 22729 14783 22763
rect 14783 22729 14792 22763
rect 14740 22720 14792 22729
rect 16028 22720 16080 22772
rect 17960 22720 18012 22772
rect 21548 22763 21600 22772
rect 21548 22729 21557 22763
rect 21557 22729 21591 22763
rect 21591 22729 21600 22763
rect 21548 22720 21600 22729
rect 23296 22720 23348 22772
rect 11060 22584 11112 22636
rect 12164 22584 12216 22636
rect 12716 22584 12768 22636
rect 16580 22584 16632 22636
rect 24216 22652 24268 22704
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 17500 22584 17552 22636
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 17408 22516 17460 22568
rect 21272 22516 21324 22568
rect 23756 22559 23808 22568
rect 13728 22448 13780 22500
rect 19248 22448 19300 22500
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 13452 22380 13504 22432
rect 16672 22380 16724 22432
rect 18512 22380 18564 22432
rect 20076 22380 20128 22432
rect 20996 22423 21048 22432
rect 20996 22389 21005 22423
rect 21005 22389 21039 22423
rect 21039 22389 21048 22423
rect 20996 22380 21048 22389
rect 22652 22423 22704 22432
rect 22652 22389 22661 22423
rect 22661 22389 22695 22423
rect 22695 22389 22704 22423
rect 22652 22380 22704 22389
rect 23756 22525 23765 22559
rect 23765 22525 23799 22559
rect 23799 22525 23808 22559
rect 23756 22516 23808 22525
rect 25044 22559 25096 22568
rect 25044 22525 25053 22559
rect 25053 22525 25087 22559
rect 25087 22525 25096 22559
rect 25044 22516 25096 22525
rect 23204 22380 23256 22432
rect 24032 22380 24084 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 11152 22176 11204 22228
rect 12716 22176 12768 22228
rect 13176 22176 13228 22228
rect 15384 22176 15436 22228
rect 17040 22176 17092 22228
rect 1400 22040 1452 22092
rect 2320 22040 2372 22092
rect 10048 22040 10100 22092
rect 11060 22083 11112 22092
rect 11060 22049 11069 22083
rect 11069 22049 11103 22083
rect 11103 22049 11112 22083
rect 11060 22040 11112 22049
rect 11796 22040 11848 22092
rect 13360 22040 13412 22092
rect 16948 22108 17000 22160
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 18604 22176 18656 22228
rect 19248 22176 19300 22228
rect 22744 22219 22796 22228
rect 22744 22185 22753 22219
rect 22753 22185 22787 22219
rect 22787 22185 22796 22219
rect 22744 22176 22796 22185
rect 20536 22151 20588 22160
rect 14004 22015 14056 22024
rect 14004 21981 14013 22015
rect 14013 21981 14047 22015
rect 14047 21981 14056 22015
rect 14004 21972 14056 21981
rect 15568 22015 15620 22024
rect 13728 21904 13780 21956
rect 9956 21836 10008 21888
rect 11244 21836 11296 21888
rect 13452 21879 13504 21888
rect 13452 21845 13461 21879
rect 13461 21845 13495 21879
rect 13495 21845 13504 21879
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 16672 21972 16724 22024
rect 18144 22015 18196 22024
rect 18144 21981 18153 22015
rect 18153 21981 18187 22015
rect 18187 21981 18196 22015
rect 20536 22117 20545 22151
rect 20545 22117 20579 22151
rect 20579 22117 20588 22151
rect 20536 22108 20588 22117
rect 18144 21972 18196 21981
rect 15476 21904 15528 21956
rect 15752 21904 15804 21956
rect 20904 22040 20956 22092
rect 21272 22083 21324 22092
rect 21272 22049 21281 22083
rect 21281 22049 21315 22083
rect 21315 22049 21324 22083
rect 21272 22040 21324 22049
rect 23940 22040 23992 22092
rect 22468 21972 22520 22024
rect 22836 22015 22888 22024
rect 22836 21981 22845 22015
rect 22845 21981 22879 22015
rect 22879 21981 22888 22015
rect 22836 21972 22888 21981
rect 23020 22015 23072 22024
rect 23020 21981 23029 22015
rect 23029 21981 23063 22015
rect 23063 21981 23072 22015
rect 23020 21972 23072 21981
rect 19432 21904 19484 21956
rect 21456 21947 21508 21956
rect 21456 21913 21465 21947
rect 21465 21913 21499 21947
rect 21499 21913 21508 21947
rect 21456 21904 21508 21913
rect 14648 21879 14700 21888
rect 13452 21836 13504 21845
rect 14648 21845 14657 21879
rect 14657 21845 14691 21879
rect 14691 21845 14700 21879
rect 14648 21836 14700 21845
rect 14832 21836 14884 21888
rect 16488 21836 16540 21888
rect 17132 21879 17184 21888
rect 17132 21845 17141 21879
rect 17141 21845 17175 21879
rect 17175 21845 17184 21879
rect 17132 21836 17184 21845
rect 22008 21879 22060 21888
rect 22008 21845 22017 21879
rect 22017 21845 22051 21879
rect 22051 21845 22060 21879
rect 22008 21836 22060 21845
rect 22652 21836 22704 21888
rect 24676 21836 24728 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 8392 21632 8444 21684
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12164 21675 12216 21684
rect 12164 21641 12173 21675
rect 12173 21641 12207 21675
rect 12207 21641 12216 21675
rect 12164 21632 12216 21641
rect 13360 21675 13412 21684
rect 13360 21641 13369 21675
rect 13369 21641 13403 21675
rect 13403 21641 13412 21675
rect 13360 21632 13412 21641
rect 9956 21496 10008 21548
rect 11152 21496 11204 21548
rect 13820 21632 13872 21684
rect 14832 21632 14884 21684
rect 15292 21632 15344 21684
rect 16672 21632 16724 21684
rect 17132 21632 17184 21684
rect 19432 21675 19484 21684
rect 19432 21641 19441 21675
rect 19441 21641 19475 21675
rect 19475 21641 19484 21675
rect 19432 21632 19484 21641
rect 22744 21632 22796 21684
rect 23020 21632 23072 21684
rect 23940 21632 23992 21684
rect 14648 21564 14700 21616
rect 15936 21564 15988 21616
rect 15384 21496 15436 21548
rect 16488 21539 16540 21548
rect 16488 21505 16497 21539
rect 16497 21505 16531 21539
rect 16531 21505 16540 21539
rect 16488 21496 16540 21505
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 17132 21428 17184 21480
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 22008 21428 22060 21480
rect 10692 21360 10744 21412
rect 15936 21403 15988 21412
rect 15936 21369 15945 21403
rect 15945 21369 15979 21403
rect 15979 21369 15988 21403
rect 15936 21360 15988 21369
rect 16580 21360 16632 21412
rect 23020 21360 23072 21412
rect 9220 21335 9272 21344
rect 9220 21301 9229 21335
rect 9229 21301 9263 21335
rect 9263 21301 9272 21335
rect 9220 21292 9272 21301
rect 9312 21292 9364 21344
rect 10968 21292 11020 21344
rect 11244 21335 11296 21344
rect 11244 21301 11253 21335
rect 11253 21301 11287 21335
rect 11287 21301 11296 21335
rect 11244 21292 11296 21301
rect 12532 21292 12584 21344
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 14004 21292 14056 21301
rect 14648 21292 14700 21344
rect 16028 21335 16080 21344
rect 16028 21301 16037 21335
rect 16037 21301 16071 21335
rect 16071 21301 16080 21335
rect 16028 21292 16080 21301
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 19524 21292 19576 21344
rect 20444 21335 20496 21344
rect 20444 21301 20453 21335
rect 20453 21301 20487 21335
rect 20487 21301 20496 21335
rect 20444 21292 20496 21301
rect 22284 21292 22336 21344
rect 22468 21335 22520 21344
rect 22468 21301 22477 21335
rect 22477 21301 22511 21335
rect 22511 21301 22520 21335
rect 22468 21292 22520 21301
rect 23940 21292 23992 21344
rect 24584 21403 24636 21412
rect 24584 21369 24593 21403
rect 24593 21369 24627 21403
rect 24627 21369 24636 21403
rect 24584 21360 24636 21369
rect 24860 21292 24912 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 11244 21088 11296 21140
rect 13452 21088 13504 21140
rect 16028 21088 16080 21140
rect 16856 21088 16908 21140
rect 18144 21088 18196 21140
rect 19984 21088 20036 21140
rect 21272 21088 21324 21140
rect 21824 21131 21876 21140
rect 21824 21097 21833 21131
rect 21833 21097 21867 21131
rect 21867 21097 21876 21131
rect 21824 21088 21876 21097
rect 13176 21020 13228 21072
rect 13912 21063 13964 21072
rect 13912 21029 13921 21063
rect 13921 21029 13955 21063
rect 13955 21029 13964 21063
rect 13912 21020 13964 21029
rect 9956 20952 10008 21004
rect 12440 20995 12492 21004
rect 12440 20961 12449 20995
rect 12449 20961 12483 20995
rect 12483 20961 12492 20995
rect 12440 20952 12492 20961
rect 13360 20952 13412 21004
rect 15384 21020 15436 21072
rect 22284 21063 22336 21072
rect 22284 21029 22318 21063
rect 22318 21029 22336 21063
rect 22284 21020 22336 21029
rect 24768 21063 24820 21072
rect 24768 21029 24777 21063
rect 24777 21029 24811 21063
rect 24811 21029 24820 21063
rect 24768 21020 24820 21029
rect 18144 20995 18196 21004
rect 18144 20961 18153 20995
rect 18153 20961 18187 20995
rect 18187 20961 18196 20995
rect 18144 20952 18196 20961
rect 19524 20995 19576 21004
rect 19524 20961 19533 20995
rect 19533 20961 19567 20995
rect 19567 20961 19576 20995
rect 19524 20952 19576 20961
rect 20352 20995 20404 21004
rect 20352 20961 20361 20995
rect 20361 20961 20395 20995
rect 20395 20961 20404 20995
rect 20352 20952 20404 20961
rect 20904 20995 20956 21004
rect 20904 20961 20913 20995
rect 20913 20961 20947 20995
rect 20947 20961 20956 20995
rect 20904 20952 20956 20961
rect 22008 20995 22060 21004
rect 22008 20961 22017 20995
rect 22017 20961 22051 20995
rect 22051 20961 22060 20995
rect 22008 20952 22060 20961
rect 24124 20952 24176 21004
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 11796 20816 11848 20868
rect 17960 20884 18012 20936
rect 7656 20791 7708 20800
rect 7656 20757 7665 20791
rect 7665 20757 7699 20791
rect 7699 20757 7708 20791
rect 7656 20748 7708 20757
rect 9312 20791 9364 20800
rect 9312 20757 9321 20791
rect 9321 20757 9355 20791
rect 9355 20757 9364 20791
rect 9312 20748 9364 20757
rect 14648 20748 14700 20800
rect 15936 20748 15988 20800
rect 16764 20748 16816 20800
rect 18788 20791 18840 20800
rect 18788 20757 18797 20791
rect 18797 20757 18831 20791
rect 18831 20757 18840 20791
rect 18788 20748 18840 20757
rect 19156 20791 19208 20800
rect 19156 20757 19165 20791
rect 19165 20757 19199 20791
rect 19199 20757 19208 20791
rect 19156 20748 19208 20757
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 21088 20791 21140 20800
rect 21088 20757 21097 20791
rect 21097 20757 21131 20791
rect 21131 20757 21140 20791
rect 21088 20748 21140 20757
rect 22008 20748 22060 20800
rect 23664 20816 23716 20868
rect 23296 20748 23348 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 9680 20544 9732 20596
rect 10048 20544 10100 20596
rect 10692 20544 10744 20596
rect 11796 20587 11848 20596
rect 11796 20553 11805 20587
rect 11805 20553 11839 20587
rect 11839 20553 11848 20587
rect 11796 20544 11848 20553
rect 15384 20544 15436 20596
rect 16028 20544 16080 20596
rect 16212 20544 16264 20596
rect 17868 20544 17920 20596
rect 23020 20587 23072 20596
rect 23020 20553 23029 20587
rect 23029 20553 23063 20587
rect 23063 20553 23072 20587
rect 23020 20544 23072 20553
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 13912 20451 13964 20460
rect 13912 20417 13921 20451
rect 13921 20417 13955 20451
rect 13955 20417 13964 20451
rect 13912 20408 13964 20417
rect 7656 20340 7708 20392
rect 12164 20340 12216 20392
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17224 20408 17276 20460
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 18788 20340 18840 20392
rect 19340 20340 19392 20392
rect 20536 20340 20588 20392
rect 7840 20315 7892 20324
rect 7840 20281 7874 20315
rect 7874 20281 7892 20315
rect 7840 20272 7892 20281
rect 12348 20272 12400 20324
rect 14188 20315 14240 20324
rect 14188 20281 14211 20315
rect 14211 20281 14240 20315
rect 14188 20272 14240 20281
rect 16212 20315 16264 20324
rect 16212 20281 16221 20315
rect 16221 20281 16255 20315
rect 16255 20281 16264 20315
rect 16212 20272 16264 20281
rect 16764 20315 16816 20324
rect 16764 20281 16773 20315
rect 16773 20281 16807 20315
rect 16807 20281 16816 20315
rect 16764 20272 16816 20281
rect 18328 20315 18380 20324
rect 18328 20281 18337 20315
rect 18337 20281 18371 20315
rect 18371 20281 18380 20315
rect 18328 20272 18380 20281
rect 20076 20272 20128 20324
rect 20812 20272 20864 20324
rect 22928 20272 22980 20324
rect 23296 20272 23348 20324
rect 8024 20204 8076 20256
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 10784 20204 10836 20256
rect 11244 20247 11296 20256
rect 11244 20213 11253 20247
rect 11253 20213 11287 20247
rect 11287 20213 11296 20247
rect 11244 20204 11296 20213
rect 13360 20204 13412 20256
rect 15936 20204 15988 20256
rect 18788 20247 18840 20256
rect 18788 20213 18797 20247
rect 18797 20213 18831 20247
rect 18831 20213 18840 20247
rect 18788 20204 18840 20213
rect 19984 20204 20036 20256
rect 20444 20204 20496 20256
rect 22008 20247 22060 20256
rect 22008 20213 22017 20247
rect 22017 20213 22051 20247
rect 22051 20213 22060 20247
rect 22008 20204 22060 20213
rect 22100 20204 22152 20256
rect 24584 20204 24636 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 7840 20043 7892 20052
rect 7840 20009 7849 20043
rect 7849 20009 7883 20043
rect 7883 20009 7892 20043
rect 7840 20000 7892 20009
rect 9956 20000 10008 20052
rect 12624 20000 12676 20052
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 16764 20000 16816 20052
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 19524 20000 19576 20052
rect 20536 20000 20588 20052
rect 22008 20000 22060 20052
rect 23296 20000 23348 20052
rect 24768 20000 24820 20052
rect 18604 19932 18656 19984
rect 21180 19975 21232 19984
rect 21180 19941 21189 19975
rect 21189 19941 21223 19975
rect 21223 19941 21232 19975
rect 21180 19932 21232 19941
rect 22100 19975 22152 19984
rect 22100 19941 22109 19975
rect 22109 19941 22143 19975
rect 22143 19941 22152 19975
rect 22100 19932 22152 19941
rect 7748 19907 7800 19916
rect 7748 19873 7757 19907
rect 7757 19873 7791 19907
rect 7791 19873 7800 19907
rect 7748 19864 7800 19873
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 9956 19907 10008 19916
rect 9956 19873 9990 19907
rect 9990 19873 10008 19907
rect 9956 19864 10008 19873
rect 11060 19864 11112 19916
rect 12164 19907 12216 19916
rect 12164 19873 12173 19907
rect 12173 19873 12207 19907
rect 12207 19873 12216 19907
rect 12164 19864 12216 19873
rect 14280 19864 14332 19916
rect 15936 19864 15988 19916
rect 18052 19864 18104 19916
rect 19156 19864 19208 19916
rect 19616 19907 19668 19916
rect 19616 19873 19625 19907
rect 19625 19873 19659 19907
rect 19659 19873 19668 19907
rect 19616 19864 19668 19873
rect 22744 19907 22796 19916
rect 8024 19839 8076 19848
rect 8024 19805 8033 19839
rect 8033 19805 8067 19839
rect 8067 19805 8076 19839
rect 8024 19796 8076 19805
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12851 19839
rect 12851 19805 12860 19839
rect 12808 19796 12860 19805
rect 11888 19728 11940 19780
rect 15568 19796 15620 19848
rect 19524 19796 19576 19848
rect 19984 19796 20036 19848
rect 22744 19873 22753 19907
rect 22753 19873 22787 19907
rect 22787 19873 22796 19907
rect 22744 19864 22796 19873
rect 24400 19907 24452 19916
rect 24400 19873 24409 19907
rect 24409 19873 24443 19907
rect 24443 19873 24452 19907
rect 24400 19864 24452 19873
rect 22928 19839 22980 19848
rect 22928 19805 22937 19839
rect 22937 19805 22971 19839
rect 22971 19805 22980 19839
rect 22928 19796 22980 19805
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 24860 19796 24912 19848
rect 24124 19728 24176 19780
rect 8208 19660 8260 19712
rect 12256 19660 12308 19712
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 13820 19703 13872 19712
rect 13820 19669 13829 19703
rect 13829 19669 13863 19703
rect 13863 19669 13872 19703
rect 13820 19660 13872 19669
rect 18420 19660 18472 19712
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 7840 19456 7892 19508
rect 9956 19499 10008 19508
rect 9956 19465 9965 19499
rect 9965 19465 9999 19499
rect 9999 19465 10008 19499
rect 9956 19456 10008 19465
rect 11888 19499 11940 19508
rect 11888 19465 11897 19499
rect 11897 19465 11931 19499
rect 11931 19465 11940 19499
rect 11888 19456 11940 19465
rect 16396 19499 16448 19508
rect 16396 19465 16405 19499
rect 16405 19465 16439 19499
rect 16439 19465 16448 19499
rect 16396 19456 16448 19465
rect 19616 19456 19668 19508
rect 22928 19456 22980 19508
rect 23664 19456 23716 19508
rect 7564 19252 7616 19304
rect 7840 19227 7892 19236
rect 7840 19193 7849 19227
rect 7849 19193 7883 19227
rect 7883 19193 7892 19227
rect 7840 19184 7892 19193
rect 8116 19252 8168 19304
rect 12624 19320 12676 19372
rect 16028 19320 16080 19372
rect 18604 19363 18656 19372
rect 18604 19329 18613 19363
rect 18613 19329 18647 19363
rect 18647 19329 18656 19363
rect 18604 19320 18656 19329
rect 22192 19388 22244 19440
rect 24032 19456 24084 19508
rect 20076 19320 20128 19372
rect 21824 19363 21876 19372
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 24032 19320 24084 19372
rect 8392 19184 8444 19236
rect 10600 19227 10652 19236
rect 10600 19193 10609 19227
rect 10609 19193 10643 19227
rect 10643 19193 10652 19227
rect 10600 19184 10652 19193
rect 13360 19252 13412 19304
rect 16856 19252 16908 19304
rect 18144 19252 18196 19304
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 19248 19252 19300 19304
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 23112 19295 23164 19304
rect 23112 19261 23121 19295
rect 23121 19261 23155 19295
rect 23155 19261 23164 19295
rect 24492 19320 24544 19372
rect 24860 19320 24912 19372
rect 25044 19295 25096 19304
rect 23112 19252 23164 19261
rect 25044 19261 25053 19295
rect 25053 19261 25087 19295
rect 25087 19261 25096 19295
rect 25044 19252 25096 19261
rect 25228 19295 25280 19304
rect 25228 19261 25237 19295
rect 25237 19261 25271 19295
rect 25271 19261 25280 19295
rect 25228 19252 25280 19261
rect 13820 19184 13872 19236
rect 21916 19184 21968 19236
rect 23480 19227 23532 19236
rect 23480 19193 23489 19227
rect 23489 19193 23523 19227
rect 23523 19193 23532 19227
rect 25504 19227 25556 19236
rect 23480 19184 23532 19193
rect 9404 19159 9456 19168
rect 9404 19125 9413 19159
rect 9413 19125 9447 19159
rect 9447 19125 9456 19159
rect 9404 19116 9456 19125
rect 10876 19116 10928 19168
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 12072 19116 12124 19168
rect 12808 19116 12860 19168
rect 14188 19159 14240 19168
rect 14188 19125 14197 19159
rect 14197 19125 14231 19159
rect 14231 19125 14240 19159
rect 14188 19116 14240 19125
rect 14280 19116 14332 19168
rect 15568 19116 15620 19168
rect 17132 19116 17184 19168
rect 17960 19116 18012 19168
rect 18144 19116 18196 19168
rect 19248 19116 19300 19168
rect 19340 19116 19392 19168
rect 20720 19116 20772 19168
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 22468 19116 22520 19168
rect 24032 19159 24084 19168
rect 24032 19125 24041 19159
rect 24041 19125 24075 19159
rect 24075 19125 24084 19159
rect 24032 19116 24084 19125
rect 25504 19193 25513 19227
rect 25513 19193 25547 19227
rect 25547 19193 25556 19227
rect 25504 19184 25556 19193
rect 24216 19116 24268 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 8024 18955 8076 18964
rect 8024 18921 8033 18955
rect 8033 18921 8067 18955
rect 8067 18921 8076 18955
rect 8024 18912 8076 18921
rect 8392 18955 8444 18964
rect 8392 18921 8401 18955
rect 8401 18921 8435 18955
rect 8435 18921 8444 18955
rect 8392 18912 8444 18921
rect 9312 18955 9364 18964
rect 9312 18921 9321 18955
rect 9321 18921 9355 18955
rect 9355 18921 9364 18955
rect 9312 18912 9364 18921
rect 11796 18912 11848 18964
rect 13360 18912 13412 18964
rect 15936 18955 15988 18964
rect 15936 18921 15945 18955
rect 15945 18921 15979 18955
rect 15979 18921 15988 18955
rect 15936 18912 15988 18921
rect 19524 18912 19576 18964
rect 21272 18912 21324 18964
rect 22100 18955 22152 18964
rect 22100 18921 22109 18955
rect 22109 18921 22143 18955
rect 22143 18921 22152 18955
rect 22100 18912 22152 18921
rect 24768 18912 24820 18964
rect 10140 18844 10192 18896
rect 11152 18844 11204 18896
rect 11888 18844 11940 18896
rect 12348 18844 12400 18896
rect 17960 18844 18012 18896
rect 19984 18844 20036 18896
rect 20076 18844 20128 18896
rect 21824 18844 21876 18896
rect 23112 18844 23164 18896
rect 24492 18887 24544 18896
rect 24492 18853 24501 18887
rect 24501 18853 24535 18887
rect 24535 18853 24544 18887
rect 24492 18844 24544 18853
rect 8392 18776 8444 18828
rect 8760 18819 8812 18828
rect 8760 18785 8769 18819
rect 8769 18785 8803 18819
rect 8803 18785 8812 18819
rect 8760 18776 8812 18785
rect 10048 18819 10100 18828
rect 10048 18785 10057 18819
rect 10057 18785 10091 18819
rect 10091 18785 10100 18819
rect 10048 18776 10100 18785
rect 11428 18776 11480 18828
rect 11796 18819 11848 18828
rect 11796 18785 11805 18819
rect 11805 18785 11839 18819
rect 11839 18785 11848 18819
rect 11796 18776 11848 18785
rect 14832 18776 14884 18828
rect 16028 18776 16080 18828
rect 17408 18776 17460 18828
rect 18420 18819 18472 18828
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 21088 18819 21140 18828
rect 21088 18785 21097 18819
rect 21097 18785 21131 18819
rect 21131 18785 21140 18819
rect 21088 18776 21140 18785
rect 21364 18776 21416 18828
rect 25044 18819 25096 18828
rect 25044 18785 25053 18819
rect 25053 18785 25087 18819
rect 25087 18785 25096 18819
rect 25044 18776 25096 18785
rect 25136 18819 25188 18828
rect 25136 18785 25145 18819
rect 25145 18785 25179 18819
rect 25179 18785 25188 18819
rect 25136 18776 25188 18785
rect 25412 18776 25464 18828
rect 9680 18708 9732 18760
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 15292 18751 15344 18760
rect 9956 18640 10008 18692
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 16580 18708 16632 18760
rect 17500 18708 17552 18760
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 20628 18708 20680 18760
rect 22100 18708 22152 18760
rect 25228 18751 25280 18760
rect 25228 18717 25237 18751
rect 25237 18717 25271 18751
rect 25271 18717 25280 18751
rect 25228 18708 25280 18717
rect 17408 18640 17460 18692
rect 9680 18615 9732 18624
rect 9680 18581 9689 18615
rect 9689 18581 9723 18615
rect 9723 18581 9732 18615
rect 9680 18572 9732 18581
rect 13728 18615 13780 18624
rect 13728 18581 13737 18615
rect 13737 18581 13771 18615
rect 13771 18581 13780 18615
rect 13728 18572 13780 18581
rect 14280 18615 14332 18624
rect 14280 18581 14289 18615
rect 14289 18581 14323 18615
rect 14323 18581 14332 18615
rect 14280 18572 14332 18581
rect 15476 18572 15528 18624
rect 16212 18615 16264 18624
rect 16212 18581 16221 18615
rect 16221 18581 16255 18615
rect 16255 18581 16264 18615
rect 16212 18572 16264 18581
rect 16488 18615 16540 18624
rect 16488 18581 16497 18615
rect 16497 18581 16531 18615
rect 16531 18581 16540 18615
rect 16488 18572 16540 18581
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 23480 18572 23532 18624
rect 24676 18615 24728 18624
rect 24676 18581 24685 18615
rect 24685 18581 24719 18615
rect 24719 18581 24728 18615
rect 24676 18572 24728 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 9956 18368 10008 18420
rect 11428 18411 11480 18420
rect 11428 18377 11437 18411
rect 11437 18377 11471 18411
rect 11471 18377 11480 18411
rect 11428 18368 11480 18377
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 12348 18368 12400 18420
rect 13912 18368 13964 18420
rect 14096 18368 14148 18420
rect 14832 18368 14884 18420
rect 20352 18368 20404 18420
rect 20536 18368 20588 18420
rect 21088 18411 21140 18420
rect 21088 18377 21097 18411
rect 21097 18377 21131 18411
rect 21131 18377 21140 18411
rect 21088 18368 21140 18377
rect 22008 18411 22060 18420
rect 22008 18377 22017 18411
rect 22017 18377 22051 18411
rect 22051 18377 22060 18411
rect 22008 18368 22060 18377
rect 23112 18411 23164 18420
rect 23112 18377 23121 18411
rect 23121 18377 23155 18411
rect 23155 18377 23164 18411
rect 23112 18368 23164 18377
rect 25228 18368 25280 18420
rect 15384 18300 15436 18352
rect 20996 18300 21048 18352
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 10140 18232 10192 18284
rect 14188 18232 14240 18284
rect 15476 18275 15528 18284
rect 15476 18241 15485 18275
rect 15485 18241 15519 18275
rect 15519 18241 15528 18275
rect 15476 18232 15528 18241
rect 15568 18232 15620 18284
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 9404 18164 9456 18216
rect 13728 18164 13780 18216
rect 16396 18164 16448 18216
rect 16580 18164 16632 18216
rect 23480 18232 23532 18284
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 23296 18164 23348 18216
rect 12348 18096 12400 18148
rect 13636 18028 13688 18080
rect 14832 18096 14884 18148
rect 17684 18096 17736 18148
rect 18604 18139 18656 18148
rect 18604 18105 18638 18139
rect 18638 18105 18656 18139
rect 18604 18096 18656 18105
rect 19156 18096 19208 18148
rect 23204 18096 23256 18148
rect 14280 18071 14332 18080
rect 14280 18037 14289 18071
rect 14289 18037 14323 18071
rect 14323 18037 14332 18071
rect 14280 18028 14332 18037
rect 14740 18028 14792 18080
rect 14924 18028 14976 18080
rect 15568 18028 15620 18080
rect 16028 18028 16080 18080
rect 17408 18028 17460 18080
rect 19984 18028 20036 18080
rect 23112 18028 23164 18080
rect 24032 18028 24084 18080
rect 25136 18028 25188 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 8300 17824 8352 17876
rect 9588 17824 9640 17876
rect 9680 17824 9732 17876
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 10876 17824 10928 17876
rect 12348 17824 12400 17876
rect 13728 17824 13780 17876
rect 14280 17824 14332 17876
rect 16580 17824 16632 17876
rect 17868 17824 17920 17876
rect 19156 17867 19208 17876
rect 19156 17833 19165 17867
rect 19165 17833 19199 17867
rect 19199 17833 19208 17867
rect 19156 17824 19208 17833
rect 23204 17824 23256 17876
rect 23940 17867 23992 17876
rect 23940 17833 23949 17867
rect 23949 17833 23983 17867
rect 23983 17833 23992 17867
rect 23940 17824 23992 17833
rect 24676 17824 24728 17876
rect 25228 17824 25280 17876
rect 12164 17756 12216 17808
rect 13820 17756 13872 17808
rect 10508 17688 10560 17740
rect 14096 17731 14148 17740
rect 14096 17697 14105 17731
rect 14105 17697 14139 17731
rect 14139 17697 14148 17731
rect 14096 17688 14148 17697
rect 16212 17756 16264 17808
rect 15568 17731 15620 17740
rect 15568 17697 15602 17731
rect 15602 17697 15620 17731
rect 15568 17688 15620 17697
rect 9956 17620 10008 17672
rect 12716 17663 12768 17672
rect 10048 17552 10100 17604
rect 9404 17484 9456 17536
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 13360 17620 13412 17672
rect 14924 17663 14976 17672
rect 14096 17552 14148 17604
rect 14924 17629 14933 17663
rect 14933 17629 14967 17663
rect 14967 17629 14976 17663
rect 14924 17620 14976 17629
rect 19064 17688 19116 17740
rect 19432 17688 19484 17740
rect 22100 17756 22152 17808
rect 22560 17756 22612 17808
rect 21180 17731 21232 17740
rect 21180 17697 21214 17731
rect 21214 17697 21232 17731
rect 21180 17688 21232 17697
rect 24032 17688 24084 17740
rect 25596 17688 25648 17740
rect 16672 17595 16724 17604
rect 16672 17561 16681 17595
rect 16681 17561 16715 17595
rect 16715 17561 16724 17595
rect 16672 17552 16724 17561
rect 13176 17527 13228 17536
rect 13176 17493 13185 17527
rect 13185 17493 13219 17527
rect 13219 17493 13228 17527
rect 13176 17484 13228 17493
rect 19524 17484 19576 17536
rect 24216 17620 24268 17672
rect 25412 17552 25464 17604
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 23296 17527 23348 17536
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23756 17527 23808 17536
rect 23296 17484 23348 17493
rect 23756 17493 23765 17527
rect 23765 17493 23799 17527
rect 23799 17493 23808 17527
rect 23756 17484 23808 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 9496 17280 9548 17332
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 12716 17280 12768 17332
rect 14280 17280 14332 17332
rect 9404 17212 9456 17264
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 11428 17212 11480 17264
rect 13820 17212 13872 17264
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 12256 17119 12308 17128
rect 12256 17085 12265 17119
rect 12265 17085 12299 17119
rect 12299 17085 12308 17119
rect 12256 17076 12308 17085
rect 12900 17119 12952 17128
rect 12900 17085 12909 17119
rect 12909 17085 12943 17119
rect 12943 17085 12952 17119
rect 12900 17076 12952 17085
rect 9496 17051 9548 17060
rect 9496 17017 9505 17051
rect 9505 17017 9539 17051
rect 9539 17017 9548 17051
rect 9496 17008 9548 17017
rect 15292 17280 15344 17332
rect 17868 17280 17920 17332
rect 19432 17280 19484 17332
rect 24676 17280 24728 17332
rect 25596 17323 25648 17332
rect 25596 17289 25605 17323
rect 25605 17289 25639 17323
rect 25639 17289 25648 17323
rect 25596 17280 25648 17289
rect 15384 17144 15436 17196
rect 16304 17144 16356 17196
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 17500 17187 17552 17196
rect 16672 17144 16724 17153
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 18696 17187 18748 17196
rect 17500 17144 17552 17153
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 16488 17119 16540 17128
rect 16488 17085 16497 17119
rect 16497 17085 16531 17119
rect 16531 17085 16540 17119
rect 16488 17076 16540 17085
rect 18512 17076 18564 17128
rect 19524 17076 19576 17128
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 23756 17076 23808 17128
rect 25504 17076 25556 17128
rect 18144 17008 18196 17060
rect 10048 16940 10100 16992
rect 12440 16940 12492 16992
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 13636 16983 13688 16992
rect 13636 16949 13645 16983
rect 13645 16949 13679 16983
rect 13679 16949 13688 16983
rect 13636 16940 13688 16949
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 15568 16940 15620 16949
rect 16212 16940 16264 16992
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 19248 17008 19300 17060
rect 20260 17008 20312 17060
rect 23940 17051 23992 17060
rect 23940 17017 23974 17051
rect 23974 17017 23992 17051
rect 23940 17008 23992 17017
rect 19064 16983 19116 16992
rect 19064 16949 19073 16983
rect 19073 16949 19107 16983
rect 19107 16949 19116 16983
rect 19064 16940 19116 16949
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 21180 16940 21232 16992
rect 23480 16983 23532 16992
rect 23480 16949 23489 16983
rect 23489 16949 23523 16983
rect 23523 16949 23532 16983
rect 23480 16940 23532 16949
rect 24216 16940 24268 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 9404 16736 9456 16788
rect 12716 16736 12768 16788
rect 13452 16736 13504 16788
rect 14740 16779 14792 16788
rect 14740 16745 14749 16779
rect 14749 16745 14783 16779
rect 14783 16745 14792 16779
rect 14740 16736 14792 16745
rect 16304 16779 16356 16788
rect 16304 16745 16313 16779
rect 16313 16745 16347 16779
rect 16347 16745 16356 16779
rect 16304 16736 16356 16745
rect 16488 16736 16540 16788
rect 18144 16736 18196 16788
rect 18420 16779 18472 16788
rect 18420 16745 18429 16779
rect 18429 16745 18463 16779
rect 18463 16745 18472 16779
rect 18420 16736 18472 16745
rect 20260 16779 20312 16788
rect 20260 16745 20269 16779
rect 20269 16745 20303 16779
rect 20303 16745 20312 16779
rect 20260 16736 20312 16745
rect 21824 16736 21876 16788
rect 22100 16736 22152 16788
rect 22468 16779 22520 16788
rect 22468 16745 22477 16779
rect 22477 16745 22511 16779
rect 22511 16745 22520 16779
rect 22468 16736 22520 16745
rect 24032 16779 24084 16788
rect 24032 16745 24041 16779
rect 24041 16745 24075 16779
rect 24075 16745 24084 16779
rect 24032 16736 24084 16745
rect 24492 16779 24544 16788
rect 24492 16745 24501 16779
rect 24501 16745 24535 16779
rect 24535 16745 24544 16779
rect 24492 16736 24544 16745
rect 14464 16668 14516 16720
rect 17592 16668 17644 16720
rect 18052 16668 18104 16720
rect 18972 16668 19024 16720
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 11704 16643 11756 16652
rect 11704 16609 11738 16643
rect 11738 16609 11756 16643
rect 11704 16600 11756 16609
rect 13912 16643 13964 16652
rect 13912 16609 13921 16643
rect 13921 16609 13955 16643
rect 13955 16609 13964 16643
rect 13912 16600 13964 16609
rect 15568 16600 15620 16652
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 16672 16600 16724 16652
rect 18144 16600 18196 16652
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 18512 16532 18564 16584
rect 19064 16575 19116 16584
rect 19064 16541 19073 16575
rect 19073 16541 19107 16575
rect 19107 16541 19116 16575
rect 19064 16532 19116 16541
rect 18420 16464 18472 16516
rect 21272 16643 21324 16652
rect 21272 16609 21281 16643
rect 21281 16609 21315 16643
rect 21315 16609 21324 16643
rect 21272 16600 21324 16609
rect 21640 16600 21692 16652
rect 22100 16600 22152 16652
rect 23940 16668 23992 16720
rect 23112 16600 23164 16652
rect 24400 16643 24452 16652
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 22744 16532 22796 16584
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 25228 16668 25280 16720
rect 23020 16532 23072 16541
rect 25504 16643 25556 16652
rect 25504 16609 25513 16643
rect 25513 16609 25547 16643
rect 25547 16609 25556 16643
rect 25504 16600 25556 16609
rect 26148 16600 26200 16652
rect 24124 16464 24176 16516
rect 11428 16396 11480 16448
rect 12716 16396 12768 16448
rect 15476 16396 15528 16448
rect 18512 16396 18564 16448
rect 20536 16439 20588 16448
rect 20536 16405 20545 16439
rect 20545 16405 20579 16439
rect 20579 16405 20588 16439
rect 20536 16396 20588 16405
rect 20720 16396 20772 16448
rect 23572 16396 23624 16448
rect 23848 16396 23900 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 11704 16192 11756 16244
rect 15384 16235 15436 16244
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 17408 16192 17460 16244
rect 17592 16192 17644 16244
rect 17960 16192 18012 16244
rect 19064 16235 19116 16244
rect 19064 16201 19073 16235
rect 19073 16201 19107 16235
rect 19107 16201 19116 16235
rect 19064 16192 19116 16201
rect 24032 16192 24084 16244
rect 24676 16235 24728 16244
rect 24676 16201 24685 16235
rect 24685 16201 24719 16235
rect 24719 16201 24728 16235
rect 24676 16192 24728 16201
rect 25228 16192 25280 16244
rect 13912 16124 13964 16176
rect 20536 16124 20588 16176
rect 23296 16124 23348 16176
rect 11428 16099 11480 16108
rect 11152 15988 11204 16040
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 13820 16056 13872 16108
rect 14004 16099 14056 16108
rect 14004 16065 14013 16099
rect 14013 16065 14047 16099
rect 14047 16065 14056 16099
rect 14004 16056 14056 16065
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 17500 16056 17552 16108
rect 12348 15988 12400 16040
rect 14280 16031 14332 16040
rect 14280 15997 14314 16031
rect 14314 15997 14332 16031
rect 14280 15988 14332 15997
rect 16304 15988 16356 16040
rect 17868 15988 17920 16040
rect 16948 15963 17000 15972
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 11980 15852 12032 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 16948 15929 16957 15963
rect 16957 15929 16991 15963
rect 16991 15929 17000 15963
rect 16948 15920 17000 15929
rect 20076 16056 20128 16108
rect 21824 16056 21876 16108
rect 23756 16056 23808 16108
rect 24584 16056 24636 16108
rect 20536 15988 20588 16040
rect 24032 16031 24084 16040
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 24032 15988 24084 15997
rect 25228 16031 25280 16040
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 16672 15852 16724 15904
rect 16764 15852 16816 15904
rect 18420 15895 18472 15904
rect 18420 15861 18429 15895
rect 18429 15861 18463 15895
rect 18463 15861 18472 15895
rect 18420 15852 18472 15861
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 20076 15895 20128 15904
rect 18512 15852 18564 15861
rect 20076 15861 20085 15895
rect 20085 15861 20119 15895
rect 20119 15861 20128 15895
rect 20076 15852 20128 15861
rect 21640 15920 21692 15972
rect 21732 15920 21784 15972
rect 22100 15963 22152 15972
rect 22100 15929 22109 15963
rect 22109 15929 22143 15963
rect 22143 15929 22152 15963
rect 25504 15963 25556 15972
rect 22100 15920 22152 15929
rect 25504 15929 25513 15963
rect 25513 15929 25547 15963
rect 25547 15929 25556 15963
rect 25504 15920 25556 15929
rect 20904 15852 20956 15904
rect 21272 15852 21324 15904
rect 21916 15852 21968 15904
rect 22744 15895 22796 15904
rect 22744 15861 22753 15895
rect 22753 15861 22787 15895
rect 22787 15861 22796 15895
rect 22744 15852 22796 15861
rect 23112 15895 23164 15904
rect 23112 15861 23121 15895
rect 23121 15861 23155 15895
rect 23155 15861 23164 15895
rect 23112 15852 23164 15861
rect 24124 15895 24176 15904
rect 24124 15861 24133 15895
rect 24133 15861 24167 15895
rect 24167 15861 24176 15895
rect 24124 15852 24176 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 11152 15648 11204 15700
rect 11428 15580 11480 15632
rect 11980 15648 12032 15700
rect 12992 15648 13044 15700
rect 13912 15648 13964 15700
rect 15844 15648 15896 15700
rect 16304 15691 16356 15700
rect 16304 15657 16313 15691
rect 16313 15657 16347 15691
rect 16347 15657 16356 15691
rect 16304 15648 16356 15657
rect 16580 15648 16632 15700
rect 17132 15648 17184 15700
rect 18144 15648 18196 15700
rect 18788 15648 18840 15700
rect 18972 15691 19024 15700
rect 18972 15657 18981 15691
rect 18981 15657 19015 15691
rect 19015 15657 19024 15691
rect 18972 15648 19024 15657
rect 19248 15691 19300 15700
rect 19248 15657 19257 15691
rect 19257 15657 19291 15691
rect 19291 15657 19300 15691
rect 19248 15648 19300 15657
rect 20904 15691 20956 15700
rect 20904 15657 20913 15691
rect 20913 15657 20947 15691
rect 20947 15657 20956 15691
rect 20904 15648 20956 15657
rect 23020 15648 23072 15700
rect 24216 15648 24268 15700
rect 24584 15648 24636 15700
rect 13084 15580 13136 15632
rect 14188 15623 14240 15632
rect 14188 15589 14197 15623
rect 14197 15589 14231 15623
rect 14231 15589 14240 15623
rect 14188 15580 14240 15589
rect 15660 15580 15712 15632
rect 11336 15555 11388 15564
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 11336 15512 11388 15521
rect 13820 15512 13872 15564
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 17224 15512 17276 15564
rect 19616 15555 19668 15564
rect 19616 15521 19625 15555
rect 19625 15521 19659 15555
rect 19659 15521 19668 15555
rect 19616 15512 19668 15521
rect 21456 15580 21508 15632
rect 24952 15580 25004 15632
rect 20904 15512 20956 15564
rect 22560 15555 22612 15564
rect 22560 15521 22569 15555
rect 22569 15521 22603 15555
rect 22603 15521 22612 15555
rect 22560 15512 22612 15521
rect 22836 15555 22888 15564
rect 22836 15521 22870 15555
rect 22870 15521 22888 15555
rect 25044 15555 25096 15564
rect 22836 15512 22888 15521
rect 25044 15521 25053 15555
rect 25053 15521 25087 15555
rect 25087 15521 25096 15555
rect 25044 15512 25096 15521
rect 10968 15444 11020 15496
rect 15660 15444 15712 15496
rect 16028 15444 16080 15496
rect 19708 15487 19760 15496
rect 10784 15419 10836 15428
rect 10784 15385 10793 15419
rect 10793 15385 10827 15419
rect 10827 15385 10836 15419
rect 10784 15376 10836 15385
rect 15568 15376 15620 15428
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 20720 15444 20772 15496
rect 21824 15444 21876 15496
rect 12440 15308 12492 15360
rect 12808 15308 12860 15360
rect 16488 15308 16540 15360
rect 21456 15376 21508 15428
rect 16856 15308 16908 15360
rect 17132 15308 17184 15360
rect 18696 15351 18748 15360
rect 18696 15317 18705 15351
rect 18705 15317 18739 15351
rect 18739 15317 18748 15351
rect 18696 15308 18748 15317
rect 21916 15351 21968 15360
rect 21916 15317 21925 15351
rect 21925 15317 21959 15351
rect 21959 15317 21968 15351
rect 21916 15308 21968 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 10876 15104 10928 15156
rect 11060 15104 11112 15156
rect 9956 15011 10008 15020
rect 9956 14977 9965 15011
rect 9965 14977 9999 15011
rect 9999 14977 10008 15011
rect 9956 14968 10008 14977
rect 10784 14968 10836 15020
rect 11244 15011 11296 15020
rect 11244 14977 11253 15011
rect 11253 14977 11287 15011
rect 11287 14977 11296 15011
rect 11244 14968 11296 14977
rect 11336 15011 11388 15020
rect 11336 14977 11345 15011
rect 11345 14977 11379 15011
rect 11379 14977 11388 15011
rect 11336 14968 11388 14977
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 13820 15104 13872 15156
rect 17224 15104 17276 15156
rect 18788 15104 18840 15156
rect 21824 15147 21876 15156
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 22376 15147 22428 15156
rect 22376 15113 22385 15147
rect 22385 15113 22419 15147
rect 22419 15113 22428 15147
rect 22376 15104 22428 15113
rect 22836 15104 22888 15156
rect 14004 15036 14056 15088
rect 12716 14968 12768 15020
rect 13728 14968 13780 15020
rect 14372 14968 14424 15020
rect 14004 14943 14056 14952
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 14004 14900 14056 14909
rect 18696 14968 18748 15020
rect 24860 15104 24912 15156
rect 26240 15147 26292 15156
rect 26240 15113 26249 15147
rect 26249 15113 26283 15147
rect 26283 15113 26292 15147
rect 26240 15104 26292 15113
rect 25044 15079 25096 15088
rect 25044 15045 25053 15079
rect 25053 15045 25087 15079
rect 25087 15045 25096 15079
rect 25044 15036 25096 15045
rect 23940 14968 23992 15020
rect 19524 14900 19576 14952
rect 19892 14900 19944 14952
rect 22376 14900 22428 14952
rect 24124 14900 24176 14952
rect 14372 14832 14424 14884
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 11152 14764 11204 14773
rect 11244 14764 11296 14816
rect 12532 14764 12584 14816
rect 13912 14764 13964 14816
rect 18788 14832 18840 14884
rect 19616 14832 19668 14884
rect 19708 14875 19760 14884
rect 19708 14841 19717 14875
rect 19717 14841 19751 14875
rect 19751 14841 19760 14875
rect 19708 14832 19760 14841
rect 23020 14832 23072 14884
rect 15752 14764 15804 14816
rect 16488 14764 16540 14816
rect 16764 14807 16816 14816
rect 16764 14773 16773 14807
rect 16773 14773 16807 14807
rect 16807 14773 16816 14807
rect 16764 14764 16816 14773
rect 18236 14807 18288 14816
rect 18236 14773 18245 14807
rect 18245 14773 18279 14807
rect 18279 14773 18288 14807
rect 18236 14764 18288 14773
rect 23848 14764 23900 14816
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 24308 14764 24360 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 10784 14560 10836 14612
rect 12716 14603 12768 14612
rect 12716 14569 12725 14603
rect 12725 14569 12759 14603
rect 12759 14569 12768 14603
rect 12716 14560 12768 14569
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 14004 14560 14056 14612
rect 14832 14560 14884 14612
rect 16488 14560 16540 14612
rect 18512 14603 18564 14612
rect 18512 14569 18521 14603
rect 18521 14569 18555 14603
rect 18555 14569 18564 14603
rect 18512 14560 18564 14569
rect 20444 14560 20496 14612
rect 20720 14603 20772 14612
rect 20720 14569 20729 14603
rect 20729 14569 20763 14603
rect 20763 14569 20772 14603
rect 20720 14560 20772 14569
rect 20904 14603 20956 14612
rect 20904 14569 20913 14603
rect 20913 14569 20947 14603
rect 20947 14569 20956 14603
rect 20904 14560 20956 14569
rect 23940 14603 23992 14612
rect 23940 14569 23949 14603
rect 23949 14569 23983 14603
rect 23983 14569 23992 14603
rect 23940 14560 23992 14569
rect 25320 14560 25372 14612
rect 19984 14492 20036 14544
rect 10784 14424 10836 14476
rect 11980 14424 12032 14476
rect 14004 14467 14056 14476
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 15936 14467 15988 14476
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 17960 14424 18012 14476
rect 19432 14424 19484 14476
rect 21272 14467 21324 14476
rect 13636 14356 13688 14408
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 15292 14356 15344 14408
rect 16764 14356 16816 14408
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 21272 14433 21281 14467
rect 21281 14433 21315 14467
rect 21315 14433 21324 14467
rect 21272 14424 21324 14433
rect 22836 14467 22888 14476
rect 22836 14433 22870 14467
rect 22870 14433 22888 14467
rect 22836 14424 22888 14433
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 20260 14356 20312 14408
rect 20904 14356 20956 14408
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 15568 14331 15620 14340
rect 15568 14297 15577 14331
rect 15577 14297 15611 14331
rect 15611 14297 15620 14331
rect 15568 14288 15620 14297
rect 12072 14263 12124 14272
rect 12072 14229 12081 14263
rect 12081 14229 12115 14263
rect 12115 14229 12124 14263
rect 12072 14220 12124 14229
rect 14188 14220 14240 14272
rect 16488 14220 16540 14272
rect 16856 14263 16908 14272
rect 16856 14229 16865 14263
rect 16865 14229 16899 14263
rect 16899 14229 16908 14263
rect 16856 14220 16908 14229
rect 23940 14288 23992 14340
rect 24032 14220 24084 14272
rect 26056 14220 26108 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 10784 14016 10836 14068
rect 11336 14016 11388 14068
rect 13452 14016 13504 14068
rect 13728 14016 13780 14068
rect 14004 14016 14056 14068
rect 16948 14016 17000 14068
rect 17224 14016 17276 14068
rect 18512 14016 18564 14068
rect 12164 13880 12216 13932
rect 13728 13880 13780 13932
rect 10968 13812 11020 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 15200 13812 15252 13864
rect 16488 13880 16540 13932
rect 18696 14016 18748 14068
rect 19984 14016 20036 14068
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 22008 14059 22060 14068
rect 22008 14025 22017 14059
rect 22017 14025 22051 14059
rect 22051 14025 22060 14059
rect 22008 14016 22060 14025
rect 24768 14016 24820 14068
rect 26056 14059 26108 14068
rect 26056 14025 26065 14059
rect 26065 14025 26099 14059
rect 26099 14025 26108 14059
rect 26056 14016 26108 14025
rect 15476 13812 15528 13864
rect 15752 13812 15804 13864
rect 9772 13744 9824 13796
rect 14280 13787 14332 13796
rect 14280 13753 14289 13787
rect 14289 13753 14323 13787
rect 14323 13753 14332 13787
rect 14280 13744 14332 13753
rect 14740 13744 14792 13796
rect 14924 13744 14976 13796
rect 15384 13744 15436 13796
rect 10784 13719 10836 13728
rect 10784 13685 10793 13719
rect 10793 13685 10827 13719
rect 10827 13685 10836 13719
rect 10784 13676 10836 13685
rect 12900 13676 12952 13728
rect 18420 13812 18472 13864
rect 20812 13880 20864 13932
rect 21824 13923 21876 13932
rect 21824 13889 21833 13923
rect 21833 13889 21867 13923
rect 21867 13889 21876 13923
rect 21824 13880 21876 13889
rect 22836 13880 22888 13932
rect 19340 13812 19392 13864
rect 20444 13812 20496 13864
rect 20904 13855 20956 13864
rect 20904 13821 20913 13855
rect 20913 13821 20947 13855
rect 20947 13821 20956 13855
rect 20904 13812 20956 13821
rect 21272 13812 21324 13864
rect 22744 13812 22796 13864
rect 16672 13744 16724 13796
rect 21824 13744 21876 13796
rect 23940 13812 23992 13864
rect 24860 13812 24912 13864
rect 24768 13744 24820 13796
rect 16488 13719 16540 13728
rect 16488 13685 16497 13719
rect 16497 13685 16531 13719
rect 16531 13685 16540 13719
rect 16488 13676 16540 13685
rect 18512 13676 18564 13728
rect 21272 13676 21324 13728
rect 21640 13676 21692 13728
rect 22376 13719 22428 13728
rect 22376 13685 22385 13719
rect 22385 13685 22419 13719
rect 22419 13685 22428 13719
rect 22376 13676 22428 13685
rect 25136 13676 25188 13728
rect 26056 13676 26108 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 9772 13515 9824 13524
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 9956 13472 10008 13524
rect 10876 13472 10928 13524
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 14832 13472 14884 13524
rect 15108 13515 15160 13524
rect 15108 13481 15117 13515
rect 15117 13481 15151 13515
rect 15151 13481 15160 13515
rect 15108 13472 15160 13481
rect 19524 13472 19576 13524
rect 20260 13515 20312 13524
rect 20260 13481 20269 13515
rect 20269 13481 20303 13515
rect 20303 13481 20312 13515
rect 20260 13472 20312 13481
rect 24308 13472 24360 13524
rect 25044 13515 25096 13524
rect 25044 13481 25053 13515
rect 25053 13481 25087 13515
rect 25087 13481 25096 13515
rect 25044 13472 25096 13481
rect 11336 13404 11388 13456
rect 12072 13404 12124 13456
rect 16120 13404 16172 13456
rect 18236 13447 18288 13456
rect 18236 13413 18245 13447
rect 18245 13413 18279 13447
rect 18279 13413 18288 13447
rect 18236 13404 18288 13413
rect 19248 13404 19300 13456
rect 21456 13404 21508 13456
rect 23296 13404 23348 13456
rect 12900 13379 12952 13388
rect 12900 13345 12909 13379
rect 12909 13345 12943 13379
rect 12943 13345 12952 13379
rect 12900 13336 12952 13345
rect 14004 13379 14056 13388
rect 14004 13345 14013 13379
rect 14013 13345 14047 13379
rect 14047 13345 14056 13379
rect 14004 13336 14056 13345
rect 15384 13336 15436 13388
rect 19156 13336 19208 13388
rect 19616 13379 19668 13388
rect 19616 13345 19625 13379
rect 19625 13345 19659 13379
rect 19659 13345 19668 13379
rect 19616 13336 19668 13345
rect 21824 13336 21876 13388
rect 24032 13336 24084 13388
rect 24676 13336 24728 13388
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15108 13268 15160 13320
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18880 13268 18932 13320
rect 19524 13268 19576 13320
rect 19892 13311 19944 13320
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 21088 13268 21140 13320
rect 23112 13311 23164 13320
rect 15292 13200 15344 13252
rect 15936 13200 15988 13252
rect 17316 13243 17368 13252
rect 17316 13209 17325 13243
rect 17325 13209 17359 13243
rect 17359 13209 17368 13243
rect 17316 13200 17368 13209
rect 17592 13200 17644 13252
rect 20536 13200 20588 13252
rect 22376 13200 22428 13252
rect 23112 13277 23121 13311
rect 23121 13277 23155 13311
rect 23155 13277 23164 13311
rect 23112 13268 23164 13277
rect 24768 13268 24820 13320
rect 23756 13200 23808 13252
rect 11152 13132 11204 13184
rect 16396 13132 16448 13184
rect 17960 13132 18012 13184
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 22468 13175 22520 13184
rect 22468 13141 22477 13175
rect 22477 13141 22511 13175
rect 22511 13141 22520 13175
rect 22468 13132 22520 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 10968 12928 11020 12980
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 14096 12928 14148 12980
rect 19616 12928 19668 12980
rect 19984 12928 20036 12980
rect 21088 12928 21140 12980
rect 24860 12928 24912 12980
rect 25136 12928 25188 12980
rect 14740 12860 14792 12912
rect 16120 12860 16172 12912
rect 24032 12903 24084 12912
rect 24032 12869 24041 12903
rect 24041 12869 24075 12903
rect 24075 12869 24084 12903
rect 24032 12860 24084 12869
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 22192 12792 22244 12844
rect 24124 12835 24176 12844
rect 24124 12801 24133 12835
rect 24133 12801 24167 12835
rect 24167 12801 24176 12835
rect 24124 12792 24176 12801
rect 11980 12724 12032 12776
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 13820 12724 13872 12776
rect 14280 12724 14332 12776
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 18696 12767 18748 12776
rect 17868 12724 17920 12733
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 19064 12724 19116 12776
rect 20904 12724 20956 12776
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 22468 12724 22520 12776
rect 12072 12656 12124 12708
rect 13636 12656 13688 12708
rect 16488 12656 16540 12708
rect 18328 12656 18380 12708
rect 19892 12656 19944 12708
rect 19984 12656 20036 12708
rect 20260 12656 20312 12708
rect 23112 12699 23164 12708
rect 23112 12665 23121 12699
rect 23121 12665 23155 12699
rect 23155 12665 23164 12699
rect 23112 12656 23164 12665
rect 24952 12656 25004 12708
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 18512 12588 18564 12640
rect 18788 12588 18840 12640
rect 20536 12588 20588 12640
rect 21088 12588 21140 12640
rect 21824 12588 21876 12640
rect 22928 12588 22980 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 11336 12384 11388 12436
rect 11980 12384 12032 12436
rect 13820 12427 13872 12436
rect 13820 12393 13829 12427
rect 13829 12393 13863 12427
rect 13863 12393 13872 12427
rect 13820 12384 13872 12393
rect 15200 12384 15252 12436
rect 15384 12384 15436 12436
rect 15936 12384 15988 12436
rect 16488 12384 16540 12436
rect 16764 12427 16816 12436
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 18420 12384 18472 12436
rect 19064 12384 19116 12436
rect 19340 12384 19392 12436
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 22836 12427 22888 12436
rect 22836 12393 22845 12427
rect 22845 12393 22879 12427
rect 22879 12393 22888 12427
rect 22836 12384 22888 12393
rect 23296 12427 23348 12436
rect 23296 12393 23305 12427
rect 23305 12393 23339 12427
rect 23339 12393 23348 12427
rect 23296 12384 23348 12393
rect 23756 12384 23808 12436
rect 24952 12427 25004 12436
rect 11612 12316 11664 12368
rect 12164 12316 12216 12368
rect 16212 12316 16264 12368
rect 15844 12248 15896 12300
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 15108 12180 15160 12189
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 17776 12316 17828 12368
rect 18512 12316 18564 12368
rect 19432 12316 19484 12368
rect 21088 12316 21140 12368
rect 24952 12393 24961 12427
rect 24961 12393 24995 12427
rect 24995 12393 25004 12427
rect 24952 12384 25004 12393
rect 24124 12316 24176 12368
rect 25320 12316 25372 12368
rect 18880 12248 18932 12300
rect 20720 12248 20772 12300
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 22836 12248 22888 12300
rect 15936 12180 15988 12189
rect 17500 12180 17552 12232
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 16764 12112 16816 12164
rect 18512 12180 18564 12232
rect 19064 12180 19116 12232
rect 11888 12044 11940 12096
rect 12992 12044 13044 12096
rect 13820 12044 13872 12096
rect 17316 12044 17368 12096
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 18880 12044 18932 12096
rect 19156 12044 19208 12096
rect 20904 12044 20956 12096
rect 22192 12044 22244 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 11612 11883 11664 11892
rect 11612 11849 11621 11883
rect 11621 11849 11655 11883
rect 11655 11849 11664 11883
rect 11612 11840 11664 11849
rect 15476 11840 15528 11892
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 17684 11840 17736 11892
rect 13360 11704 13412 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 16764 11679 16816 11688
rect 16764 11645 16773 11679
rect 16773 11645 16807 11679
rect 16807 11645 16816 11679
rect 16764 11636 16816 11645
rect 17960 11636 18012 11688
rect 18420 11840 18472 11892
rect 21088 11840 21140 11892
rect 23756 11840 23808 11892
rect 25320 11883 25372 11892
rect 25320 11849 25329 11883
rect 25329 11849 25363 11883
rect 25363 11849 25372 11883
rect 25320 11840 25372 11849
rect 20536 11772 20588 11824
rect 23020 11772 23072 11824
rect 20720 11704 20772 11756
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 24584 11704 24636 11756
rect 24952 11747 25004 11756
rect 24952 11713 24961 11747
rect 24961 11713 24995 11747
rect 24995 11713 25004 11747
rect 24952 11704 25004 11713
rect 22192 11636 22244 11688
rect 13728 11611 13780 11620
rect 13728 11577 13737 11611
rect 13737 11577 13771 11611
rect 13771 11577 13780 11611
rect 13728 11568 13780 11577
rect 18696 11568 18748 11620
rect 24860 11568 24912 11620
rect 11888 11543 11940 11552
rect 11888 11509 11897 11543
rect 11897 11509 11931 11543
rect 11931 11509 11940 11543
rect 11888 11500 11940 11509
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 16304 11500 16356 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 17776 11543 17828 11552
rect 16856 11500 16908 11509
rect 17776 11509 17785 11543
rect 17785 11509 17819 11543
rect 17819 11509 17828 11543
rect 17776 11500 17828 11509
rect 19340 11500 19392 11552
rect 21732 11500 21784 11552
rect 23664 11500 23716 11552
rect 24216 11500 24268 11552
rect 24584 11500 24636 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 13728 11296 13780 11348
rect 14832 11296 14884 11348
rect 15936 11296 15988 11348
rect 16948 11296 17000 11348
rect 18236 11296 18288 11348
rect 19064 11296 19116 11348
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 20904 11339 20956 11348
rect 20904 11305 20913 11339
rect 20913 11305 20947 11339
rect 20947 11305 20956 11339
rect 20904 11296 20956 11305
rect 21456 11296 21508 11348
rect 22008 11296 22060 11348
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 22836 11296 22888 11348
rect 23756 11296 23808 11348
rect 24952 11296 25004 11348
rect 25688 11296 25740 11348
rect 11888 11160 11940 11212
rect 15384 11228 15436 11280
rect 16028 11228 16080 11280
rect 20168 11228 20220 11280
rect 12716 11203 12768 11212
rect 12716 11169 12750 11203
rect 12750 11169 12768 11203
rect 12716 11160 12768 11169
rect 13820 11160 13872 11212
rect 16488 11160 16540 11212
rect 17316 11203 17368 11212
rect 17316 11169 17350 11203
rect 17350 11169 17368 11203
rect 17316 11160 17368 11169
rect 19340 11160 19392 11212
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 16948 11092 17000 11144
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 22652 11160 22704 11212
rect 23020 11228 23072 11280
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 10968 11024 11020 11076
rect 11704 11024 11756 11076
rect 11888 10999 11940 11008
rect 11888 10965 11897 10999
rect 11897 10965 11931 10999
rect 11931 10965 11940 10999
rect 11888 10956 11940 10965
rect 12348 10999 12400 11008
rect 12348 10965 12357 10999
rect 12357 10965 12391 10999
rect 12391 10965 12400 10999
rect 12348 10956 12400 10965
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 18512 11024 18564 11076
rect 14004 10956 14056 11008
rect 19340 10956 19392 11008
rect 19892 10956 19944 11008
rect 21640 10956 21692 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 16028 10752 16080 10804
rect 17316 10752 17368 10804
rect 17684 10752 17736 10804
rect 11428 10659 11480 10668
rect 11428 10625 11437 10659
rect 11437 10625 11471 10659
rect 11471 10625 11480 10659
rect 11428 10616 11480 10625
rect 11060 10548 11112 10600
rect 16580 10684 16632 10736
rect 12348 10616 12400 10668
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 10876 10412 10928 10464
rect 11796 10455 11848 10464
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 13452 10412 13504 10464
rect 14556 10616 14608 10668
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 16120 10616 16172 10668
rect 16672 10616 16724 10668
rect 16856 10548 16908 10600
rect 18052 10548 18104 10600
rect 19156 10752 19208 10804
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 19708 10795 19760 10804
rect 19708 10761 19717 10795
rect 19717 10761 19751 10795
rect 19751 10761 19760 10795
rect 19708 10752 19760 10761
rect 23204 10752 23256 10804
rect 21364 10684 21416 10736
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 15844 10480 15896 10532
rect 16396 10480 16448 10532
rect 18696 10480 18748 10532
rect 14004 10412 14056 10464
rect 14832 10412 14884 10464
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 19432 10616 19484 10668
rect 19892 10591 19944 10600
rect 19892 10557 19901 10591
rect 19901 10557 19935 10591
rect 19935 10557 19944 10591
rect 19892 10548 19944 10557
rect 21640 10659 21692 10668
rect 21640 10625 21649 10659
rect 21649 10625 21683 10659
rect 21683 10625 21692 10659
rect 21640 10616 21692 10625
rect 22100 10616 22152 10668
rect 23940 10752 23992 10804
rect 25228 10752 25280 10804
rect 25320 10752 25372 10804
rect 24308 10659 24360 10668
rect 24308 10625 24317 10659
rect 24317 10625 24351 10659
rect 24351 10625 24360 10659
rect 24308 10616 24360 10625
rect 24860 10616 24912 10668
rect 19340 10412 19392 10464
rect 20444 10412 20496 10464
rect 21180 10412 21232 10464
rect 21456 10412 21508 10464
rect 24216 10548 24268 10600
rect 23112 10480 23164 10532
rect 23296 10480 23348 10532
rect 22836 10412 22888 10464
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 23664 10412 23716 10464
rect 24216 10455 24268 10464
rect 24216 10421 24225 10455
rect 24225 10421 24259 10455
rect 24259 10421 24268 10455
rect 24216 10412 24268 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 11428 10208 11480 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 14740 10251 14792 10260
rect 14740 10217 14749 10251
rect 14749 10217 14783 10251
rect 14783 10217 14792 10251
rect 14740 10208 14792 10217
rect 16028 10208 16080 10260
rect 16212 10208 16264 10260
rect 16580 10208 16632 10260
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 18236 10251 18288 10260
rect 18236 10217 18245 10251
rect 18245 10217 18279 10251
rect 18279 10217 18288 10251
rect 18236 10208 18288 10217
rect 18972 10208 19024 10260
rect 20168 10208 20220 10260
rect 21088 10208 21140 10260
rect 21272 10208 21324 10260
rect 21548 10208 21600 10260
rect 22008 10208 22060 10260
rect 22652 10208 22704 10260
rect 22928 10251 22980 10260
rect 11244 10004 11296 10056
rect 11888 10140 11940 10192
rect 14648 10140 14700 10192
rect 17500 10140 17552 10192
rect 22928 10217 22937 10251
rect 22937 10217 22971 10251
rect 22971 10217 22980 10251
rect 22928 10208 22980 10217
rect 23848 10251 23900 10260
rect 23848 10217 23857 10251
rect 23857 10217 23891 10251
rect 23891 10217 23900 10251
rect 23848 10208 23900 10217
rect 24216 10208 24268 10260
rect 24308 10208 24360 10260
rect 12348 10072 12400 10124
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 16028 10115 16080 10124
rect 16028 10081 16037 10115
rect 16037 10081 16071 10115
rect 16071 10081 16080 10115
rect 16028 10072 16080 10081
rect 19248 10072 19300 10124
rect 19984 10072 20036 10124
rect 21088 10072 21140 10124
rect 21456 10072 21508 10124
rect 24952 10072 25004 10124
rect 16672 10004 16724 10056
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 16580 9936 16632 9988
rect 20076 10004 20128 10056
rect 21640 10004 21692 10056
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 13820 9868 13872 9920
rect 14188 9868 14240 9920
rect 15844 9868 15896 9920
rect 16948 9868 17000 9920
rect 17684 9868 17736 9920
rect 20628 9911 20680 9920
rect 20628 9877 20637 9911
rect 20637 9877 20671 9911
rect 20671 9877 20680 9911
rect 20628 9868 20680 9877
rect 20996 9868 21048 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 10876 9664 10928 9716
rect 11796 9528 11848 9580
rect 10140 9392 10192 9444
rect 10600 9392 10652 9444
rect 13084 9664 13136 9716
rect 12808 9528 12860 9580
rect 13176 9596 13228 9648
rect 16212 9664 16264 9716
rect 17316 9664 17368 9716
rect 20168 9664 20220 9716
rect 19432 9639 19484 9648
rect 19432 9605 19441 9639
rect 19441 9605 19475 9639
rect 19475 9605 19484 9639
rect 19432 9596 19484 9605
rect 21548 9664 21600 9716
rect 21640 9664 21692 9716
rect 22652 9707 22704 9716
rect 22652 9673 22661 9707
rect 22661 9673 22695 9707
rect 22695 9673 22704 9707
rect 22652 9664 22704 9673
rect 22836 9664 22888 9716
rect 23848 9707 23900 9716
rect 13268 9528 13320 9580
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 16396 9528 16448 9580
rect 13176 9460 13228 9512
rect 16580 9528 16632 9580
rect 17776 9528 17828 9580
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 21088 9571 21140 9580
rect 21088 9537 21097 9571
rect 21097 9537 21131 9571
rect 21131 9537 21140 9571
rect 21088 9528 21140 9537
rect 21456 9528 21508 9580
rect 23848 9673 23857 9707
rect 23857 9673 23891 9707
rect 23891 9673 23900 9707
rect 23848 9664 23900 9673
rect 24952 9707 25004 9716
rect 24952 9673 24961 9707
rect 24961 9673 24995 9707
rect 24995 9673 25004 9707
rect 24952 9664 25004 9673
rect 24952 9528 25004 9580
rect 25412 9571 25464 9580
rect 25412 9537 25421 9571
rect 25421 9537 25455 9571
rect 25455 9537 25464 9571
rect 25412 9528 25464 9537
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 17868 9460 17920 9512
rect 17960 9460 18012 9512
rect 20628 9460 20680 9512
rect 23388 9460 23440 9512
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 12348 9324 12400 9376
rect 12532 9392 12584 9444
rect 15752 9392 15804 9444
rect 18236 9392 18288 9444
rect 23020 9435 23072 9444
rect 23020 9401 23029 9435
rect 23029 9401 23063 9435
rect 23063 9401 23072 9435
rect 23020 9392 23072 9401
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 15292 9324 15344 9376
rect 16028 9324 16080 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 20628 9324 20680 9376
rect 23480 9367 23532 9376
rect 23480 9333 23489 9367
rect 23489 9333 23523 9367
rect 23523 9333 23532 9367
rect 24216 9367 24268 9376
rect 23480 9324 23532 9333
rect 24216 9333 24225 9367
rect 24225 9333 24259 9367
rect 24259 9333 24268 9367
rect 24216 9324 24268 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 12348 9120 12400 9172
rect 12808 9120 12860 9172
rect 14096 9120 14148 9172
rect 15752 9120 15804 9172
rect 17868 9120 17920 9172
rect 19340 9120 19392 9172
rect 20076 9163 20128 9172
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 20168 9120 20220 9172
rect 20444 9120 20496 9172
rect 21180 9120 21232 9172
rect 21824 9120 21876 9172
rect 24032 9120 24084 9172
rect 16120 9052 16172 9104
rect 16672 9052 16724 9104
rect 22008 9052 22060 9104
rect 11428 8984 11480 9036
rect 16212 8984 16264 9036
rect 18328 9027 18380 9036
rect 18328 8993 18362 9027
rect 18362 8993 18380 9027
rect 20720 9027 20772 9036
rect 18328 8984 18380 8993
rect 20720 8993 20729 9027
rect 20729 8993 20763 9027
rect 20763 8993 20772 9027
rect 20720 8984 20772 8993
rect 20904 9027 20956 9036
rect 20904 8993 20913 9027
rect 20913 8993 20947 9027
rect 20947 8993 20956 9027
rect 20904 8984 20956 8993
rect 20996 8984 21048 9036
rect 21640 8984 21692 9036
rect 23112 8984 23164 9036
rect 24768 8984 24820 9036
rect 10324 8916 10376 8968
rect 11244 8916 11296 8968
rect 14188 8916 14240 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 17684 8916 17736 8968
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 20076 8916 20128 8968
rect 20260 8916 20312 8968
rect 14096 8848 14148 8900
rect 14556 8848 14608 8900
rect 23940 8848 23992 8900
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 11428 8780 11480 8789
rect 15476 8780 15528 8832
rect 15752 8780 15804 8832
rect 16488 8780 16540 8832
rect 17960 8823 18012 8832
rect 17960 8789 17969 8823
rect 17969 8789 18003 8823
rect 18003 8789 18012 8823
rect 17960 8780 18012 8789
rect 20260 8780 20312 8832
rect 22284 8823 22336 8832
rect 22284 8789 22293 8823
rect 22293 8789 22327 8823
rect 22327 8789 22336 8823
rect 22284 8780 22336 8789
rect 23388 8823 23440 8832
rect 23388 8789 23397 8823
rect 23397 8789 23431 8823
rect 23431 8789 23440 8823
rect 23388 8780 23440 8789
rect 23848 8823 23900 8832
rect 23848 8789 23857 8823
rect 23857 8789 23891 8823
rect 23891 8789 23900 8823
rect 23848 8780 23900 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 10324 8619 10376 8628
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 12532 8619 12584 8628
rect 12532 8585 12541 8619
rect 12541 8585 12575 8619
rect 12575 8585 12584 8619
rect 12532 8576 12584 8585
rect 13084 8576 13136 8628
rect 13268 8576 13320 8628
rect 16120 8619 16172 8628
rect 16120 8585 16129 8619
rect 16129 8585 16163 8619
rect 16163 8585 16172 8619
rect 16120 8576 16172 8585
rect 16212 8576 16264 8628
rect 17592 8576 17644 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 20812 8576 20864 8628
rect 23112 8619 23164 8628
rect 23112 8585 23121 8619
rect 23121 8585 23155 8619
rect 23155 8585 23164 8619
rect 23112 8576 23164 8585
rect 24032 8576 24084 8628
rect 24952 8576 25004 8628
rect 12900 8508 12952 8560
rect 15936 8508 15988 8560
rect 11428 8483 11480 8492
rect 11428 8449 11437 8483
rect 11437 8449 11471 8483
rect 11471 8449 11480 8483
rect 11428 8440 11480 8449
rect 12532 8440 12584 8492
rect 11336 8372 11388 8424
rect 13268 8372 13320 8424
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 14740 8372 14792 8424
rect 12624 8304 12676 8356
rect 12900 8347 12952 8356
rect 12900 8313 12909 8347
rect 12909 8313 12943 8347
rect 12943 8313 12952 8347
rect 12900 8304 12952 8313
rect 16488 8304 16540 8356
rect 21088 8372 21140 8424
rect 22284 8440 22336 8492
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 22560 8372 22612 8424
rect 23388 8372 23440 8424
rect 20260 8304 20312 8356
rect 10876 8236 10928 8288
rect 11980 8236 12032 8288
rect 17040 8236 17092 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 20444 8236 20496 8288
rect 24124 8347 24176 8356
rect 24124 8313 24158 8347
rect 24158 8313 24176 8347
rect 24124 8304 24176 8313
rect 20996 8279 21048 8288
rect 20996 8245 21005 8279
rect 21005 8245 21039 8279
rect 21039 8245 21048 8279
rect 20996 8236 21048 8245
rect 21456 8279 21508 8288
rect 21456 8245 21465 8279
rect 21465 8245 21499 8279
rect 21499 8245 21508 8279
rect 21456 8236 21508 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 14280 8032 14332 8084
rect 16120 8032 16172 8084
rect 16488 8032 16540 8084
rect 17868 8032 17920 8084
rect 18052 8075 18104 8084
rect 18052 8041 18061 8075
rect 18061 8041 18095 8075
rect 18095 8041 18104 8075
rect 18052 8032 18104 8041
rect 18788 8032 18840 8084
rect 20720 8032 20772 8084
rect 22192 8032 22244 8084
rect 23940 8075 23992 8084
rect 23940 8041 23949 8075
rect 23949 8041 23983 8075
rect 23983 8041 23992 8075
rect 23940 8032 23992 8041
rect 24860 8032 24912 8084
rect 11152 7964 11204 8016
rect 14096 8007 14148 8016
rect 14096 7973 14105 8007
rect 14105 7973 14139 8007
rect 14139 7973 14148 8007
rect 14096 7964 14148 7973
rect 15108 7964 15160 8016
rect 15844 7964 15896 8016
rect 19248 8007 19300 8016
rect 19248 7973 19257 8007
rect 19257 7973 19291 8007
rect 19291 7973 19300 8007
rect 19248 7964 19300 7973
rect 21456 7964 21508 8016
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 11244 7896 11296 7948
rect 15568 7896 15620 7948
rect 18052 7896 18104 7948
rect 18604 7939 18656 7948
rect 18604 7905 18613 7939
rect 18613 7905 18647 7939
rect 18647 7905 18656 7939
rect 18604 7896 18656 7905
rect 22468 7896 22520 7948
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 14372 7828 14424 7880
rect 16396 7828 16448 7880
rect 18328 7760 18380 7812
rect 19432 7828 19484 7880
rect 20812 7828 20864 7880
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 22560 7871 22612 7880
rect 22560 7837 22569 7871
rect 22569 7837 22603 7871
rect 22603 7837 22612 7871
rect 22560 7828 22612 7837
rect 22100 7803 22152 7812
rect 22100 7769 22109 7803
rect 22109 7769 22143 7803
rect 22143 7769 22152 7803
rect 22100 7760 22152 7769
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 12900 7692 12952 7744
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 14004 7692 14056 7744
rect 15752 7692 15804 7744
rect 18512 7692 18564 7744
rect 20628 7692 20680 7744
rect 20904 7735 20956 7744
rect 20904 7701 20913 7735
rect 20913 7701 20947 7735
rect 20947 7701 20956 7735
rect 20904 7692 20956 7701
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 22744 7692 22796 7744
rect 24124 7692 24176 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 9864 7488 9916 7540
rect 11244 7531 11296 7540
rect 11244 7497 11253 7531
rect 11253 7497 11287 7531
rect 11287 7497 11296 7531
rect 11244 7488 11296 7497
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 14096 7531 14148 7540
rect 12440 7488 12492 7497
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 18604 7488 18656 7540
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 21824 7531 21876 7540
rect 21824 7497 21833 7531
rect 21833 7497 21867 7531
rect 21867 7497 21876 7531
rect 21824 7488 21876 7497
rect 22008 7488 22060 7540
rect 14372 7420 14424 7472
rect 15844 7420 15896 7472
rect 20352 7463 20404 7472
rect 20352 7429 20361 7463
rect 20361 7429 20395 7463
rect 20395 7429 20404 7463
rect 20352 7420 20404 7429
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 15752 7352 15804 7404
rect 8300 7284 8352 7336
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 10600 7284 10652 7336
rect 11060 7216 11112 7268
rect 11244 7284 11296 7336
rect 12072 7284 12124 7336
rect 12440 7284 12492 7336
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 17960 7284 18012 7336
rect 19248 7327 19300 7336
rect 16028 7216 16080 7268
rect 12072 7148 12124 7200
rect 14372 7191 14424 7200
rect 14372 7157 14381 7191
rect 14381 7157 14415 7191
rect 14415 7157 14424 7191
rect 14372 7148 14424 7157
rect 15292 7148 15344 7200
rect 16948 7191 17000 7200
rect 16948 7157 16957 7191
rect 16957 7157 16991 7191
rect 16991 7157 17000 7191
rect 16948 7148 17000 7157
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 18696 7148 18748 7200
rect 18880 7191 18932 7200
rect 18880 7157 18889 7191
rect 18889 7157 18923 7191
rect 18923 7157 18932 7191
rect 18880 7148 18932 7157
rect 19248 7293 19257 7327
rect 19257 7293 19291 7327
rect 19291 7293 19300 7327
rect 19248 7284 19300 7293
rect 19340 7284 19392 7336
rect 20628 7352 20680 7404
rect 20996 7352 21048 7404
rect 21456 7352 21508 7404
rect 22468 7352 22520 7404
rect 21916 7284 21968 7336
rect 22008 7284 22060 7336
rect 20720 7216 20772 7268
rect 21364 7216 21416 7268
rect 20076 7148 20128 7200
rect 22008 7191 22060 7200
rect 22008 7157 22017 7191
rect 22017 7157 22051 7191
rect 22051 7157 22060 7191
rect 22008 7148 22060 7157
rect 22376 7191 22428 7200
rect 22376 7157 22385 7191
rect 22385 7157 22419 7191
rect 22419 7157 22428 7191
rect 22376 7148 22428 7157
rect 22744 7148 22796 7200
rect 23940 7327 23992 7336
rect 23940 7293 23974 7327
rect 23974 7293 23992 7327
rect 23940 7284 23992 7293
rect 23204 7148 23256 7200
rect 23940 7148 23992 7200
rect 24124 7148 24176 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 12072 6987 12124 6996
rect 12072 6953 12081 6987
rect 12081 6953 12115 6987
rect 12115 6953 12124 6987
rect 12072 6944 12124 6953
rect 12256 6944 12308 6996
rect 14280 6987 14332 6996
rect 14280 6953 14289 6987
rect 14289 6953 14323 6987
rect 14323 6953 14332 6987
rect 14280 6944 14332 6953
rect 14556 6987 14608 6996
rect 14556 6953 14565 6987
rect 14565 6953 14599 6987
rect 14599 6953 14608 6987
rect 14556 6944 14608 6953
rect 15476 6944 15528 6996
rect 15752 6944 15804 6996
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 11888 6876 11940 6928
rect 9956 6851 10008 6860
rect 9956 6817 9990 6851
rect 9990 6817 10008 6851
rect 9956 6808 10008 6817
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 14004 6876 14056 6928
rect 14372 6876 14424 6928
rect 15384 6808 15436 6860
rect 15936 6808 15988 6860
rect 23204 6944 23256 6996
rect 18880 6876 18932 6928
rect 18144 6851 18196 6860
rect 18144 6817 18153 6851
rect 18153 6817 18187 6851
rect 18187 6817 18196 6851
rect 18144 6808 18196 6817
rect 18328 6808 18380 6860
rect 20720 6876 20772 6928
rect 21088 6808 21140 6860
rect 22100 6808 22152 6860
rect 23848 6851 23900 6860
rect 23848 6817 23857 6851
rect 23857 6817 23891 6851
rect 23891 6817 23900 6851
rect 23848 6808 23900 6817
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 20260 6740 20312 6792
rect 23296 6740 23348 6792
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 25044 6783 25096 6792
rect 24032 6740 24084 6749
rect 25044 6749 25053 6783
rect 25053 6749 25087 6783
rect 25087 6749 25096 6783
rect 25044 6740 25096 6749
rect 22560 6672 22612 6724
rect 9864 6604 9916 6656
rect 11152 6604 11204 6656
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 19340 6604 19392 6656
rect 23572 6604 23624 6656
rect 23940 6604 23992 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 572 6400 624 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 12256 6443 12308 6452
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 15936 6443 15988 6452
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 17500 6443 17552 6452
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 18328 6400 18380 6452
rect 21088 6443 21140 6452
rect 11060 6332 11112 6384
rect 12716 6375 12768 6384
rect 12716 6341 12725 6375
rect 12725 6341 12759 6375
rect 12759 6341 12768 6375
rect 12716 6332 12768 6341
rect 9956 6264 10008 6316
rect 11428 6307 11480 6316
rect 11428 6273 11437 6307
rect 11437 6273 11471 6307
rect 11471 6273 11480 6307
rect 11428 6264 11480 6273
rect 12624 6264 12676 6316
rect 14004 6307 14056 6316
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 15292 6264 15344 6316
rect 15568 6307 15620 6316
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 21088 6409 21097 6443
rect 21097 6409 21131 6443
rect 21131 6409 21140 6443
rect 21088 6400 21140 6409
rect 22192 6400 22244 6452
rect 23848 6400 23900 6452
rect 24032 6332 24084 6384
rect 23204 6264 23256 6316
rect 24584 6264 24636 6316
rect 9680 6196 9732 6248
rect 11612 6196 11664 6248
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 13728 6239 13780 6248
rect 13728 6205 13737 6239
rect 13737 6205 13771 6239
rect 13771 6205 13780 6239
rect 13728 6196 13780 6205
rect 10784 6128 10836 6180
rect 11336 6128 11388 6180
rect 8208 6060 8260 6112
rect 18880 6196 18932 6248
rect 17868 6128 17920 6180
rect 18236 6128 18288 6180
rect 20260 6196 20312 6248
rect 22100 6196 22152 6248
rect 24768 6196 24820 6248
rect 14004 6060 14056 6112
rect 14740 6103 14792 6112
rect 14740 6069 14749 6103
rect 14749 6069 14783 6103
rect 14783 6069 14792 6103
rect 14740 6060 14792 6069
rect 15384 6060 15436 6112
rect 15476 6060 15528 6112
rect 15752 6060 15804 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 18144 6103 18196 6112
rect 18144 6069 18153 6103
rect 18153 6069 18187 6103
rect 18187 6069 18196 6103
rect 18144 6060 18196 6069
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 19340 6060 19392 6112
rect 23388 6060 23440 6112
rect 24860 6060 24912 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 8208 5856 8260 5908
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 12348 5856 12400 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 13728 5856 13780 5908
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 15292 5856 15344 5908
rect 16488 5788 16540 5840
rect 18052 5856 18104 5908
rect 18328 5856 18380 5908
rect 20260 5899 20312 5908
rect 20260 5865 20269 5899
rect 20269 5865 20303 5899
rect 20303 5865 20312 5899
rect 20260 5856 20312 5865
rect 18420 5788 18472 5840
rect 11704 5720 11756 5772
rect 12072 5763 12124 5772
rect 12072 5729 12081 5763
rect 12081 5729 12115 5763
rect 12115 5729 12124 5763
rect 12072 5720 12124 5729
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12716 5652 12768 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 13820 5584 13872 5636
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 21456 5856 21508 5908
rect 23756 5856 23808 5908
rect 24584 5899 24636 5908
rect 24584 5865 24593 5899
rect 24593 5865 24627 5899
rect 24627 5865 24636 5899
rect 24584 5856 24636 5865
rect 21180 5788 21232 5840
rect 23296 5831 23348 5840
rect 23296 5797 23305 5831
rect 23305 5797 23339 5831
rect 23339 5797 23348 5831
rect 23296 5788 23348 5797
rect 23480 5788 23532 5840
rect 23940 5788 23992 5840
rect 25596 5720 25648 5772
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 23572 5652 23624 5704
rect 24032 5695 24084 5704
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 15568 5584 15620 5636
rect 13912 5516 13964 5568
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 23848 5516 23900 5568
rect 26148 5516 26200 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 12164 5312 12216 5364
rect 13728 5355 13780 5364
rect 13728 5321 13737 5355
rect 13737 5321 13771 5355
rect 13771 5321 13780 5355
rect 13728 5312 13780 5321
rect 14004 5355 14056 5364
rect 14004 5321 14013 5355
rect 14013 5321 14047 5355
rect 14047 5321 14056 5355
rect 14004 5312 14056 5321
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 23572 5312 23624 5364
rect 12072 5244 12124 5296
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 12808 5176 12860 5228
rect 11428 5040 11480 5092
rect 13360 5176 13412 5228
rect 24032 5312 24084 5364
rect 25596 5312 25648 5364
rect 18328 5176 18380 5228
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 20352 5219 20404 5228
rect 19616 5176 19668 5185
rect 13268 4972 13320 5024
rect 14832 5108 14884 5160
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 20352 5185 20361 5219
rect 20361 5185 20395 5219
rect 20395 5185 20404 5219
rect 20352 5176 20404 5185
rect 21180 5176 21232 5228
rect 23572 5176 23624 5228
rect 16856 5108 16908 5117
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 23848 5151 23900 5160
rect 18788 5040 18840 5092
rect 23848 5117 23857 5151
rect 23857 5117 23891 5151
rect 23891 5117 23900 5151
rect 23848 5108 23900 5117
rect 23204 5040 23256 5092
rect 24124 5083 24176 5092
rect 24124 5049 24158 5083
rect 24158 5049 24176 5083
rect 24124 5040 24176 5049
rect 15752 4972 15804 5024
rect 16764 4972 16816 5024
rect 17040 5015 17092 5024
rect 17040 4981 17049 5015
rect 17049 4981 17083 5015
rect 17083 4981 17092 5015
rect 17040 4972 17092 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 18696 5015 18748 5024
rect 18696 4981 18705 5015
rect 18705 4981 18739 5015
rect 18739 4981 18748 5015
rect 18696 4972 18748 4981
rect 19984 4972 20036 5024
rect 20260 5015 20312 5024
rect 20260 4981 20269 5015
rect 20269 4981 20303 5015
rect 20303 4981 20312 5015
rect 20260 4972 20312 4981
rect 21548 5015 21600 5024
rect 21548 4981 21557 5015
rect 21557 4981 21591 5015
rect 21591 4981 21600 5015
rect 21548 4972 21600 4981
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 24860 4972 24912 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 12164 4768 12216 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14096 4768 14148 4820
rect 14832 4811 14884 4820
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 15384 4768 15436 4820
rect 18604 4768 18656 4820
rect 20260 4768 20312 4820
rect 23112 4768 23164 4820
rect 23296 4768 23348 4820
rect 24676 4768 24728 4820
rect 24768 4768 24820 4820
rect 25044 4811 25096 4820
rect 25044 4777 25053 4811
rect 25053 4777 25087 4811
rect 25087 4777 25096 4811
rect 25044 4768 25096 4777
rect 12716 4700 12768 4752
rect 12808 4743 12860 4752
rect 12808 4709 12817 4743
rect 12817 4709 12851 4743
rect 12851 4709 12860 4743
rect 12808 4700 12860 4709
rect 16396 4700 16448 4752
rect 18420 4700 18472 4752
rect 18512 4700 18564 4752
rect 20168 4700 20220 4752
rect 23848 4700 23900 4752
rect 24952 4743 25004 4752
rect 24952 4709 24961 4743
rect 24961 4709 24995 4743
rect 24995 4709 25004 4743
rect 24952 4700 25004 4709
rect 14464 4632 14516 4684
rect 15292 4632 15344 4684
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 13360 4564 13412 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 16488 4564 16540 4616
rect 14280 4539 14332 4548
rect 14280 4505 14289 4539
rect 14289 4505 14323 4539
rect 14323 4505 14332 4539
rect 14280 4496 14332 4505
rect 22008 4632 22060 4684
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 18236 4564 18288 4616
rect 18972 4607 19024 4616
rect 18972 4573 18981 4607
rect 18981 4573 19015 4607
rect 19015 4573 19024 4607
rect 18972 4564 19024 4573
rect 19248 4564 19300 4616
rect 21456 4564 21508 4616
rect 23112 4564 23164 4616
rect 23572 4564 23624 4616
rect 24860 4564 24912 4616
rect 25136 4607 25188 4616
rect 25136 4573 25145 4607
rect 25145 4573 25179 4607
rect 25179 4573 25188 4607
rect 25136 4564 25188 4573
rect 16764 4471 16816 4480
rect 16764 4437 16773 4471
rect 16773 4437 16807 4471
rect 16807 4437 16816 4471
rect 16764 4428 16816 4437
rect 19524 4428 19576 4480
rect 20352 4428 20404 4480
rect 22100 4471 22152 4480
rect 22100 4437 22109 4471
rect 22109 4437 22143 4471
rect 22143 4437 22152 4471
rect 22560 4471 22612 4480
rect 22100 4428 22152 4437
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 22560 4428 22612 4437
rect 22836 4471 22888 4480
rect 22836 4437 22845 4471
rect 22845 4437 22879 4471
rect 22879 4437 22888 4471
rect 22836 4428 22888 4437
rect 24124 4471 24176 4480
rect 24124 4437 24133 4471
rect 24133 4437 24167 4471
rect 24167 4437 24176 4471
rect 24124 4428 24176 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 12808 4224 12860 4276
rect 13360 4267 13412 4276
rect 13360 4233 13369 4267
rect 13369 4233 13403 4267
rect 13403 4233 13412 4267
rect 13360 4224 13412 4233
rect 14096 4224 14148 4276
rect 15936 4267 15988 4276
rect 15936 4233 15945 4267
rect 15945 4233 15979 4267
rect 15979 4233 15988 4267
rect 15936 4224 15988 4233
rect 18236 4224 18288 4276
rect 18972 4267 19024 4276
rect 18972 4233 18981 4267
rect 18981 4233 19015 4267
rect 19015 4233 19024 4267
rect 18972 4224 19024 4233
rect 21456 4267 21508 4276
rect 21456 4233 21465 4267
rect 21465 4233 21499 4267
rect 21499 4233 21508 4267
rect 21456 4224 21508 4233
rect 22008 4224 22060 4276
rect 23296 4224 23348 4276
rect 24952 4224 25004 4276
rect 940 4156 992 4208
rect 9588 4156 9640 4208
rect 12900 4156 12952 4208
rect 14464 4156 14516 4208
rect 14924 4156 14976 4208
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 9128 4020 9180 4072
rect 9588 4020 9640 4072
rect 11336 4020 11388 4072
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 13636 4020 13688 4072
rect 17868 4088 17920 4140
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 22560 4088 22612 4097
rect 23572 4088 23624 4140
rect 18144 4063 18196 4072
rect 18144 4029 18153 4063
rect 18153 4029 18187 4063
rect 18187 4029 18196 4063
rect 18144 4020 18196 4029
rect 20168 4020 20220 4072
rect 21456 4020 21508 4072
rect 13820 3995 13872 4004
rect 13820 3961 13829 3995
rect 13829 3961 13863 3995
rect 13863 3961 13872 3995
rect 13820 3952 13872 3961
rect 16672 3995 16724 4004
rect 16672 3961 16681 3995
rect 16681 3961 16715 3995
rect 16715 3961 16724 3995
rect 16672 3952 16724 3961
rect 22100 3952 22152 4004
rect 22836 4020 22888 4072
rect 23756 4020 23808 4072
rect 23848 3952 23900 4004
rect 11152 3927 11204 3936
rect 11152 3893 11161 3927
rect 11161 3893 11195 3927
rect 11195 3893 11204 3927
rect 11152 3884 11204 3893
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 19524 3884 19576 3936
rect 20720 3884 20772 3936
rect 21916 3884 21968 3936
rect 22928 3884 22980 3936
rect 23756 3884 23808 3936
rect 25044 3927 25096 3936
rect 25044 3893 25053 3927
rect 25053 3893 25087 3927
rect 25087 3893 25096 3927
rect 25044 3884 25096 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 11520 3680 11572 3732
rect 12992 3723 13044 3732
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 13544 3680 13596 3732
rect 13912 3680 13964 3732
rect 15108 3680 15160 3732
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 18512 3680 18564 3732
rect 19248 3723 19300 3732
rect 19248 3689 19257 3723
rect 19257 3689 19291 3723
rect 19291 3689 19300 3723
rect 19248 3680 19300 3689
rect 19432 3680 19484 3732
rect 19984 3680 20036 3732
rect 22560 3680 22612 3732
rect 23848 3680 23900 3732
rect 24400 3723 24452 3732
rect 24400 3689 24409 3723
rect 24409 3689 24443 3723
rect 24443 3689 24452 3723
rect 24400 3680 24452 3689
rect 24952 3680 25004 3732
rect 25136 3680 25188 3732
rect 15568 3655 15620 3664
rect 15568 3621 15577 3655
rect 15577 3621 15611 3655
rect 15611 3621 15620 3655
rect 15568 3612 15620 3621
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 12532 3544 12584 3596
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 14464 3544 14516 3596
rect 20168 3612 20220 3664
rect 17316 3544 17368 3596
rect 22284 3612 22336 3664
rect 23940 3612 23992 3664
rect 24676 3612 24728 3664
rect 21824 3587 21876 3596
rect 21824 3553 21858 3587
rect 21858 3553 21876 3587
rect 21824 3544 21876 3553
rect 12348 3476 12400 3528
rect 14004 3519 14056 3528
rect 14004 3485 14013 3519
rect 14013 3485 14047 3519
rect 14047 3485 14056 3519
rect 14004 3476 14056 3485
rect 16764 3519 16816 3528
rect 11704 3340 11756 3392
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 13636 3340 13688 3392
rect 15384 3340 15436 3392
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 20720 3476 20772 3528
rect 24124 3408 24176 3460
rect 25044 3476 25096 3528
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 18512 3340 18564 3392
rect 23112 3340 23164 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12348 3136 12400 3188
rect 12532 3136 12584 3188
rect 14004 3136 14056 3188
rect 10876 3068 10928 3120
rect 11428 3111 11480 3120
rect 11428 3077 11437 3111
rect 11437 3077 11471 3111
rect 11471 3077 11480 3111
rect 11428 3068 11480 3077
rect 16948 3136 17000 3188
rect 18052 3179 18104 3188
rect 10784 2932 10836 2984
rect 11796 2932 11848 2984
rect 12164 2932 12216 2984
rect 12992 2932 13044 2984
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 19432 3136 19484 3188
rect 21824 3179 21876 3188
rect 21824 3145 21833 3179
rect 21833 3145 21867 3179
rect 21867 3145 21876 3179
rect 21824 3136 21876 3145
rect 22192 3136 22244 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 24124 3136 24176 3188
rect 24216 3136 24268 3188
rect 24676 3136 24728 3188
rect 25412 3136 25464 3188
rect 26884 3068 26936 3120
rect 18144 3000 18196 3052
rect 13268 2864 13320 2916
rect 18880 2932 18932 2984
rect 20168 2932 20220 2984
rect 20720 2975 20772 2984
rect 20720 2941 20754 2975
rect 20754 2941 20772 2975
rect 20720 2932 20772 2941
rect 23480 2932 23532 2984
rect 25412 2932 25464 2984
rect 23940 2907 23992 2916
rect 23940 2873 23949 2907
rect 23949 2873 23983 2907
rect 23983 2873 23992 2907
rect 23940 2864 23992 2873
rect 15384 2796 15436 2848
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 18512 2839 18564 2848
rect 18512 2805 18521 2839
rect 18521 2805 18555 2839
rect 18555 2805 18564 2839
rect 18512 2796 18564 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 12440 2592 12492 2644
rect 13728 2592 13780 2644
rect 15384 2592 15436 2644
rect 16304 2635 16356 2644
rect 16304 2601 16313 2635
rect 16313 2601 16347 2635
rect 16347 2601 16356 2635
rect 16304 2592 16356 2601
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19524 2592 19576 2644
rect 22008 2592 22060 2644
rect 22192 2635 22244 2644
rect 22192 2601 22201 2635
rect 22201 2601 22235 2635
rect 22235 2601 22244 2635
rect 22192 2592 22244 2601
rect 22284 2592 22336 2644
rect 23480 2592 23532 2644
rect 13268 2524 13320 2576
rect 11520 2456 11572 2508
rect 12532 2456 12584 2508
rect 14832 2456 14884 2508
rect 16120 2456 16172 2508
rect 18880 2524 18932 2576
rect 23204 2524 23256 2576
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 15660 2388 15712 2440
rect 16764 2431 16816 2440
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 17316 2388 17368 2440
rect 18144 2388 18196 2440
rect 20904 2499 20956 2508
rect 20904 2465 20913 2499
rect 20913 2465 20947 2499
rect 20947 2465 20956 2499
rect 20904 2456 20956 2465
rect 22744 2499 22796 2508
rect 22744 2465 22753 2499
rect 22753 2465 22787 2499
rect 22787 2465 22796 2499
rect 22744 2456 22796 2465
rect 23664 2456 23716 2508
rect 25320 2499 25372 2508
rect 25320 2465 25329 2499
rect 25329 2465 25363 2499
rect 25363 2465 25372 2499
rect 25320 2456 25372 2465
rect 20536 2388 20588 2440
rect 21640 2431 21692 2440
rect 21640 2397 21649 2431
rect 21649 2397 21683 2431
rect 21683 2397 21692 2431
rect 21640 2388 21692 2397
rect 22192 2388 22244 2440
rect 13728 2363 13780 2372
rect 13728 2329 13737 2363
rect 13737 2329 13771 2363
rect 13771 2329 13780 2363
rect 13728 2320 13780 2329
rect 21364 2320 21416 2372
rect 27528 2320 27580 2372
rect 10784 2252 10836 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 12532 2252 12584 2304
rect 13084 2252 13136 2304
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 16120 2295 16172 2304
rect 16120 2261 16129 2295
rect 16129 2261 16163 2295
rect 16163 2261 16172 2295
rect 16120 2252 16172 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 21548 552 21600 604
rect 24124 552 24176 604
<< metal2 >>
rect 294 27520 350 28000
rect 938 27520 994 28000
rect 1582 27520 1638 28000
rect 2318 27520 2374 28000
rect 2962 27520 3018 28000
rect 3698 27520 3754 28000
rect 4342 27520 4398 28000
rect 4986 27520 5042 28000
rect 5722 27520 5778 28000
rect 6366 27520 6422 28000
rect 7102 27520 7158 28000
rect 7746 27520 7802 28000
rect 8390 27520 8446 28000
rect 9126 27520 9182 28000
rect 9770 27520 9826 28000
rect 10506 27520 10562 28000
rect 11150 27520 11206 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13174 27520 13230 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15290 27520 15346 28000
rect 15934 27520 15990 28000
rect 16578 27520 16634 28000
rect 17314 27520 17370 28000
rect 17958 27520 18014 28000
rect 18694 27520 18750 28000
rect 19338 27520 19394 28000
rect 20074 27520 20130 28000
rect 20718 27520 20774 28000
rect 21362 27520 21418 28000
rect 22098 27520 22154 28000
rect 22742 27520 22798 28000
rect 23478 27520 23534 28000
rect 24122 27520 24178 28000
rect 24582 27704 24638 27713
rect 24582 27639 24638 27648
rect 308 27418 336 27520
rect 308 27390 428 27418
rect 400 15473 428 27390
rect 952 23089 980 27520
rect 938 23080 994 23089
rect 938 23015 994 23024
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 386 15464 442 15473
rect 386 15399 442 15408
rect 294 7440 350 7449
rect 294 7375 350 7384
rect 308 480 336 7375
rect 570 7032 626 7041
rect 570 6967 626 6976
rect 584 6458 612 6967
rect 572 6452 624 6458
rect 572 6394 624 6400
rect 940 4208 992 4214
rect 940 4150 992 4156
rect 952 480 980 4150
rect 1412 4049 1440 22034
rect 1596 19281 1624 27520
rect 2332 22098 2360 27520
rect 2976 22545 3004 27520
rect 2962 22536 3018 22545
rect 2962 22471 3018 22480
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 3712 19961 3740 27520
rect 4066 21040 4122 21049
rect 4066 20975 4122 20984
rect 3698 19952 3754 19961
rect 3698 19887 3754 19896
rect 1582 19272 1638 19281
rect 1582 19207 1638 19216
rect 4080 13977 4108 20975
rect 4356 19009 4384 27520
rect 5000 22681 5028 27520
rect 5736 25242 5764 27520
rect 5736 25214 6040 25242
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 4986 22672 5042 22681
rect 4986 22607 5042 22616
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 20097 6040 25214
rect 6380 23497 6408 27520
rect 7116 23633 7144 27520
rect 7760 24313 7788 27520
rect 7746 24304 7802 24313
rect 7746 24239 7802 24248
rect 7102 23624 7158 23633
rect 7102 23559 7158 23568
rect 6366 23488 6422 23497
rect 6366 23423 6422 23432
rect 7746 23488 7802 23497
rect 7746 23423 7802 23432
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 20398 7696 20742
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 5998 20088 6054 20097
rect 5998 20023 6054 20032
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 7564 19304 7616 19310
rect 7668 19292 7696 20334
rect 7760 19922 7788 23423
rect 8404 21690 8432 27520
rect 9140 24721 9168 27520
rect 9126 24712 9182 24721
rect 9126 24647 9182 24656
rect 9784 24041 9812 27520
rect 10520 27418 10548 27520
rect 10520 27390 10916 27418
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10690 24304 10746 24313
rect 10690 24239 10746 24248
rect 9770 24032 9826 24041
rect 9770 23967 9826 23976
rect 9310 23624 9366 23633
rect 9310 23559 9366 23568
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 9324 21350 9352 23559
rect 10704 23526 10732 24239
rect 10782 24168 10838 24177
rect 10782 24103 10838 24112
rect 10796 23866 10824 24103
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10888 22273 10916 27390
rect 11164 23662 11192 27520
rect 11900 24313 11928 27520
rect 11886 24304 11942 24313
rect 11886 24239 11942 24248
rect 12544 24154 12572 27520
rect 12714 24848 12770 24857
rect 13188 24834 13216 27520
rect 12714 24783 12770 24792
rect 13004 24806 13216 24834
rect 12728 24614 12756 24783
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12544 24126 12664 24154
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 11348 23730 11376 24006
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 11164 23474 11192 23598
rect 10980 23446 11192 23474
rect 11244 23520 11296 23526
rect 11244 23462 11296 23468
rect 10980 23322 11008 23446
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 11152 23248 11204 23254
rect 11256 23225 11284 23462
rect 12544 23322 12572 24006
rect 12636 23769 12664 24126
rect 12622 23760 12678 23769
rect 12622 23695 12678 23704
rect 12728 23610 12756 24210
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12636 23582 12756 23610
rect 12636 23526 12664 23582
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 11152 23190 11204 23196
rect 11242 23216 11298 23225
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11072 22642 11100 23054
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10874 22264 10930 22273
rect 10874 22199 10930 22208
rect 11072 22098 11100 22578
rect 11164 22438 11192 23190
rect 11242 23151 11298 23160
rect 12346 22672 12402 22681
rect 12164 22636 12216 22642
rect 12346 22607 12402 22616
rect 12164 22578 12216 22584
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 11886 22400 11942 22409
rect 11164 22234 11192 22374
rect 11886 22335 11942 22344
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21554 9996 21830
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9312 21344 9364 21350
rect 9312 21286 9364 21292
rect 9232 21049 9260 21286
rect 9218 21040 9274 21049
rect 9218 20975 9274 20984
rect 9324 20806 9352 21286
rect 9968 21010 9996 21490
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 7838 20360 7894 20369
rect 7838 20295 7840 20304
rect 7892 20295 7894 20304
rect 7840 20266 7892 20272
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 7838 20088 7894 20097
rect 7838 20023 7840 20032
rect 7892 20023 7894 20032
rect 7840 19994 7892 20000
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7616 19264 7696 19292
rect 7564 19246 7616 19252
rect 7760 19224 7788 19858
rect 7852 19514 7880 19994
rect 8036 19854 8064 20198
rect 8024 19848 8076 19854
rect 9324 19825 9352 20742
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9692 19922 9720 20538
rect 9968 20262 9996 20946
rect 10060 20942 10088 22034
rect 11164 21554 11192 22170
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 10060 20602 10088 20878
rect 10704 20602 10732 21354
rect 11256 21350 11284 21830
rect 11808 21690 11836 22034
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 9968 20058 9996 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 8024 19790 8076 19796
rect 9310 19816 9366 19825
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 8036 19292 8064 19790
rect 9310 19751 9366 19760
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8116 19304 8168 19310
rect 8036 19264 8116 19292
rect 7840 19236 7892 19242
rect 7760 19196 7840 19224
rect 4342 19000 4398 19009
rect 4342 18935 4398 18944
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 7760 15994 7788 19196
rect 7840 19178 7892 19184
rect 8036 18970 8064 19264
rect 8116 19246 8168 19252
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8220 17898 8248 19654
rect 9692 19360 9720 19858
rect 9968 19514 9996 19858
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9600 19332 9720 19360
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8404 18970 8432 19178
rect 9404 19168 9456 19174
rect 9310 19136 9366 19145
rect 9600 19145 9628 19332
rect 9404 19110 9456 19116
rect 9586 19136 9642 19145
rect 9310 19071 9366 19080
rect 9324 18970 9352 19071
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 8404 18834 8432 18906
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8772 18290 8800 18770
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 9416 18222 9444 19110
rect 9586 19071 9642 19080
rect 9680 18760 9732 18766
rect 9508 18708 9680 18714
rect 9508 18702 9732 18708
rect 9508 18686 9720 18702
rect 9968 18698 9996 19450
rect 10598 19272 10654 19281
rect 10598 19207 10600 19216
rect 10652 19207 10654 19216
rect 10600 19178 10652 19184
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10138 19000 10194 19009
rect 10289 18992 10585 19012
rect 10138 18935 10194 18944
rect 10152 18902 10180 18935
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9956 18692 10008 18698
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 8220 17882 8340 17898
rect 8220 17876 8352 17882
rect 8220 17870 8300 17876
rect 8300 17818 8352 17824
rect 9416 17542 9444 18158
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9416 17270 9444 17478
rect 9508 17338 9536 18686
rect 9956 18634 10008 18640
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9692 17882 9720 18566
rect 9968 18426 9996 18634
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9416 16794 9444 17206
rect 9600 17202 9628 17818
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9494 17096 9550 17105
rect 9494 17031 9496 17040
rect 9548 17031 9550 17040
rect 9496 17002 9548 17008
rect 9968 16980 9996 17614
rect 10060 17610 10088 18770
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10152 18290 10180 18702
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10520 17338 10548 17682
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10704 17134 10732 17818
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10048 16992 10100 16998
rect 9968 16952 10048 16980
rect 10048 16934 10100 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 10060 16017 10088 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 7576 15966 7788 15994
rect 10046 16008 10102 16017
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 4066 13968 4122 13977
rect 4066 13903 4122 13912
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 7576 12322 7604 15966
rect 10046 15943 10102 15952
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15026 9996 15846
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9784 13530 9812 13738
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9968 12986 9996 13466
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 7576 12294 7696 12322
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 3698 8392 3754 8401
rect 3698 8327 3754 8336
rect 2318 5672 2374 5681
rect 2318 5607 2374 5616
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1582 2544 1638 2553
rect 1582 2479 1638 2488
rect 1596 480 1624 2479
rect 2332 480 2360 5607
rect 2962 5264 3018 5273
rect 2962 5199 3018 5208
rect 2976 480 3004 5199
rect 3712 480 3740 8327
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4342 6760 4398 6769
rect 4342 6695 4398 6704
rect 4356 480 4384 6695
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 7668 5137 7696 12294
rect 7746 11112 7802 11121
rect 7746 11047 7802 11056
rect 7654 5128 7710 5137
rect 7654 5063 7710 5072
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6366 3904 6422 3913
rect 6366 3839 6422 3848
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 4986 3088 5042 3097
rect 4986 3023 5042 3032
rect 5000 480 5028 3023
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5722 1456 5778 1465
rect 5722 1391 5778 1400
rect 5736 480 5764 1391
rect 6380 480 6408 3839
rect 7102 3632 7158 3641
rect 7102 3567 7158 3576
rect 7116 480 7144 3567
rect 7760 480 7788 11047
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9876 7857 9904 7890
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9876 7546 9904 7783
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5930 8248 6054
rect 8312 5930 8340 7278
rect 9876 6662 9904 7278
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9968 6322 9996 6802
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 8220 5914 8340 5930
rect 8208 5908 8340 5914
rect 8260 5902 8340 5908
rect 8208 5850 8260 5856
rect 9588 4208 9640 4214
rect 9586 4176 9588 4185
rect 9640 4176 9642 4185
rect 9586 4111 9642 4120
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9588 4072 9640 4078
rect 9692 4060 9720 6190
rect 9968 5914 9996 6258
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9770 5536 9826 5545
rect 9770 5471 9826 5480
rect 9640 4032 9720 4060
rect 9588 4014 9640 4020
rect 8390 2952 8446 2961
rect 8390 2887 8446 2896
rect 8404 480 8432 2887
rect 9140 480 9168 4014
rect 9784 480 9812 5471
rect 10060 3913 10088 15943
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10796 15552 10824 20198
rect 10980 19938 11008 21286
rect 11256 21146 11284 21286
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11808 20874 11836 21626
rect 11796 20868 11848 20874
rect 11796 20810 11848 20816
rect 11808 20602 11836 20810
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11242 20496 11298 20505
rect 11242 20431 11298 20440
rect 11256 20262 11284 20431
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11900 19938 11928 22335
rect 12176 21690 12204 22578
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12360 21185 12388 22607
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12346 21176 12402 21185
rect 12346 21111 12402 21120
rect 12438 21040 12494 21049
rect 12438 20975 12440 20984
rect 12492 20975 12494 20984
rect 12440 20946 12492 20952
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 10980 19922 11100 19938
rect 10980 19916 11112 19922
rect 10980 19910 11060 19916
rect 11060 19858 11112 19864
rect 11716 19910 11928 19938
rect 12176 19922 12204 20334
rect 12348 20324 12400 20330
rect 12544 20312 12572 21286
rect 12400 20284 12572 20312
rect 12348 20266 12400 20272
rect 12636 20058 12664 23462
rect 12728 22642 12756 23462
rect 12820 23254 12848 24006
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12820 22778 12848 23190
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12728 22234 12756 22578
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12714 21584 12770 21593
rect 12714 21519 12770 21528
rect 12728 20466 12756 21519
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12164 19916 12216 19922
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 10888 17882 10916 19110
rect 11164 18902 11192 19110
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11440 18426 11468 18770
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 10966 18320 11022 18329
rect 10966 18255 11022 18264
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10980 17202 11008 18255
rect 11610 18184 11666 18193
rect 11610 18119 11666 18128
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11440 16658 11468 17206
rect 11428 16652 11480 16658
rect 11348 16612 11428 16640
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11164 15910 11192 15982
rect 11152 15904 11204 15910
rect 10874 15872 10930 15881
rect 11152 15846 11204 15852
rect 10874 15807 10930 15816
rect 10704 15524 10824 15552
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10232 14408 10284 14414
rect 10230 14376 10232 14385
rect 10284 14376 10286 14385
rect 10230 14311 10286 14320
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12458 10732 15524
rect 10782 15464 10838 15473
rect 10782 15399 10784 15408
rect 10836 15399 10838 15408
rect 10784 15370 10836 15376
rect 10782 15192 10838 15201
rect 10888 15162 10916 15807
rect 11164 15706 11192 15846
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11348 15570 11376 16612
rect 11428 16594 11480 16600
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11440 16114 11468 16390
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11440 15638 11468 16050
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11242 15464 11298 15473
rect 10782 15127 10838 15136
rect 10876 15156 10928 15162
rect 10796 15026 10824 15127
rect 10980 15144 11008 15438
rect 11242 15399 11298 15408
rect 11060 15156 11112 15162
rect 10980 15116 11060 15144
rect 10876 15098 10928 15104
rect 11060 15098 11112 15104
rect 11256 15026 11284 15399
rect 11348 15201 11376 15506
rect 11624 15314 11652 18119
rect 11716 16776 11744 19910
rect 12164 19858 12216 19864
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11900 19514 11928 19722
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11808 18834 11836 18906
rect 11900 18902 11928 19450
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11900 18426 11928 18838
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11716 16748 11836 16776
rect 11702 16688 11758 16697
rect 11702 16623 11704 16632
rect 11756 16623 11758 16632
rect 11704 16594 11756 16600
rect 11716 16250 11744 16594
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11440 15286 11652 15314
rect 11334 15192 11390 15201
rect 11334 15127 11390 15136
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 10796 14618 10824 14962
rect 11256 14822 11284 14962
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 10784 14612 10836 14618
rect 10836 14572 10916 14600
rect 10784 14554 10836 14560
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10796 14074 10824 14418
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10796 12889 10824 13670
rect 10888 13530 10916 14572
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10980 12986 11008 13806
rect 11164 13190 11192 14758
rect 11348 14074 11376 14962
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10782 12880 10838 12889
rect 11348 12850 11376 13398
rect 10782 12815 10838 12824
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 10704 12430 10824 12458
rect 11348 12442 11376 12786
rect 10796 11744 10824 12430
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 10704 11716 10824 11744
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10248 10732 11716
rect 10782 11656 10838 11665
rect 10782 11591 10838 11600
rect 10796 10810 10824 11591
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10980 10690 11008 11018
rect 11440 10826 11468 15286
rect 11808 12458 11836 16748
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15706 12020 15846
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11992 14482 12020 15642
rect 12084 15586 12112 19110
rect 12268 18714 12296 19654
rect 12636 19378 12664 19994
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12176 18686 12296 18714
rect 12176 17814 12204 18686
rect 12254 18592 12310 18601
rect 12254 18527 12310 18536
rect 12268 18426 12296 18527
rect 12360 18426 12388 18838
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12268 17134 12296 18362
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12360 17882 12388 18090
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16130 12480 16934
rect 12636 16833 12664 19314
rect 12820 19174 12848 19790
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 17338 12756 17614
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12820 17116 12848 19110
rect 12912 18193 12940 24550
rect 12898 18184 12954 18193
rect 12898 18119 12954 18128
rect 12900 17128 12952 17134
rect 12820 17096 12900 17116
rect 12952 17096 12954 17105
rect 12820 17088 12898 17096
rect 12898 17031 12954 17040
rect 13004 16998 13032 24806
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 13096 23322 13124 23598
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 13188 22658 13216 24686
rect 13268 24200 13320 24206
rect 13266 24168 13268 24177
rect 13360 24200 13412 24206
rect 13320 24168 13322 24177
rect 13360 24142 13412 24148
rect 13266 24103 13322 24112
rect 13280 23322 13308 24103
rect 13372 23526 13400 24142
rect 13924 23866 13952 27520
rect 14568 24857 14596 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14554 24848 14610 24857
rect 14554 24783 14610 24792
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14922 24712 14978 24721
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13280 22778 13308 23054
rect 13372 22982 13400 23462
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13832 23066 13860 23122
rect 13740 23038 13860 23066
rect 14094 23080 14150 23089
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13188 22630 13308 22658
rect 13176 22228 13228 22234
rect 13176 22170 13228 22176
rect 13188 21078 13216 22170
rect 13176 21072 13228 21078
rect 13176 21014 13228 21020
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17202 13216 17478
rect 13280 17252 13308 22630
rect 13372 22386 13400 22918
rect 13648 22545 13676 22918
rect 13450 22536 13506 22545
rect 13634 22536 13690 22545
rect 13506 22494 13584 22522
rect 13450 22471 13506 22480
rect 13452 22432 13504 22438
rect 13372 22380 13452 22386
rect 13372 22374 13504 22380
rect 13372 22358 13492 22374
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13372 21690 13400 22034
rect 13464 21894 13492 22358
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 13464 21146 13492 21830
rect 13556 21672 13584 22494
rect 13740 22506 13768 23038
rect 14094 23015 14150 23024
rect 13634 22471 13690 22480
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13740 21962 13768 22442
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 13820 21684 13872 21690
rect 13556 21644 13820 21672
rect 13820 21626 13872 21632
rect 14016 21350 14044 21966
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20262 13400 20946
rect 13924 20466 13952 21014
rect 14016 20913 14044 21286
rect 14002 20904 14058 20913
rect 14002 20839 14058 20848
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13372 20097 13400 20198
rect 13358 20088 13414 20097
rect 13924 20058 13952 20402
rect 13358 20023 13414 20032
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13372 19310 13400 19654
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13372 18970 13400 19246
rect 13832 19242 13860 19654
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13372 17678 13400 18906
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13740 18222 13768 18566
rect 13728 18216 13780 18222
rect 13634 18184 13690 18193
rect 13728 18158 13780 18164
rect 13634 18119 13690 18128
rect 13648 18086 13676 18119
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13740 17882 13768 18158
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13832 17814 13860 19178
rect 14108 18426 14136 23015
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 14200 19174 14228 20266
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14292 19174 14320 19858
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17354 13400 17614
rect 13372 17326 13492 17354
rect 13280 17224 13400 17252
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13188 17105 13216 17138
rect 13174 17096 13230 17105
rect 13174 17031 13230 17040
rect 12992 16992 13044 16998
rect 12990 16960 12992 16969
rect 13044 16960 13046 16969
rect 12990 16895 13046 16904
rect 12622 16824 12678 16833
rect 12622 16759 12678 16768
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12728 16454 12756 16730
rect 13188 16697 13216 17031
rect 13174 16688 13230 16697
rect 13174 16623 13230 16632
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12360 16102 12480 16130
rect 12360 16046 12388 16102
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12084 15558 12388 15586
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 13462 12112 14214
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 13530 12204 13874
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11716 12430 11836 12458
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11624 11898 11652 12310
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11716 11778 11744 12430
rect 11900 12102 11928 12582
rect 11992 12481 12020 12718
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 11978 12472 12034 12481
rect 11978 12407 11980 12416
rect 12032 12407 12034 12416
rect 11980 12378 12032 12384
rect 11992 12347 12020 12378
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11164 10798 11468 10826
rect 11624 11750 11744 11778
rect 10980 10662 11100 10690
rect 11072 10606 11100 10662
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10966 10432 11022 10441
rect 10612 10220 10732 10248
rect 10612 9450 10640 10220
rect 10888 9926 10916 10406
rect 10966 10367 11022 10376
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9722 10916 9862
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10046 3904 10102 3913
rect 10046 3839 10102 3848
rect 10152 3641 10180 9386
rect 10782 9344 10838 9353
rect 10289 9276 10585 9296
rect 10782 9279 10838 9288
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8634 10364 8910
rect 10796 8634 10824 9279
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10980 8480 11008 10367
rect 10796 8452 11008 8480
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10598 7440 10654 7449
rect 10598 7375 10654 7384
rect 10612 7342 10640 7375
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 6610 10824 8452
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 7750 10916 8230
rect 11164 8022 11192 10798
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11440 10266 11468 10610
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9382 11284 9998
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 8974 11284 9318
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11440 8838 11468 8978
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11440 8498 11468 8774
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11336 8424 11388 8430
rect 11334 8392 11336 8401
rect 11388 8392 11390 8401
rect 11334 8327 11390 8336
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7449 10916 7686
rect 10874 7440 10930 7449
rect 10874 7375 10930 7384
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11072 7002 11100 7210
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10796 6582 11008 6610
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10796 5710 10824 6122
rect 10784 5704 10836 5710
rect 10782 5672 10784 5681
rect 10836 5672 10838 5681
rect 10782 5607 10838 5616
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10138 3632 10194 3641
rect 10138 3567 10194 3576
rect 10782 3496 10838 3505
rect 10782 3431 10838 3440
rect 10796 3194 10824 3431
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10796 2990 10824 3130
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10888 2825 10916 3062
rect 10874 2816 10930 2825
rect 10289 2748 10585 2768
rect 10874 2751 10930 2760
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10874 2680 10930 2689
rect 10874 2615 10876 2624
rect 10928 2615 10930 2624
rect 10876 2586 10928 2592
rect 10980 2530 11008 6582
rect 11072 6390 11100 6938
rect 11164 6662 11192 7822
rect 11256 7546 11284 7890
rect 11334 7712 11390 7721
rect 11334 7647 11390 7656
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11058 5672 11114 5681
rect 11058 5607 11114 5616
rect 11072 3097 11100 5607
rect 11152 3936 11204 3942
rect 11150 3904 11152 3913
rect 11204 3904 11206 3913
rect 11150 3839 11206 3848
rect 11150 3632 11206 3641
rect 11150 3567 11152 3576
rect 11204 3567 11206 3576
rect 11152 3538 11204 3544
rect 11164 3194 11192 3538
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11058 3088 11114 3097
rect 11256 3074 11284 7278
rect 11348 6186 11376 7647
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11334 6080 11390 6089
rect 11334 6015 11390 6024
rect 11348 5234 11376 6015
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11440 5098 11468 6258
rect 11624 6254 11652 11750
rect 11900 11558 11928 12038
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11900 11218 11928 11494
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11716 6746 11744 11018
rect 11900 11014 11928 11154
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 9586 11836 10406
rect 11900 10198 11928 10950
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11716 6718 11836 6746
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11716 5778 11744 6598
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11610 4992 11666 5001
rect 11610 4927 11666 4936
rect 11336 4072 11388 4078
rect 11334 4040 11336 4049
rect 11388 4040 11390 4049
rect 11334 3975 11390 3984
rect 11518 4040 11574 4049
rect 11518 3975 11574 3984
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3233 11468 3878
rect 11532 3738 11560 3975
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11624 3618 11652 4927
rect 11532 3590 11652 3618
rect 11426 3224 11482 3233
rect 11426 3159 11482 3168
rect 11428 3120 11480 3126
rect 11058 3023 11114 3032
rect 11164 3046 11284 3074
rect 11426 3088 11428 3097
rect 11480 3088 11482 3097
rect 10520 2502 11008 2530
rect 10520 480 10548 2502
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 1737 10824 2246
rect 10782 1728 10838 1737
rect 10782 1663 10838 1672
rect 11164 480 11192 3046
rect 11426 3023 11482 3032
rect 11532 2514 11560 3590
rect 11716 3398 11744 5714
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11808 3194 11836 6718
rect 11900 6458 11928 6870
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 3482 12020 8230
rect 12084 7342 12112 12650
rect 12176 12374 12204 13466
rect 12254 13016 12310 13025
rect 12254 12951 12256 12960
rect 12308 12951 12310 12960
rect 12256 12922 12308 12928
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12360 11098 12388 15558
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 15162 12480 15302
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12728 15026 12756 16390
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15366 12848 15846
rect 13004 15706 13032 16050
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12438 12880 12494 12889
rect 12438 12815 12494 12824
rect 12452 12782 12480 12815
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12544 12345 12572 14758
rect 12728 14618 12756 14962
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13433 12940 13670
rect 12898 13424 12954 13433
rect 12898 13359 12900 13368
rect 12952 13359 12954 13368
rect 12900 13330 12952 13336
rect 13096 13297 13124 15574
rect 13174 15464 13230 15473
rect 13174 15399 13230 15408
rect 13188 14618 13216 15399
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13082 13288 13138 13297
rect 13082 13223 13138 13232
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12440 11688 12492 11694
rect 12438 11656 12440 11665
rect 12492 11656 12494 11665
rect 12438 11591 12494 11600
rect 12360 11070 12480 11098
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 10674 12388 10950
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 7002 12112 7142
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12176 5794 12204 10406
rect 12360 10130 12388 10610
rect 12452 10305 12480 11070
rect 12438 10296 12494 10305
rect 12438 10231 12494 10240
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12360 9382 12388 10066
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 9178 12388 9318
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12452 7970 12480 10231
rect 12544 9568 12572 12271
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12728 10266 12756 11154
rect 12898 10704 12954 10713
rect 12898 10639 12954 10648
rect 12912 10606 12940 10639
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12808 9580 12860 9586
rect 12544 9540 12756 9568
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12544 8634 12572 9386
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12452 7942 12572 7970
rect 12438 7848 12494 7857
rect 12438 7783 12494 7792
rect 12452 7546 12480 7783
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12268 6458 12296 6938
rect 12452 6746 12480 7278
rect 12360 6718 12480 6746
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12360 5914 12388 6718
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12438 5808 12494 5817
rect 12072 5772 12124 5778
rect 12176 5766 12388 5794
rect 12072 5714 12124 5720
rect 12084 5302 12112 5714
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12176 5370 12204 5646
rect 12360 5545 12388 5766
rect 12438 5743 12494 5752
rect 12346 5536 12402 5545
rect 12346 5471 12402 5480
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12084 4826 12112 5238
rect 12176 4826 12204 5306
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12452 4078 12480 5743
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12544 3602 12572 7942
rect 12636 6322 12664 8298
rect 12728 7188 12756 9540
rect 12808 9522 12860 9528
rect 12820 9178 12848 9522
rect 12900 9376 12952 9382
rect 12898 9344 12900 9353
rect 12952 9344 12954 9353
rect 12898 9279 12954 9288
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12898 8936 12954 8945
rect 12898 8871 12954 8880
rect 12912 8566 12940 8871
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12912 8362 12940 8502
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7342 12940 7686
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12728 7160 12940 7188
rect 12806 7032 12862 7041
rect 12806 6967 12862 6976
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 6390 12756 6734
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12728 5710 12756 6326
rect 12820 5914 12848 6967
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 4758 12756 5646
rect 12820 5234 12848 5850
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12820 4282 12848 4694
rect 12912 4622 12940 7160
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12912 4214 12940 4558
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3777 12664 3878
rect 12622 3768 12678 3777
rect 13004 3738 13032 12038
rect 13096 9722 13124 13223
rect 13174 12880 13230 12889
rect 13174 12815 13230 12824
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13188 9654 13216 12815
rect 13280 11665 13308 13806
rect 13372 11762 13400 17224
rect 13464 16794 13492 17326
rect 13832 17270 13860 17750
rect 13924 17649 13952 18362
rect 14200 18290 14228 19110
rect 14292 18630 14320 19110
rect 14280 18624 14332 18630
rect 14278 18592 14280 18601
rect 14332 18592 14334 18601
rect 14278 18527 14334 18536
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17882 14320 18022
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14094 17776 14150 17785
rect 14094 17711 14096 17720
rect 14148 17711 14150 17720
rect 14096 17682 14148 17688
rect 13910 17640 13966 17649
rect 13910 17575 13966 17584
rect 14096 17604 14148 17610
rect 14096 17546 14148 17552
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13648 16833 13676 16934
rect 13634 16824 13690 16833
rect 13452 16788 13504 16794
rect 13634 16759 13690 16768
rect 13452 16730 13504 16736
rect 13832 16114 13860 17206
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 16182 13952 16594
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13924 15706 13952 16118
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13450 15600 13506 15609
rect 13450 15535 13506 15544
rect 13820 15564 13872 15570
rect 13464 14074 13492 15535
rect 13820 15506 13872 15512
rect 13832 15162 13860 15506
rect 13820 15156 13872 15162
rect 13556 15116 13820 15144
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13266 11656 13322 11665
rect 13266 11591 13322 11600
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12622 3703 12678 3712
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12348 3528 12400 3534
rect 11992 3454 12112 3482
rect 12348 3470 12400 3476
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11808 2990 11836 3130
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 12084 2666 12112 3454
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 2990 12204 3334
rect 12360 3194 12388 3470
rect 12544 3194 12572 3538
rect 12348 3188 12400 3194
rect 12532 3188 12584 3194
rect 12400 3148 12480 3176
rect 12348 3130 12400 3136
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 11900 2638 12112 2666
rect 12452 2650 12480 3148
rect 12532 3130 12584 3136
rect 13004 2990 13032 3674
rect 12992 2984 13044 2990
rect 12530 2952 12586 2961
rect 12992 2926 13044 2932
rect 12530 2887 12586 2896
rect 12440 2644 12492 2650
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 2009 11652 2246
rect 11610 2000 11666 2009
rect 11610 1935 11666 1944
rect 11900 480 11928 2638
rect 12440 2586 12492 2592
rect 12544 2514 12572 2887
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 13096 2310 13124 8570
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12544 480 12572 2246
rect 13188 480 13216 9454
rect 13280 8634 13308 9522
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13266 8528 13322 8537
rect 13266 8463 13322 8472
rect 13280 8430 13308 8463
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13464 6769 13492 10406
rect 13450 6760 13506 6769
rect 13450 6695 13506 6704
rect 13268 6248 13320 6254
rect 13266 6216 13268 6225
rect 13320 6216 13322 6225
rect 13266 6151 13322 6160
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13266 5128 13322 5137
rect 13266 5063 13322 5072
rect 13280 5030 13308 5063
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13372 4622 13400 5170
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13372 4282 13400 4558
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13556 3738 13584 15116
rect 13820 15098 13872 15104
rect 13832 15033 13860 15098
rect 14016 15094 14044 16050
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13648 13530 13676 14350
rect 13740 14074 13768 14962
rect 14004 14952 14056 14958
rect 13818 14920 13874 14929
rect 14004 14894 14056 14900
rect 13818 14855 13874 14864
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13740 13841 13768 13874
rect 13726 13832 13782 13841
rect 13726 13767 13782 13776
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13832 12866 13860 14855
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14498 13952 14758
rect 14016 14618 14044 14894
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13924 14482 14044 14498
rect 13924 14476 14056 14482
rect 13924 14470 14004 14476
rect 14004 14418 14056 14424
rect 14016 14074 14044 14418
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14108 13954 14136 17546
rect 14292 17338 14320 17818
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14278 16144 14334 16153
rect 14278 16079 14334 16088
rect 14292 16046 14320 16079
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14186 15736 14242 15745
rect 14186 15671 14242 15680
rect 14200 15638 14228 15671
rect 14188 15632 14240 15638
rect 14188 15574 14240 15580
rect 14384 15026 14412 24686
rect 15304 24698 15332 27520
rect 15474 24848 15530 24857
rect 15474 24783 15530 24792
rect 15120 24682 15332 24698
rect 14922 24647 14978 24656
rect 15108 24676 15332 24682
rect 14936 24614 14964 24647
rect 15160 24670 15332 24676
rect 15108 24618 15160 24624
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14752 23866 14780 24210
rect 14832 24064 14884 24070
rect 14832 24006 14884 24012
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14844 23730 14872 24006
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 14554 23352 14610 23361
rect 14554 23287 14610 23296
rect 14462 19408 14518 19417
rect 14462 19343 14518 19352
rect 14476 16726 14504 19343
rect 14568 17202 14596 23287
rect 15212 23118 15240 23530
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 14752 22778 14780 23054
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 15290 22536 15346 22545
rect 15290 22471 15346 22480
rect 15304 22098 15332 22471
rect 15396 22234 15424 23122
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14660 21622 14688 21830
rect 14844 21690 14872 21830
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21690 15332 22034
rect 15396 21842 15424 22170
rect 15488 21962 15516 24783
rect 15948 24721 15976 27520
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 15934 24712 15990 24721
rect 15934 24647 15990 24656
rect 15842 24440 15898 24449
rect 15842 24375 15844 24384
rect 15896 24375 15898 24384
rect 15844 24346 15896 24352
rect 15658 23488 15714 23497
rect 15658 23423 15714 23432
rect 15568 22024 15620 22030
rect 15566 21992 15568 22001
rect 15620 21992 15622 22001
rect 15476 21956 15528 21962
rect 15566 21927 15622 21936
rect 15476 21898 15528 21904
rect 15396 21814 15608 21842
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14660 21185 14688 21286
rect 14646 21176 14702 21185
rect 14646 21111 14702 21120
rect 14660 20806 14688 21111
rect 15396 21078 15424 21490
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 13924 13926 14136 13954
rect 13924 13002 13952 13926
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14016 13161 14044 13330
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14002 13152 14058 13161
rect 14002 13087 14058 13096
rect 13924 12974 14044 13002
rect 14108 12986 14136 13262
rect 13832 12838 13952 12866
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13648 11393 13676 12650
rect 13740 12084 13768 12718
rect 13832 12442 13860 12718
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13820 12096 13872 12102
rect 13740 12056 13820 12084
rect 13820 12038 13872 12044
rect 13832 11694 13860 12038
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13634 11384 13690 11393
rect 13740 11354 13768 11562
rect 13634 11319 13690 11328
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13832 11218 13860 11630
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13832 9926 13860 11154
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13636 7744 13688 7750
rect 13924 7721 13952 12838
rect 14016 11014 14044 12974
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14200 10810 14228 14214
rect 14292 13802 14320 14350
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12782 14320 13262
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14004 10464 14056 10470
rect 14002 10432 14004 10441
rect 14056 10432 14058 10441
rect 14002 10367 14058 10376
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14108 9178 14136 10066
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14108 8906 14136 9114
rect 14200 8974 14228 9862
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14096 8424 14148 8430
rect 14200 8412 14228 8910
rect 14148 8384 14228 8412
rect 14096 8366 14148 8372
rect 14384 8276 14412 14826
rect 14568 13784 14596 17138
rect 14476 13756 14596 13784
rect 14476 12696 14504 13756
rect 14660 13705 14688 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15396 20602 15424 21014
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 14738 19952 14794 19961
rect 14738 19887 14794 19896
rect 14752 18086 14780 19887
rect 15580 19854 15608 21814
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15580 19174 15608 19790
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 14830 18864 14886 18873
rect 14830 18799 14832 18808
rect 14884 18799 14886 18808
rect 14832 18770 14884 18776
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14844 18154 14872 18362
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14936 17678 14964 18022
rect 14924 17672 14976 17678
rect 14738 17640 14794 17649
rect 14924 17614 14976 17620
rect 14738 17575 14794 17584
rect 14752 17202 14780 17575
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17338 15332 18702
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15396 17202 15424 18294
rect 15488 18290 15516 18566
rect 15580 18290 15608 19110
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15488 18068 15516 18226
rect 15568 18080 15620 18086
rect 15488 18040 15568 18068
rect 15568 18022 15620 18028
rect 15580 17746 15608 18022
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 14752 16794 14780 17138
rect 15382 17096 15438 17105
rect 15382 17031 15438 17040
rect 15290 16960 15346 16969
rect 15290 16895 15346 16904
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16130 15332 16895
rect 15396 16250 15424 17031
rect 15580 16998 15608 17682
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15304 16102 15424 16130
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14646 13696 14702 13705
rect 14646 13631 14702 13640
rect 14646 13560 14702 13569
rect 14646 13495 14702 13504
rect 14476 12668 14596 12696
rect 14462 12608 14518 12617
rect 14462 12543 14518 12552
rect 14476 11121 14504 12543
rect 14462 11112 14518 11121
rect 14462 11047 14518 11056
rect 14462 10976 14518 10985
rect 14462 10911 14518 10920
rect 14200 8248 14412 8276
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14004 7744 14056 7750
rect 13636 7686 13688 7692
rect 13910 7712 13966 7721
rect 13648 4826 13676 7686
rect 14004 7686 14056 7692
rect 13910 7647 13966 7656
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13740 6254 13768 7375
rect 14016 6934 14044 7686
rect 14108 7546 14136 7958
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 14016 6322 14044 6870
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 14016 6202 14044 6258
rect 13740 5914 13768 6190
rect 14016 6174 14136 6202
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5914 14044 6054
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14108 5794 14136 6174
rect 14016 5766 14136 5794
rect 13740 5642 13860 5658
rect 13740 5636 13872 5642
rect 13740 5630 13820 5636
rect 13740 5370 13768 5630
rect 13820 5578 13872 5584
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13648 4078 13676 4762
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13832 3641 13860 3946
rect 13924 3738 13952 5510
rect 14016 5370 14044 5766
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14108 4826 14136 5646
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14108 4282 14136 4762
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13818 3632 13874 3641
rect 13728 3596 13780 3602
rect 14200 3618 14228 8248
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14292 7002 14320 8026
rect 14372 7880 14424 7886
rect 14370 7848 14372 7857
rect 14424 7848 14426 7857
rect 14370 7783 14426 7792
rect 14384 7478 14412 7783
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14384 6934 14412 7142
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14476 4690 14504 10911
rect 14568 10674 14596 12668
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14660 10198 14688 13495
rect 14752 12918 14780 13738
rect 14844 13530 14872 14554
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13954 15332 14350
rect 15396 14226 15424 16102
rect 15488 15570 15516 16390
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15488 15473 15516 15506
rect 15474 15464 15530 15473
rect 15580 15434 15608 16594
rect 15672 15638 15700 23423
rect 15856 23322 15884 24346
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 16040 23866 16068 24142
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 16040 23322 16068 23802
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 15856 22273 15884 23258
rect 16040 22778 16068 23258
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15842 22264 15898 22273
rect 15842 22199 15898 22208
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15764 19417 15792 21898
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15948 21418 15976 21558
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 15948 20806 15976 21354
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16040 21146 16068 21286
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15948 20262 15976 20742
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19922 15976 20198
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 15842 19816 15898 19825
rect 15842 19751 15898 19760
rect 15750 19408 15806 19417
rect 15750 19343 15806 19352
rect 15856 18850 15884 19751
rect 15948 18970 15976 19858
rect 16040 19378 16068 20538
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15856 18822 15976 18850
rect 15750 16688 15806 16697
rect 15750 16623 15752 16632
rect 15804 16623 15806 16632
rect 15752 16594 15804 16600
rect 15844 16584 15896 16590
rect 15750 16552 15806 16561
rect 15844 16526 15896 16532
rect 15750 16487 15806 16496
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15474 15399 15530 15408
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 14346 15608 15370
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15396 14198 15608 14226
rect 15382 14104 15438 14113
rect 15382 14039 15438 14048
rect 15120 13926 15332 13954
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14936 13410 14964 13738
rect 15120 13530 15148 13926
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15212 13410 15240 13806
rect 15396 13802 15424 14039
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 14844 13382 14964 13410
rect 15120 13382 15240 13410
rect 15384 13388 15436 13394
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14844 12617 14872 13382
rect 15120 13326 15148 13382
rect 15384 13330 15436 13336
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12968 15332 13194
rect 15212 12940 15332 12968
rect 14830 12608 14886 12617
rect 14830 12543 14886 12552
rect 15212 12442 15240 12940
rect 15396 12442 15424 13330
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15108 12232 15160 12238
rect 15106 12200 15108 12209
rect 15160 12200 15162 12209
rect 15106 12135 15162 12144
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15488 11898 15516 13806
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14738 11248 14794 11257
rect 14738 11183 14794 11192
rect 14752 10266 14780 11183
rect 14844 10674 14872 11290
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14830 10568 14886 10577
rect 14830 10503 14886 10512
rect 14844 10470 14872 10503
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14568 7342 14596 8842
rect 14752 8430 14780 9522
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14740 8424 14792 8430
rect 15304 8378 15332 9318
rect 14740 8366 14792 8372
rect 15120 8350 15332 8378
rect 15120 8022 15148 8350
rect 15108 8016 15160 8022
rect 15396 7993 15424 11222
rect 15580 9058 15608 14198
rect 15488 9030 15608 9058
rect 15488 8838 15516 9030
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15474 8664 15530 8673
rect 15474 8599 15530 8608
rect 15108 7958 15160 7964
rect 15382 7984 15438 7993
rect 15382 7919 15438 7928
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15488 7410 15516 8599
rect 15580 7954 15608 8910
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14568 7002 14596 7278
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6322 15332 7142
rect 15488 7002 15516 7346
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15384 6860 15436 6866
rect 15436 6820 15516 6848
rect 15384 6802 15436 6808
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 14740 6112 14792 6118
rect 14738 6080 14740 6089
rect 14792 6080 14794 6089
rect 14738 6015 14794 6024
rect 15304 5914 15332 6258
rect 15488 6118 15516 6820
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14844 4826 14872 5102
rect 15396 4826 15424 6054
rect 15580 5642 15608 6258
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15580 5370 15608 5578
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14278 4584 14334 4593
rect 14278 4519 14280 4528
rect 14332 4519 14334 4528
rect 14280 4490 14332 4496
rect 14476 4214 14504 4626
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14844 4162 14872 4762
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14924 4208 14976 4214
rect 14844 4156 14924 4162
rect 15304 4162 15332 4626
rect 14844 4150 14976 4156
rect 13818 3567 13874 3576
rect 13924 3590 14228 3618
rect 14476 3602 14504 4150
rect 14844 4134 14964 4150
rect 15120 4134 15332 4162
rect 15120 3738 15148 4134
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15566 3904 15622 3913
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15212 3641 15240 3878
rect 15566 3839 15622 3848
rect 15580 3670 15608 3839
rect 15568 3664 15620 3670
rect 15198 3632 15254 3641
rect 14464 3596 14516 3602
rect 13728 3538 13780 3544
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 2961 13676 3334
rect 13634 2952 13690 2961
rect 13268 2916 13320 2922
rect 13634 2887 13690 2896
rect 13268 2858 13320 2864
rect 13280 2582 13308 2858
rect 13740 2650 13768 3538
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13280 2446 13308 2518
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13726 2408 13782 2417
rect 13726 2343 13728 2352
rect 13780 2343 13782 2352
rect 13728 2314 13780 2320
rect 13924 480 13952 3590
rect 15568 3606 15620 3612
rect 15198 3567 15254 3576
rect 14464 3538 14516 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 3194 14044 3470
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14554 3224 14610 3233
rect 14004 3188 14056 3194
rect 14956 3216 15252 3236
rect 14554 3159 14610 3168
rect 14004 3130 14056 3136
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 1873 14504 2246
rect 14462 1864 14518 1873
rect 14462 1799 14518 1808
rect 14568 480 14596 3159
rect 15396 2854 15424 3334
rect 15384 2848 15436 2854
rect 15290 2816 15346 2825
rect 15384 2790 15436 2796
rect 15290 2751 15346 2760
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 14844 2310 14872 2450
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 1601 14872 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14830 1592 14886 1601
rect 14830 1527 14886 1536
rect 15304 480 15332 2751
rect 15396 2650 15424 2790
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15672 2446 15700 15438
rect 15764 15065 15792 16487
rect 15856 15706 15884 16526
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15856 15337 15884 15642
rect 15842 15328 15898 15337
rect 15948 15314 15976 18822
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16040 18086 16068 18770
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16040 15502 16068 18022
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15948 15286 16068 15314
rect 15842 15263 15898 15272
rect 15750 15056 15806 15065
rect 15750 14991 15806 15000
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 13870 15792 14758
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15752 13864 15804 13870
rect 15750 13832 15752 13841
rect 15804 13832 15806 13841
rect 15750 13767 15806 13776
rect 15948 13258 15976 14418
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15948 12345 15976 12378
rect 15934 12336 15990 12345
rect 15844 12300 15896 12306
rect 15934 12271 15990 12280
rect 15844 12242 15896 12248
rect 15856 11558 15884 12242
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 10538 15884 11494
rect 15948 11354 15976 12174
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16040 11286 16068 15286
rect 16132 13462 16160 26386
rect 16396 25356 16448 25362
rect 16396 25298 16448 25304
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16316 24614 16344 24686
rect 16304 24608 16356 24614
rect 16304 24550 16356 24556
rect 16408 24562 16436 25298
rect 16592 24698 16620 27520
rect 16500 24682 16620 24698
rect 16488 24676 16620 24682
rect 16540 24670 16620 24676
rect 16488 24618 16540 24624
rect 16580 24608 16632 24614
rect 16408 24556 16580 24562
rect 16408 24550 16632 24556
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 16224 20369 16252 20538
rect 16210 20360 16266 20369
rect 16210 20295 16212 20304
rect 16264 20295 16266 20304
rect 16212 20266 16264 20272
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16224 17814 16252 18566
rect 16212 17808 16264 17814
rect 16212 17750 16264 17756
rect 16316 17354 16344 24550
rect 16408 24534 16620 24550
rect 16408 23361 16436 24534
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16394 23352 16450 23361
rect 16394 23287 16450 23296
rect 16500 22624 16528 24006
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 16684 23186 16712 23598
rect 16960 23526 16988 24210
rect 16948 23520 17000 23526
rect 16946 23488 16948 23497
rect 17000 23488 17002 23497
rect 16946 23423 17002 23432
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16580 22636 16632 22642
rect 16500 22596 16580 22624
rect 16580 22578 16632 22584
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16684 22030 16712 22374
rect 17052 22234 17080 22578
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 17038 22128 17094 22137
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16500 21554 16528 21830
rect 16684 21690 16712 21966
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16394 20224 16450 20233
rect 16394 20159 16450 20168
rect 16408 19514 16436 20159
rect 16592 20097 16620 21354
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16776 20330 16804 20742
rect 16868 20466 16896 21082
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16578 20088 16634 20097
rect 16776 20058 16804 20266
rect 16578 20023 16634 20032
rect 16764 20052 16816 20058
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16592 18766 16620 20023
rect 16764 19994 16816 20000
rect 16960 19394 16988 22102
rect 17038 22063 17094 22072
rect 17052 20369 17080 22063
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17144 21690 17172 21830
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17144 21486 17172 21626
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17236 20618 17264 24550
rect 17328 24410 17356 27520
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17604 23526 17632 24210
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17512 22642 17540 22918
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17420 21350 17448 22510
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17144 20590 17264 20618
rect 17038 20360 17094 20369
rect 17038 20295 17094 20304
rect 16868 19366 16988 19394
rect 16868 19310 16896 19366
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16396 18216 16448 18222
rect 16394 18184 16396 18193
rect 16448 18184 16450 18193
rect 16394 18119 16450 18128
rect 16316 17326 16436 17354
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16114 16252 16934
rect 16316 16794 16344 17138
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16316 15706 16344 15982
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16408 14929 16436 17326
rect 16500 17134 16528 18566
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16592 17882 16620 18158
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16684 17202 16712 17546
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16500 16794 16528 17070
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 15910 16712 16594
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16394 14920 16450 14929
rect 16394 14855 16450 14864
rect 16500 14822 16528 15302
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16592 14634 16620 15642
rect 16500 14618 16620 14634
rect 16488 14612 16620 14618
rect 16540 14606 16620 14612
rect 16488 14554 16540 14560
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 13938 16528 14214
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16684 13802 16712 15846
rect 16776 14822 16804 15846
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14414 16804 14758
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16868 14278 16896 15302
rect 16960 14521 16988 15914
rect 17052 14793 17080 20295
rect 17144 19174 17172 20590
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17236 20058 17264 20402
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17222 19952 17278 19961
rect 17222 19887 17278 19896
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 15706 17172 19110
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17144 15366 17172 15642
rect 17236 15570 17264 19887
rect 17314 18864 17370 18873
rect 17420 18834 17448 21286
rect 17314 18799 17370 18808
rect 17408 18828 17460 18834
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17236 15162 17264 15506
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17038 14784 17094 14793
rect 17038 14719 17094 14728
rect 16946 14512 17002 14521
rect 16946 14447 17002 14456
rect 17132 14408 17184 14414
rect 17130 14376 17132 14385
rect 17184 14376 17186 14385
rect 17130 14311 17186 14320
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16500 13569 16528 13670
rect 16486 13560 16542 13569
rect 16486 13495 16542 13504
rect 16120 13456 16172 13462
rect 16120 13398 16172 13404
rect 16132 12918 16160 13398
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 16118 12744 16174 12753
rect 16118 12679 16174 12688
rect 16132 12646 16160 12679
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16028 11280 16080 11286
rect 15934 11248 15990 11257
rect 16028 11222 16080 11228
rect 15934 11183 15990 11192
rect 15948 11150 15976 11183
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16040 10810 16068 11086
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 9450 15792 10406
rect 16040 10266 16068 10746
rect 16132 10674 16160 12582
rect 16224 12374 16252 12405
rect 16212 12368 16264 12374
rect 16210 12336 16212 12345
rect 16264 12336 16266 12345
rect 16210 12271 16266 12280
rect 16224 11898 16252 12271
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16132 10169 16160 10406
rect 16224 10266 16252 11834
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16118 10160 16174 10169
rect 16028 10124 16080 10130
rect 16118 10095 16174 10104
rect 16028 10066 16080 10072
rect 16040 10033 16068 10066
rect 16026 10024 16082 10033
rect 16026 9959 16082 9968
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15764 9178 15792 9386
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15764 8129 15792 8774
rect 15750 8120 15806 8129
rect 15750 8055 15806 8064
rect 15856 8022 15884 9862
rect 16040 9382 16068 9959
rect 16224 9722 16252 10202
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7410 15792 7686
rect 15856 7478 15884 7958
rect 15948 7857 15976 8502
rect 15934 7848 15990 7857
rect 15934 7783 15990 7792
rect 15844 7472 15896 7478
rect 15844 7414 15896 7420
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15764 7002 15792 7346
rect 15842 7168 15898 7177
rect 15842 7103 15898 7112
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5710 15792 6054
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15764 5030 15792 5646
rect 15856 5137 15884 7103
rect 15948 6866 15976 7783
rect 16040 7274 16068 9318
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16132 8634 16160 9046
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16224 8634 16252 8978
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16210 8120 16266 8129
rect 16120 8084 16172 8090
rect 16210 8055 16266 8064
rect 16120 8026 16172 8032
rect 16132 7546 16160 8026
rect 16224 7585 16252 8055
rect 16210 7576 16266 7585
rect 16120 7540 16172 7546
rect 16210 7511 16266 7520
rect 16120 7482 16172 7488
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6458 15976 6802
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15842 5128 15898 5137
rect 15842 5063 15898 5072
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15948 4282 15976 4558
rect 16118 4312 16174 4321
rect 15936 4276 15988 4282
rect 16118 4247 16174 4256
rect 15936 4218 15988 4224
rect 15934 4040 15990 4049
rect 15934 3975 15990 3984
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15948 480 15976 3975
rect 16132 3738 16160 4247
rect 16316 4146 16344 11494
rect 16408 10538 16436 13126
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16500 12442 16528 12650
rect 16776 12442 16804 12786
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16868 12322 16896 14214
rect 17236 14074 17264 15098
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 16684 12294 16896 12322
rect 16684 11540 16712 12294
rect 16762 12200 16818 12209
rect 16762 12135 16764 12144
rect 16816 12135 16818 12144
rect 16764 12106 16816 12112
rect 16776 11694 16804 12106
rect 16960 11914 16988 14010
rect 17328 13258 17356 18799
rect 17408 18770 17460 18776
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17420 18086 17448 18634
rect 17408 18080 17460 18086
rect 17406 18048 17408 18057
rect 17460 18048 17462 18057
rect 17406 17983 17462 17992
rect 17512 17202 17540 18702
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17512 16590 17540 17138
rect 17604 16726 17632 23462
rect 17880 23338 17908 24754
rect 17972 24410 18000 27520
rect 18708 25498 18736 27520
rect 18696 25492 18748 25498
rect 18696 25434 18748 25440
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 18236 23588 18288 23594
rect 18236 23530 18288 23536
rect 17880 23322 18000 23338
rect 17880 23316 18012 23322
rect 17880 23310 17960 23316
rect 17774 23216 17830 23225
rect 17774 23151 17830 23160
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17130 12200 17186 12209
rect 17130 12135 17186 12144
rect 16960 11886 17080 11914
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16856 11552 16908 11558
rect 16684 11512 16804 11540
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10690 16528 11154
rect 16580 10736 16632 10742
rect 16500 10684 16580 10690
rect 16500 10678 16632 10684
rect 16500 10662 16620 10678
rect 16672 10668 16724 10674
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16500 10282 16528 10662
rect 16672 10610 16724 10616
rect 16500 10266 16620 10282
rect 16500 10260 16632 10266
rect 16500 10254 16580 10260
rect 16580 10202 16632 10208
rect 16684 10062 16712 10610
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16592 9586 16620 9930
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16408 8820 16436 9522
rect 16684 9518 16712 9998
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 9110 16712 9454
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16488 8832 16540 8838
rect 16408 8792 16488 8820
rect 16408 7886 16436 8792
rect 16488 8774 16540 8780
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 8090 16528 8298
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16408 7546 16436 7822
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16394 5400 16450 5409
rect 16394 5335 16450 5344
rect 16408 4758 16436 5335
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16500 4622 16528 5782
rect 16776 5681 16804 11512
rect 16856 11494 16908 11500
rect 16868 11082 16896 11494
rect 16960 11354 16988 11698
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16868 9489 16896 10542
rect 16960 9926 16988 11086
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16854 9480 16910 9489
rect 16854 9415 16910 9424
rect 16762 5672 16818 5681
rect 16762 5607 16818 5616
rect 16868 5166 16896 9415
rect 17052 8294 17080 11886
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16776 4486 16804 4966
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16578 3768 16634 3777
rect 16120 3732 16172 3738
rect 16578 3703 16634 3712
rect 16120 3674 16172 3680
rect 16302 2816 16358 2825
rect 16302 2751 16358 2760
rect 16316 2650 16344 2751
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 16132 2310 16160 2450
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 1465 16160 2246
rect 16118 1456 16174 1465
rect 16118 1391 16174 1400
rect 16592 480 16620 3703
rect 16684 3505 16712 3946
rect 16776 3534 16804 4422
rect 16764 3528 16816 3534
rect 16670 3496 16726 3505
rect 16764 3470 16816 3476
rect 16670 3431 16726 3440
rect 16960 3194 16988 7142
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5681 17080 6054
rect 17038 5672 17094 5681
rect 17038 5607 17094 5616
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 17052 4729 17080 4966
rect 17038 4720 17094 4729
rect 17038 4655 17094 4664
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17052 2689 17080 4558
rect 17038 2680 17094 2689
rect 17038 2615 17094 2624
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16776 2281 16804 2382
rect 16762 2272 16818 2281
rect 16762 2207 16818 2216
rect 17144 921 17172 12135
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11529 17356 12038
rect 17314 11520 17370 11529
rect 17314 11455 17370 11464
rect 17328 11218 17356 11455
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17328 10810 17356 11154
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17314 10296 17370 10305
rect 17314 10231 17370 10240
rect 17328 9722 17356 10231
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17420 8945 17448 16186
rect 17512 16114 17540 16526
rect 17604 16250 17632 16662
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17696 15201 17724 18090
rect 17682 15192 17738 15201
rect 17682 15127 17738 15136
rect 17498 13424 17554 13433
rect 17498 13359 17554 13368
rect 17512 12238 17540 13359
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17498 12064 17554 12073
rect 17498 11999 17554 12008
rect 17512 10198 17540 11999
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17512 9382 17540 10134
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17406 8936 17462 8945
rect 17406 8871 17462 8880
rect 17512 8537 17540 9318
rect 17604 8634 17632 13194
rect 17788 12594 17816 23151
rect 17880 22794 17908 23310
rect 17960 23258 18012 23264
rect 18248 22982 18276 23530
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 17880 22778 18000 22794
rect 17880 22772 18012 22778
rect 17880 22766 17960 22772
rect 17960 22714 18012 22720
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 18156 21146 18184 21966
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18144 21004 18196 21010
rect 18144 20946 18196 20952
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17972 20618 18000 20878
rect 17880 20602 18000 20618
rect 17868 20596 18000 20602
rect 17920 20590 18000 20596
rect 17868 20538 17920 20544
rect 17972 19174 18000 20590
rect 18156 20233 18184 20946
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 18142 20224 18198 20233
rect 18142 20159 18198 20168
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17960 18896 18012 18902
rect 18064 18873 18092 19858
rect 18340 19417 18368 20266
rect 18432 19961 18460 24550
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18524 22438 18552 23054
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18512 22432 18564 22438
rect 18510 22400 18512 22409
rect 18564 22400 18566 22409
rect 18510 22335 18566 22344
rect 18510 22264 18566 22273
rect 18616 22234 18644 22918
rect 18510 22199 18566 22208
rect 18604 22228 18656 22234
rect 18524 20777 18552 22199
rect 18604 22170 18656 22176
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18510 20768 18566 20777
rect 18510 20703 18566 20712
rect 18616 19990 18644 21490
rect 18604 19984 18656 19990
rect 18418 19952 18474 19961
rect 18604 19926 18656 19932
rect 18418 19887 18474 19896
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18326 19408 18382 19417
rect 18326 19343 18382 19352
rect 18432 19310 18460 19654
rect 18616 19378 18644 19926
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18144 19304 18196 19310
rect 18420 19304 18472 19310
rect 18144 19246 18196 19252
rect 18418 19272 18420 19281
rect 18472 19272 18474 19281
rect 18156 19174 18184 19246
rect 18474 19230 18552 19258
rect 18418 19207 18474 19216
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17960 18838 18012 18844
rect 18050 18864 18106 18873
rect 17868 17876 17920 17882
rect 17972 17864 18000 18838
rect 18050 18799 18106 18808
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17920 17836 18000 17864
rect 17868 17818 17920 17824
rect 17880 17338 17908 17818
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 18064 17082 18092 18566
rect 17972 17054 18092 17082
rect 18156 17066 18184 19110
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18144 17060 18196 17066
rect 17972 16776 18000 17054
rect 18144 17002 18196 17008
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17880 16748 18000 16776
rect 17880 16046 17908 16748
rect 18064 16726 18092 16934
rect 18432 16794 18460 18770
rect 18524 17134 18552 19230
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18616 18154 18644 18702
rect 18604 18148 18656 18154
rect 18604 18090 18656 18096
rect 18602 18048 18658 18057
rect 18602 17983 18658 17992
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18052 16720 18104 16726
rect 17958 16688 18014 16697
rect 18052 16662 18104 16668
rect 18156 16658 18184 16730
rect 17958 16623 18014 16632
rect 18144 16652 18196 16658
rect 17972 16250 18000 16623
rect 18144 16594 18196 16600
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 18156 15706 18184 16594
rect 18524 16590 18552 17070
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18432 15910 18460 16458
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 15910 18552 16390
rect 18420 15904 18472 15910
rect 18512 15904 18564 15910
rect 18420 15846 18472 15852
rect 18510 15872 18512 15881
rect 18564 15872 18566 15881
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18432 15609 18460 15846
rect 18510 15807 18566 15816
rect 18418 15600 18474 15609
rect 18418 15535 18474 15544
rect 18510 15328 18566 15337
rect 18510 15263 18566 15272
rect 18326 15056 18382 15065
rect 18326 14991 18382 15000
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17972 13190 18000 14418
rect 18248 13462 18276 14758
rect 18340 13841 18368 14991
rect 18524 14618 18552 15263
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18524 14074 18552 14554
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18420 13864 18472 13870
rect 18326 13832 18382 13841
rect 18420 13806 18472 13812
rect 18326 13767 18382 13776
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17866 12880 17922 12889
rect 17866 12815 17922 12824
rect 17880 12782 17908 12815
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 18340 12714 18368 13767
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 17788 12566 18092 12594
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11898 17724 12174
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17682 11656 17738 11665
rect 17682 11591 17738 11600
rect 17696 10810 17724 11591
rect 17788 11558 17816 12310
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17682 10296 17738 10305
rect 17682 10231 17684 10240
rect 17736 10231 17738 10240
rect 17684 10202 17736 10208
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17696 8974 17724 9862
rect 17788 9586 17816 11494
rect 17972 11121 18000 11630
rect 17958 11112 18014 11121
rect 17958 11047 18014 11056
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17880 9625 17908 9998
rect 17866 9616 17922 9625
rect 17776 9580 17828 9586
rect 17866 9551 17922 9560
rect 17776 9522 17828 9528
rect 17880 9518 17908 9551
rect 17972 9518 18000 11047
rect 18064 10606 18092 12566
rect 18432 12442 18460 13806
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18524 13326 18552 13670
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18432 11898 18460 12378
rect 18524 12374 18552 12582
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18248 10266 18276 11290
rect 18524 11082 18552 12174
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18616 10713 18644 17983
rect 18708 17354 18736 24686
rect 18892 24614 18920 25298
rect 19352 24698 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19260 24682 19380 24698
rect 19248 24676 19380 24682
rect 19300 24670 19380 24676
rect 19248 24618 19300 24624
rect 18880 24608 18932 24614
rect 18880 24550 18932 24556
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20088 24410 20116 27520
rect 20260 25356 20312 25362
rect 20260 25298 20312 25304
rect 20272 24614 20300 25298
rect 20732 24698 20760 27520
rect 20640 24682 20760 24698
rect 20628 24676 20760 24682
rect 20680 24670 20760 24676
rect 20628 24618 20680 24624
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20720 24608 20772 24614
rect 21088 24608 21140 24614
rect 20720 24550 20772 24556
rect 21086 24576 21088 24585
rect 21140 24576 21142 24585
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 18878 24168 18934 24177
rect 18878 24103 18934 24112
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18800 22982 18828 23598
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 22642 18828 22918
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 20398 18828 20742
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18788 20256 18840 20262
rect 18786 20224 18788 20233
rect 18840 20224 18842 20233
rect 18786 20159 18842 20168
rect 18892 18873 18920 24103
rect 20180 23526 20208 24210
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 19260 22506 19288 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19248 22500 19300 22506
rect 19248 22442 19300 22448
rect 19260 22234 19288 22442
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19248 22228 19300 22234
rect 19248 22170 19300 22176
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19444 21690 19472 21898
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19982 21584 20038 21593
rect 19982 21519 20038 21528
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21010 19564 21286
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19996 21146 20024 21519
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 19156 20800 19208 20806
rect 19156 20742 19208 20748
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19168 19922 19196 20742
rect 19352 20398 19380 20742
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19536 20058 19564 20946
rect 20088 20330 20116 22374
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 20052 19576 20058
rect 19444 20012 19524 20040
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19260 19174 19288 19246
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 18878 18864 18934 18873
rect 18878 18799 18934 18808
rect 18708 17326 18828 17354
rect 18694 17232 18750 17241
rect 18694 17167 18696 17176
rect 18748 17167 18750 17176
rect 18696 17138 18748 17144
rect 18800 16017 18828 17326
rect 18786 16008 18842 16017
rect 18786 15943 18842 15952
rect 18800 15706 18828 15943
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 15026 18736 15302
rect 18800 15162 18828 15642
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18786 15056 18842 15065
rect 18696 15020 18748 15026
rect 18786 14991 18842 15000
rect 18696 14962 18748 14968
rect 18708 14074 18736 14962
rect 18800 14890 18828 14991
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18892 14770 18920 18799
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19168 17882 19196 18090
rect 19352 18057 19380 19110
rect 19338 18048 19394 18057
rect 19338 17983 19394 17992
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 19444 17746 19472 20012
rect 19524 19994 19576 20000
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19536 18970 19564 19790
rect 19628 19514 19656 19858
rect 19996 19854 20024 20198
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19996 18902 20024 19790
rect 20088 19378 20116 20266
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20088 18902 20116 19314
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 20076 18896 20128 18902
rect 20076 18838 20128 18844
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19076 16998 19104 17682
rect 19444 17338 19472 17682
rect 19996 17649 20024 18022
rect 19982 17640 20038 17649
rect 19982 17575 20038 17584
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19536 17134 19564 17478
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 19260 16946 19288 17002
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18984 15706 19012 16662
rect 19076 16590 19104 16934
rect 19260 16918 19380 16946
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 19076 16250 19104 16526
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19260 15609 19288 15642
rect 19246 15600 19302 15609
rect 19246 15535 19302 15544
rect 18970 15328 19026 15337
rect 18970 15263 19026 15272
rect 18800 14742 18920 14770
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 18708 12782 18736 12951
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18800 12730 18828 14742
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18892 12889 18920 13262
rect 18878 12880 18934 12889
rect 18878 12815 18880 12824
rect 18932 12815 18934 12824
rect 18880 12786 18932 12792
rect 18800 12702 18920 12730
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11626 18736 12038
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18602 10704 18658 10713
rect 18708 10674 18736 11562
rect 18602 10639 18658 10648
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17880 9178 17908 9454
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17972 9081 18000 9454
rect 18248 9450 18276 10202
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 18328 9036 18380 9042
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17972 8838 18000 9007
rect 18328 8978 18380 8984
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8832 18012 8838
rect 17866 8800 17922 8809
rect 17960 8774 18012 8780
rect 17866 8735 17922 8744
rect 17880 8634 17908 8735
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17498 8528 17554 8537
rect 17972 8514 18000 8774
rect 17498 8463 17554 8472
rect 17880 8486 18000 8514
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7002 17448 8230
rect 17880 8090 17908 8486
rect 18064 8090 18092 8910
rect 18340 8634 18368 8978
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18064 7954 18092 8026
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18616 7857 18644 7890
rect 18602 7848 18658 7857
rect 18328 7812 18380 7818
rect 18602 7783 18658 7792
rect 18328 7754 18380 7760
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17512 6458 17540 7142
rect 17880 7041 17908 7482
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17972 7177 18000 7278
rect 17958 7168 18014 7177
rect 17958 7103 18014 7112
rect 17866 7032 17922 7041
rect 17866 6967 17922 6976
rect 18142 6896 18198 6905
rect 18340 6866 18368 7754
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18064 6840 18142 6848
rect 18064 6820 18144 6840
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 17880 4146 17908 6122
rect 18064 5914 18092 6820
rect 18196 6831 18198 6840
rect 18328 6860 18380 6866
rect 18144 6802 18196 6808
rect 18328 6802 18380 6808
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18248 6186 18276 6734
rect 18340 6458 18368 6802
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18156 4078 18184 6054
rect 18248 5778 18276 6122
rect 18340 5914 18368 6394
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18340 5234 18368 5850
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4622 18276 4966
rect 18432 4758 18460 5782
rect 18524 4758 18552 7686
rect 18616 7546 18644 7783
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18708 7313 18736 10474
rect 18800 10146 18828 12582
rect 18892 12306 18920 12702
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11257 18920 12038
rect 18878 11248 18934 11257
rect 18878 11183 18934 11192
rect 18984 10266 19012 15263
rect 19352 13870 19380 16918
rect 19430 15736 19486 15745
rect 19430 15671 19486 15680
rect 19444 14482 19472 15671
rect 19536 14958 19564 17070
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20088 16114 20116 16934
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20074 16008 20130 16017
rect 20074 15943 20130 15952
rect 20088 15910 20116 15943
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19524 14952 19576 14958
rect 19628 14929 19656 15506
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19524 14894 19576 14900
rect 19614 14920 19670 14929
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19536 14385 19564 14894
rect 19720 14890 19748 15438
rect 19904 14958 19932 15438
rect 19892 14952 19944 14958
rect 19944 14912 20024 14940
rect 19892 14894 19944 14900
rect 19614 14855 19616 14864
rect 19668 14855 19670 14864
rect 19708 14884 19760 14890
rect 19616 14826 19668 14832
rect 19708 14826 19760 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14550 20024 14912
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19522 14376 19578 14385
rect 19522 14311 19578 14320
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19076 12442 19104 12718
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11354 19104 12174
rect 19168 12102 19196 13330
rect 19260 13274 19288 13398
rect 19536 13326 19564 13466
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19524 13320 19576 13326
rect 19260 13246 19380 13274
rect 19628 13297 19656 13330
rect 19892 13320 19944 13326
rect 19524 13262 19576 13268
rect 19614 13288 19670 13297
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19260 11098 19288 13126
rect 19352 12442 19380 13246
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19340 11552 19392 11558
rect 19338 11520 19340 11529
rect 19392 11520 19394 11529
rect 19338 11455 19394 11464
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19352 11098 19380 11154
rect 19260 11070 19380 11098
rect 19154 10976 19210 10985
rect 19154 10911 19210 10920
rect 19168 10810 19196 10911
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18800 10118 19104 10146
rect 19260 10130 19288 11070
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10554 19380 10950
rect 19444 10674 19472 12310
rect 19536 10810 19564 13262
rect 19892 13262 19944 13268
rect 19614 13223 19670 13232
rect 19628 12986 19656 13223
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19904 12714 19932 13262
rect 19996 12986 20024 14010
rect 20074 13560 20130 13569
rect 20074 13495 20130 13504
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19996 12714 20024 12922
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19706 11112 19762 11121
rect 19706 11047 19762 11056
rect 19720 10810 19748 11047
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19904 10606 19932 10950
rect 20088 10690 20116 13495
rect 20180 11286 20208 23462
rect 20272 20890 20300 24550
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 22166 20576 22918
rect 20626 22264 20682 22273
rect 20626 22199 20682 22208
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 20548 21486 20576 22102
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20350 21040 20406 21049
rect 20350 20975 20352 20984
rect 20404 20975 20406 20984
rect 20352 20946 20404 20952
rect 20272 20862 20392 20890
rect 20258 20768 20314 20777
rect 20258 20703 20314 20712
rect 20272 18170 20300 20703
rect 20364 18426 20392 20862
rect 20456 20262 20484 21286
rect 20548 20398 20576 21422
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20548 20058 20576 20334
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 18850 20668 22199
rect 20732 19174 20760 24550
rect 21086 24511 21142 24520
rect 20810 24304 20866 24313
rect 20810 24239 20866 24248
rect 20996 24268 21048 24274
rect 20824 22681 20852 24239
rect 20996 24210 21048 24216
rect 21008 23594 21036 24210
rect 20996 23588 21048 23594
rect 20996 23530 21048 23536
rect 21178 23352 21234 23361
rect 21376 23322 21404 27520
rect 21640 26716 21692 26722
rect 21640 26658 21692 26664
rect 21546 24440 21602 24449
rect 21546 24375 21602 24384
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 21178 23287 21234 23296
rect 21364 23316 21416 23322
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20810 22672 20866 22681
rect 20810 22607 20866 22616
rect 21008 22438 21036 23122
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 20904 22092 20956 22098
rect 20904 22034 20956 22040
rect 20916 21010 20944 22034
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20902 20904 20958 20913
rect 20902 20839 20958 20848
rect 20810 20360 20866 20369
rect 20810 20295 20812 20304
rect 20864 20295 20866 20304
rect 20812 20266 20864 20272
rect 20916 20210 20944 20839
rect 21008 20505 21036 22374
rect 21088 20800 21140 20806
rect 21086 20768 21088 20777
rect 21140 20768 21142 20777
rect 21086 20703 21142 20712
rect 20994 20496 21050 20505
rect 20994 20431 21050 20440
rect 20824 20182 20944 20210
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20456 18822 20668 18850
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20350 18320 20406 18329
rect 20350 18255 20352 18264
rect 20404 18255 20406 18264
rect 20352 18226 20404 18232
rect 20272 18142 20392 18170
rect 20260 17060 20312 17066
rect 20260 17002 20312 17008
rect 20272 16794 20300 17002
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20272 13530 20300 14350
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 20272 11354 20300 12650
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20088 10662 20300 10690
rect 19892 10600 19944 10606
rect 19352 10526 19564 10554
rect 19892 10542 19944 10548
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18694 7304 18750 7313
rect 18694 7239 18750 7248
rect 18696 7200 18748 7206
rect 18800 7188 18828 8026
rect 18748 7160 18828 7188
rect 18880 7200 18932 7206
rect 18696 7142 18748 7148
rect 18880 7142 18932 7148
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18616 4826 18644 6054
rect 18708 5409 18736 7142
rect 18892 6934 18920 7142
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18892 6254 18920 6870
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18694 5400 18750 5409
rect 18694 5335 18750 5344
rect 18786 5128 18842 5137
rect 18786 5063 18788 5072
rect 18840 5063 18842 5072
rect 18788 5034 18840 5040
rect 18696 5024 18748 5030
rect 18694 4992 18696 5001
rect 18748 4992 18750 5001
rect 18694 4927 18750 4936
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18248 4282 18276 4558
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18524 3738 18552 4694
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18984 4282 19012 4558
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17328 2854 17356 3538
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18050 3224 18106 3233
rect 18050 3159 18052 3168
rect 18104 3159 18106 3168
rect 18052 3130 18104 3136
rect 17958 3088 18014 3097
rect 18156 3058 18184 3334
rect 17958 3023 18014 3032
rect 18144 3052 18196 3058
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17328 2650 17356 2790
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17328 2446 17356 2586
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17314 1728 17370 1737
rect 17314 1663 17370 1672
rect 17130 912 17186 921
rect 17130 847 17186 856
rect 17328 480 17356 1663
rect 17972 480 18000 3023
rect 18144 2994 18196 3000
rect 18156 2650 18184 2994
rect 18524 2854 18552 3334
rect 18880 2984 18932 2990
rect 18694 2952 18750 2961
rect 18880 2926 18932 2932
rect 18694 2887 18750 2896
rect 18512 2848 18564 2854
rect 18510 2816 18512 2825
rect 18564 2816 18566 2825
rect 18510 2751 18566 2760
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18156 2446 18184 2586
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18708 480 18736 2887
rect 18892 2582 18920 2926
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 19076 2417 19104 10118
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19352 9178 19380 10406
rect 19432 9648 19484 9654
rect 19430 9616 19432 9625
rect 19484 9616 19486 9625
rect 19430 9551 19486 9560
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19260 7342 19288 7958
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19352 6662 19380 7278
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6118 19380 6598
rect 19340 6112 19392 6118
rect 19260 6072 19340 6100
rect 19260 4622 19288 6072
rect 19340 6054 19392 6060
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19338 4584 19394 4593
rect 19338 4519 19394 4528
rect 19246 4040 19302 4049
rect 19246 3975 19302 3984
rect 19260 3738 19288 3975
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19062 2408 19118 2417
rect 19062 2343 19118 2352
rect 19076 1465 19104 2343
rect 19062 1456 19118 1465
rect 19062 1391 19118 1400
rect 19352 480 19380 4519
rect 19444 3738 19472 7822
rect 19536 5545 19564 10526
rect 20074 10432 20130 10441
rect 19622 10364 19918 10384
rect 20074 10367 20130 10376
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9194 20024 10066
rect 20088 10062 20116 10367
rect 20166 10296 20222 10305
rect 20166 10231 20168 10240
rect 20220 10231 20222 10240
rect 20168 10202 20220 10208
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20180 9722 20208 10202
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20074 9208 20130 9217
rect 19996 9166 20074 9194
rect 20074 9143 20076 9152
rect 20128 9143 20130 9152
rect 20168 9172 20220 9178
rect 20076 9114 20128 9120
rect 20168 9114 20220 9120
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19982 8528 20038 8537
rect 19982 8463 20038 8472
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19996 6633 20024 8463
rect 20088 7206 20116 8910
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20180 6905 20208 9114
rect 20272 8974 20300 10662
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20272 8362 20300 8774
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20364 7478 20392 18142
rect 20456 14618 20484 18822
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20548 16833 20576 18362
rect 20640 16969 20668 18702
rect 20626 16960 20682 16969
rect 20626 16895 20682 16904
rect 20534 16824 20590 16833
rect 20590 16782 20668 16810
rect 20534 16759 20590 16768
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20548 16182 20576 16390
rect 20536 16176 20588 16182
rect 20536 16118 20588 16124
rect 20548 16046 20576 16118
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20456 11676 20484 13806
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20548 12866 20576 13194
rect 20640 13025 20668 16782
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 15502 20760 16390
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20732 14618 20760 15438
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20824 14113 20852 20182
rect 20902 19680 20958 19689
rect 20902 19615 20958 19624
rect 20916 16028 20944 19615
rect 21008 19553 21036 20431
rect 21192 19990 21220 23287
rect 21364 23258 21416 23264
rect 21468 23202 21496 23598
rect 21376 23174 21496 23202
rect 21272 22568 21324 22574
rect 21270 22536 21272 22545
rect 21324 22536 21326 22545
rect 21270 22471 21326 22480
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21284 21146 21312 22034
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 20994 19544 21050 19553
rect 20994 19479 21050 19488
rect 21086 19408 21142 19417
rect 21086 19343 21142 19352
rect 21100 18850 21128 19343
rect 21180 19304 21232 19310
rect 21376 19281 21404 23174
rect 21560 22778 21588 24375
rect 21652 23866 21680 26658
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21454 22536 21510 22545
rect 21454 22471 21510 22480
rect 21468 21962 21496 22471
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21652 20913 21680 23530
rect 21638 20904 21694 20913
rect 21638 20839 21694 20848
rect 21180 19246 21232 19252
rect 21362 19272 21418 19281
rect 21192 18873 21220 19246
rect 21362 19207 21418 19216
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18970 21312 19110
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21008 18834 21128 18850
rect 21178 18864 21234 18873
rect 21008 18828 21140 18834
rect 21008 18822 21088 18828
rect 21008 18358 21036 18822
rect 21376 18834 21404 19207
rect 21178 18799 21234 18808
rect 21364 18828 21416 18834
rect 21088 18770 21140 18776
rect 21364 18770 21416 18776
rect 21086 18728 21142 18737
rect 21086 18663 21142 18672
rect 21100 18426 21128 18663
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 21284 18057 21312 18566
rect 21270 18048 21326 18057
rect 21744 18034 21772 24686
rect 21836 24682 21864 25298
rect 21824 24676 21876 24682
rect 21824 24618 21876 24624
rect 22112 24426 22140 27520
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22020 24410 22140 24426
rect 22008 24404 22140 24410
rect 22060 24398 22140 24404
rect 22008 24346 22060 24352
rect 22204 24070 22232 24686
rect 22756 24682 22784 27520
rect 23386 26616 23442 26625
rect 23386 26551 23442 26560
rect 23294 26072 23350 26081
rect 23294 26007 23350 26016
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22744 24676 22796 24682
rect 22744 24618 22796 24624
rect 22848 24614 22876 25298
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22282 24304 22338 24313
rect 22282 24239 22338 24248
rect 22376 24268 22428 24274
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22020 21486 22048 21830
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 21822 21176 21878 21185
rect 21822 21111 21824 21120
rect 21876 21111 21878 21120
rect 21824 21082 21876 21088
rect 22020 21010 22048 21422
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22020 20806 22048 20946
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22020 20058 22048 20198
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 22020 19530 22048 19994
rect 22112 19990 22140 20198
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22112 19666 22140 19926
rect 22204 19802 22232 24006
rect 22296 22273 22324 24239
rect 22376 24210 22428 24216
rect 22388 23730 22416 24210
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22742 22400 22798 22409
rect 22282 22264 22338 22273
rect 22282 22199 22338 22208
rect 22664 22137 22692 22374
rect 22742 22335 22798 22344
rect 22756 22234 22784 22335
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 22650 22128 22706 22137
rect 22650 22063 22706 22072
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22480 21350 22508 21966
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22664 21570 22692 21830
rect 22756 21690 22784 22170
rect 22848 22030 22876 24550
rect 23308 23866 23336 26007
rect 23400 24410 23428 26551
rect 23492 24449 23520 27520
rect 23662 25392 23718 25401
rect 23662 25327 23718 25336
rect 24032 25356 24084 25362
rect 23478 24440 23534 24449
rect 23388 24404 23440 24410
rect 23676 24410 23704 25327
rect 24032 25298 24084 25304
rect 24044 24614 24072 25298
rect 24136 25226 24164 27520
rect 24596 26450 24624 27639
rect 24766 27520 24822 28000
rect 25502 27520 25558 28000
rect 26146 27520 26202 28000
rect 26882 27520 26938 28000
rect 27526 27520 27582 28000
rect 24780 27282 24808 27520
rect 24688 27254 24808 27282
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 24688 25498 24716 27254
rect 24766 27160 24822 27169
rect 24766 27095 24822 27104
rect 24780 26722 24808 27095
rect 24768 26716 24820 26722
rect 24768 26658 24820 26664
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24780 24857 24808 25094
rect 24582 24848 24638 24857
rect 24582 24783 24638 24792
rect 24766 24848 24822 24857
rect 24766 24783 24822 24792
rect 24596 24750 24624 24783
rect 24584 24744 24636 24750
rect 24584 24686 24636 24692
rect 24032 24608 24084 24614
rect 24032 24550 24084 24556
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 23478 24375 23534 24384
rect 23664 24404 23716 24410
rect 23388 24346 23440 24352
rect 23664 24346 23716 24352
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 23492 23866 23520 24210
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23400 23576 23428 23666
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23400 23548 23520 23576
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23124 23254 23152 23462
rect 23492 23254 23520 23548
rect 23112 23248 23164 23254
rect 23112 23190 23164 23196
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23308 22778 23336 23122
rect 23584 22982 23612 23598
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 23032 21690 23060 21966
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 22664 21542 22784 21570
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22296 21078 22324 21286
rect 22284 21072 22336 21078
rect 22284 21014 22336 21020
rect 22204 19774 22324 19802
rect 22112 19638 22232 19666
rect 22020 19502 22140 19530
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21836 18902 21864 19314
rect 22006 19272 22062 19281
rect 21916 19236 21968 19242
rect 22006 19207 22062 19216
rect 21916 19178 21968 19184
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21270 17983 21326 17992
rect 21376 18006 21772 18034
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21192 16998 21220 17682
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21376 16776 21404 18006
rect 21546 17912 21602 17921
rect 21546 17847 21602 17856
rect 21100 16748 21404 16776
rect 20916 16000 21036 16028
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20916 15706 20944 15846
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20916 14618 20944 15506
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20810 14104 20866 14113
rect 20810 14039 20866 14048
rect 20824 13938 20852 14039
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20916 13870 20944 14350
rect 20904 13864 20956 13870
rect 20902 13832 20904 13841
rect 20956 13832 20958 13841
rect 20902 13767 20958 13776
rect 20626 13016 20682 13025
rect 20626 12951 20682 12960
rect 20548 12838 20668 12866
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 11830 20576 12582
rect 20640 12442 20668 12838
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20916 12306 20944 12718
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20732 11762 20760 12242
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20456 11648 20576 11676
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 9178 20484 10406
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 7546 20484 8230
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20166 6896 20222 6905
rect 20166 6831 20222 6840
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 19982 6624 20038 6633
rect 19982 6559 20038 6568
rect 20272 6254 20300 6734
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20272 5914 20300 6190
rect 20260 5908 20312 5914
rect 20180 5868 20260 5896
rect 20074 5672 20130 5681
rect 20074 5607 20130 5616
rect 19522 5536 19578 5545
rect 19522 5471 19578 5480
rect 19614 5264 19670 5273
rect 19614 5199 19616 5208
rect 19668 5199 19670 5208
rect 19616 5170 19668 5176
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19536 3942 19564 4422
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19444 3194 19472 3674
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19536 2650 19564 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19996 3738 20024 4966
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20088 480 20116 5607
rect 20180 4758 20208 5868
rect 20260 5850 20312 5856
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20272 4865 20300 4966
rect 20258 4856 20314 4865
rect 20258 4791 20260 4800
rect 20312 4791 20314 4800
rect 20260 4762 20312 4768
rect 20168 4752 20220 4758
rect 20272 4731 20300 4762
rect 20168 4694 20220 4700
rect 20180 4078 20208 4694
rect 20364 4486 20392 5170
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20180 3670 20208 4014
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 20180 2990 20208 3606
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20548 2446 20576 11648
rect 20916 11354 20944 12038
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 21008 10577 21036 16000
rect 21100 13326 21128 16748
rect 21270 16688 21326 16697
rect 21270 16623 21272 16632
rect 21324 16623 21326 16632
rect 21272 16594 21324 16600
rect 21284 15910 21312 16594
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21272 15904 21324 15910
rect 21192 15864 21272 15892
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21100 13161 21128 13262
rect 21086 13152 21142 13161
rect 21086 13087 21142 13096
rect 21100 12986 21128 13087
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21086 12880 21142 12889
rect 21086 12815 21142 12824
rect 21100 12646 21128 12815
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21100 12374 21128 12582
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21100 11898 21128 12310
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21192 11778 21220 15864
rect 21272 15846 21324 15852
rect 21468 15638 21496 16526
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21468 15434 21496 15574
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21362 15056 21418 15065
rect 21362 14991 21418 15000
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21284 14074 21312 14418
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21284 13870 21312 14010
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21100 11750 21220 11778
rect 20994 10568 21050 10577
rect 20994 10503 21050 10512
rect 21100 10266 21128 11750
rect 21284 10588 21312 13670
rect 21376 12594 21404 14991
rect 21468 14414 21496 15370
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21468 13462 21496 14350
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21356 12566 21404 12594
rect 21356 12424 21384 12566
rect 21356 12396 21404 12424
rect 21376 11540 21404 12396
rect 21560 11914 21588 17847
rect 21824 16788 21876 16794
rect 21928 16776 21956 19178
rect 22020 18426 22048 19207
rect 22112 18970 22140 19502
rect 22204 19446 22232 19638
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22112 17814 22140 18702
rect 22100 17808 22152 17814
rect 22100 17750 22152 17756
rect 22296 17626 22324 19774
rect 22480 19689 22508 21286
rect 22756 19922 22784 21542
rect 23032 21418 23060 21626
rect 23020 21412 23072 21418
rect 23020 21354 23072 21360
rect 23032 20602 23060 21354
rect 23020 20596 23072 20602
rect 23020 20538 23072 20544
rect 22928 20324 22980 20330
rect 22928 20266 22980 20272
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 22466 19680 22522 19689
rect 22466 19615 22522 19624
rect 22756 19417 22784 19858
rect 22940 19854 22968 20266
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22940 19514 22968 19790
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 22742 19408 22798 19417
rect 22742 19343 22798 19352
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22480 18222 22508 19110
rect 23124 18902 23152 19246
rect 23216 19009 23244 22374
rect 23308 20890 23336 22714
rect 23478 22672 23534 22681
rect 23478 22607 23534 22616
rect 23308 20862 23428 20890
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23308 20330 23336 20742
rect 23296 20324 23348 20330
rect 23296 20266 23348 20272
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23202 19000 23258 19009
rect 23202 18935 23258 18944
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23124 18426 23152 18838
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23308 18306 23336 19994
rect 23216 18278 23336 18306
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 23216 18154 23244 18278
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23204 18148 23256 18154
rect 23204 18090 23256 18096
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 22560 17808 22612 17814
rect 22466 17776 22522 17785
rect 22560 17750 22612 17756
rect 22466 17711 22522 17720
rect 22204 17598 22324 17626
rect 22100 16788 22152 16794
rect 21928 16748 22100 16776
rect 21824 16730 21876 16736
rect 22100 16730 22152 16736
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21652 15978 21680 16594
rect 21836 16114 21864 16730
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21640 15972 21692 15978
rect 21640 15914 21692 15920
rect 21732 15972 21784 15978
rect 21732 15914 21784 15920
rect 21652 13734 21680 15914
rect 21744 15609 21772 15914
rect 21730 15600 21786 15609
rect 21730 15535 21786 15544
rect 21836 15502 21864 16050
rect 22112 15978 22140 16594
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15162 21864 15438
rect 21928 15366 21956 15846
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21836 13802 21864 13874
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21836 12646 21864 13330
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21928 12424 21956 15302
rect 22006 14240 22062 14249
rect 22006 14175 22062 14184
rect 22020 14074 22048 14175
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22204 12850 22232 17598
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22296 17241 22324 17478
rect 22282 17232 22338 17241
rect 22282 17167 22338 17176
rect 22480 16794 22508 17711
rect 22572 17134 22600 17750
rect 23018 17640 23074 17649
rect 23018 17575 23074 17584
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22572 15570 22600 17070
rect 23032 16590 23060 17575
rect 23124 16658 23152 18022
rect 23216 17882 23244 18090
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23308 17542 23336 18158
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22756 15910 22784 16526
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22374 15464 22430 15473
rect 22374 15399 22430 15408
rect 22388 15162 22416 15399
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22388 14958 22416 15098
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22756 13870 22784 15846
rect 23032 15706 23060 16526
rect 23124 15910 23152 16594
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23124 15586 23152 15846
rect 23202 15736 23258 15745
rect 23202 15671 23258 15680
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 23032 15558 23152 15586
rect 22848 15162 22876 15506
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 23032 14890 23060 15558
rect 23216 15065 23244 15671
rect 23202 15056 23258 15065
rect 23202 14991 23258 15000
rect 23020 14884 23072 14890
rect 23020 14826 23072 14832
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22848 13938 22876 14418
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22388 13258 22416 13670
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 21928 12396 22140 12424
rect 21560 11886 21956 11914
rect 21732 11552 21784 11558
rect 21376 11512 21588 11540
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21376 10742 21404 11086
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21284 10560 21384 10588
rect 21356 10554 21384 10560
rect 21356 10526 21404 10554
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21100 10033 21128 10066
rect 21086 10024 21142 10033
rect 21086 9959 21142 9968
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 20640 9518 20668 9862
rect 21008 9586 21036 9862
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 8072 20668 9318
rect 20902 9072 20958 9081
rect 20720 9036 20772 9042
rect 20902 9007 20904 9016
rect 20720 8978 20772 8984
rect 20956 9007 20958 9016
rect 20996 9036 21048 9042
rect 20904 8978 20956 8984
rect 20996 8978 21048 8984
rect 20732 8809 20760 8978
rect 20718 8800 20774 8809
rect 20718 8735 20774 8744
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 8084 20772 8090
rect 20640 8044 20720 8072
rect 20720 8026 20772 8032
rect 20824 7886 20852 8570
rect 21008 8294 21036 8978
rect 21100 8430 21128 9522
rect 21192 9178 21220 10406
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20640 7410 20668 7686
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20732 6934 20760 7210
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 20732 5817 20760 6870
rect 20718 5808 20774 5817
rect 20718 5743 20774 5752
rect 20916 4321 20944 7686
rect 21008 7410 21036 8230
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21100 6458 21128 6802
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21192 5234 21220 5782
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 20902 4312 20958 4321
rect 20902 4247 20958 4256
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 3534 20760 3878
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20732 2990 20760 3470
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 21284 2689 21312 10202
rect 21376 7274 21404 10526
rect 21468 10470 21496 11290
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21560 10266 21588 11512
rect 21732 11494 21784 11500
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21652 10674 21680 10950
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21468 9586 21496 10066
rect 21560 9722 21588 10202
rect 21652 10062 21680 10610
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21652 9722 21680 9998
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21652 9042 21680 9658
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21468 8022 21496 8230
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21468 7546 21496 7822
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21468 5914 21496 7346
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21362 5536 21418 5545
rect 21362 5471 21418 5480
rect 21376 5166 21404 5471
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21468 4282 21496 4558
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 21468 4078 21496 4218
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21270 2680 21326 2689
rect 21270 2615 21326 2624
rect 20902 2544 20958 2553
rect 20902 2479 20904 2488
rect 20956 2479 20958 2488
rect 20904 2450 20956 2456
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 20718 2000 20774 2009
rect 20718 1935 20774 1944
rect 20732 480 20760 1935
rect 21376 480 21404 2314
rect 21560 610 21588 4966
rect 21744 4049 21772 11494
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 21836 8430 21864 9114
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21822 7576 21878 7585
rect 21822 7511 21824 7520
rect 21876 7511 21878 7520
rect 21824 7482 21876 7488
rect 21928 7426 21956 11886
rect 22006 11792 22062 11801
rect 22006 11727 22062 11736
rect 22020 11354 22048 11727
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22112 10674 22140 12396
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 11694 22232 12038
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22296 11354 22324 12718
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22020 9110 22048 10202
rect 22388 9625 22416 13194
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12782 22508 13126
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22558 12744 22614 12753
rect 22558 12679 22614 12688
rect 22374 9616 22430 9625
rect 22572 9602 22600 12679
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22664 10266 22692 11154
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22664 9722 22692 10202
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22572 9574 22692 9602
rect 22374 9551 22430 9560
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22296 8498 22324 8774
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22098 7984 22154 7993
rect 22098 7919 22154 7928
rect 22112 7818 22140 7919
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21836 7398 21956 7426
rect 21730 4040 21786 4049
rect 21730 3975 21786 3984
rect 21836 3720 21864 7398
rect 22020 7342 22048 7482
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21928 6746 21956 7278
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22020 6882 22048 7142
rect 22020 6866 22140 6882
rect 22020 6860 22152 6866
rect 22020 6854 22100 6860
rect 22100 6802 22152 6808
rect 21928 6718 22140 6746
rect 22006 6624 22062 6633
rect 22006 6559 22062 6568
rect 21914 6352 21970 6361
rect 21914 6287 21970 6296
rect 21928 3942 21956 6287
rect 22020 4690 22048 6559
rect 22112 6254 22140 6718
rect 22204 6458 22232 8026
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22480 7750 22508 7890
rect 22572 7886 22600 8366
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22480 7410 22508 7686
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22388 7041 22416 7142
rect 22374 7032 22430 7041
rect 22374 6967 22430 6976
rect 22572 6730 22600 7822
rect 22664 6769 22692 9574
rect 22756 7834 22784 13806
rect 22834 13288 22890 13297
rect 22834 13223 22890 13232
rect 22848 12442 22876 13223
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 23032 12594 23060 14826
rect 23202 13968 23258 13977
rect 23202 13903 23258 13912
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 23124 12714 23152 13262
rect 23112 12708 23164 12714
rect 23112 12650 23164 12656
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22848 11354 22876 12242
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 9722 22876 10406
rect 22940 10266 22968 12582
rect 23032 12566 23152 12594
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 23032 11286 23060 11766
rect 23020 11280 23072 11286
rect 23020 11222 23072 11228
rect 23032 10470 23060 11222
rect 23124 10538 23152 12566
rect 23216 10810 23244 13903
rect 23308 13462 23336 16118
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23308 12442 23336 13398
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 23400 10656 23428 20862
rect 23492 19242 23520 22607
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 18290 23520 18566
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23492 16153 23520 16934
rect 23584 16538 23612 22918
rect 23756 22568 23808 22574
rect 23756 22510 23808 22516
rect 23952 22522 23980 23122
rect 24044 22642 24072 24550
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23676 20466 23704 20810
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23676 19514 23704 19654
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23768 19394 23796 22510
rect 23952 22494 24072 22522
rect 24044 22438 24072 22494
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 23952 21729 23980 22034
rect 23938 21720 23994 21729
rect 23938 21655 23940 21664
rect 23992 21655 23994 21664
rect 23940 21626 23992 21632
rect 23952 21595 23980 21626
rect 24044 21434 24072 22374
rect 24136 21457 24164 24006
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23225 24716 24550
rect 24768 24268 24820 24274
rect 24768 24210 24820 24216
rect 24780 23526 24808 24210
rect 25134 23760 25190 23769
rect 25134 23695 25190 23704
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 24768 23520 24820 23526
rect 24768 23462 24820 23468
rect 24674 23216 24730 23225
rect 24674 23151 24730 23160
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 23676 19366 23796 19394
rect 23860 21406 24072 21434
rect 24122 21448 24178 21457
rect 23676 17921 23704 19366
rect 23662 17912 23718 17921
rect 23662 17847 23718 17856
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23768 17134 23796 17478
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 23584 16510 23704 16538
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23478 16144 23534 16153
rect 23478 16079 23534 16088
rect 23478 14920 23534 14929
rect 23478 14855 23534 14864
rect 23492 13433 23520 14855
rect 23478 13424 23534 13433
rect 23478 13359 23534 13368
rect 23216 10628 23428 10656
rect 23112 10532 23164 10538
rect 23112 10474 23164 10480
rect 23020 10464 23072 10470
rect 23018 10432 23020 10441
rect 23072 10432 23074 10441
rect 23018 10367 23074 10376
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 23018 9480 23074 9489
rect 23018 9415 23020 9424
rect 23072 9415 23074 9424
rect 23020 9386 23072 9392
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23124 8634 23152 8978
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22756 7806 22876 7834
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22756 7206 22784 7686
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22650 6760 22706 6769
rect 22560 6724 22612 6730
rect 22650 6695 22706 6704
rect 22560 6666 22612 6672
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22190 4720 22246 4729
rect 22008 4684 22060 4690
rect 22190 4655 22246 4664
rect 22008 4626 22060 4632
rect 22020 4282 22048 4626
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22112 4185 22140 4422
rect 22098 4176 22154 4185
rect 22098 4111 22154 4120
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 21916 3936 21968 3942
rect 22112 3890 22140 3946
rect 21916 3878 21968 3884
rect 21744 3692 21864 3720
rect 22020 3862 22140 3890
rect 21744 3233 21772 3692
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21730 3224 21786 3233
rect 21836 3194 21864 3538
rect 21730 3159 21786 3168
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 22020 2650 22048 3862
rect 22204 3754 22232 4655
rect 22664 4593 22692 4966
rect 22650 4584 22706 4593
rect 22650 4519 22706 4528
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22572 4146 22600 4422
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22112 3726 22232 3754
rect 22572 3738 22600 4082
rect 22560 3732 22612 3738
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 21640 2440 21692 2446
rect 21638 2408 21640 2417
rect 21692 2408 21694 2417
rect 21638 2343 21694 2352
rect 21548 604 21600 610
rect 21548 546 21600 552
rect 22112 480 22140 3726
rect 22560 3674 22612 3680
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22204 2650 22232 3130
rect 22296 2650 22324 3606
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22204 2446 22232 2586
rect 22756 2514 22784 7142
rect 22848 4865 22876 7806
rect 23216 7426 23244 10628
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23308 7834 23336 10474
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23400 9058 23428 9454
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23492 9217 23520 9318
rect 23478 9208 23534 9217
rect 23478 9143 23534 9152
rect 23400 9030 23520 9058
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23400 8430 23428 8774
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23492 7993 23520 9030
rect 23478 7984 23534 7993
rect 23478 7919 23534 7928
rect 23308 7806 23520 7834
rect 23032 7398 23244 7426
rect 23032 6361 23060 7398
rect 23110 7304 23166 7313
rect 23110 7239 23166 7248
rect 23018 6352 23074 6361
rect 23018 6287 23074 6296
rect 22834 4856 22890 4865
rect 22890 4814 22968 4842
rect 23124 4826 23152 7239
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23216 7002 23244 7142
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23216 6322 23244 6938
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23308 5846 23336 6734
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 23294 5672 23350 5681
rect 23294 5607 23350 5616
rect 23204 5092 23256 5098
rect 23204 5034 23256 5040
rect 22834 4791 22890 4800
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22848 4078 22876 4422
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22940 3942 22968 4814
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 23124 3398 23152 4558
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23124 3194 23152 3334
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23216 2582 23244 5034
rect 23308 4826 23336 5607
rect 23296 4820 23348 4826
rect 23296 4762 23348 4768
rect 23308 4282 23336 4762
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 23204 2576 23256 2582
rect 23204 2518 23256 2524
rect 23400 2530 23428 6054
rect 23492 5846 23520 7806
rect 23584 7313 23612 16390
rect 23676 11558 23704 16510
rect 23860 16454 23888 21406
rect 24122 21383 24178 21392
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23952 17882 23980 21286
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24030 19952 24086 19961
rect 24030 19887 24086 19896
rect 24044 19514 24072 19887
rect 24136 19786 24164 20946
rect 24228 19825 24256 22646
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24584 21412 24636 21418
rect 24584 21354 24636 21360
rect 24596 21185 24624 21354
rect 24582 21176 24638 21185
rect 24582 21111 24638 21120
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24584 20256 24636 20262
rect 24584 20198 24636 20204
rect 24398 19952 24454 19961
rect 24398 19887 24400 19896
rect 24452 19887 24454 19896
rect 24400 19858 24452 19864
rect 24596 19854 24624 20198
rect 24584 19848 24636 19854
rect 24214 19816 24270 19825
rect 24124 19780 24176 19786
rect 24584 19790 24636 19796
rect 24214 19751 24270 19760
rect 24124 19722 24176 19728
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24122 19544 24178 19553
rect 24032 19508 24084 19514
rect 24289 19536 24585 19556
rect 24122 19479 24178 19488
rect 24032 19450 24084 19456
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 24044 19174 24072 19314
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 24044 18086 24072 19110
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 23940 17060 23992 17066
rect 23940 17002 23992 17008
rect 23952 16726 23980 17002
rect 24044 16794 24072 17682
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23940 16720 23992 16726
rect 23940 16662 23992 16668
rect 24136 16640 24164 19479
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 24228 18873 24256 19110
rect 24504 18902 24532 19314
rect 24688 19145 24716 21830
rect 24780 21078 24808 23462
rect 25056 23361 25084 23598
rect 25042 23352 25098 23361
rect 25042 23287 25098 23296
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 25056 22273 25084 22510
rect 25042 22264 25098 22273
rect 25042 22199 25098 22208
rect 24860 21344 24912 21350
rect 24860 21286 24912 21292
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24768 20052 24820 20058
rect 24872 20040 24900 21286
rect 24950 21040 25006 21049
rect 24950 20975 25006 20984
rect 24820 20012 24900 20040
rect 24768 19994 24820 20000
rect 24674 19136 24730 19145
rect 24674 19071 24730 19080
rect 24780 18970 24808 19994
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24872 19378 24900 19790
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24492 18896 24544 18902
rect 24214 18864 24270 18873
rect 24492 18838 24544 18844
rect 24214 18799 24270 18808
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 17882 24716 18566
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24228 16998 24256 17614
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17338 24716 17818
rect 24766 17504 24822 17513
rect 24766 17439 24822 17448
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24398 16960 24454 16969
rect 24398 16895 24454 16904
rect 24412 16658 24440 16895
rect 24490 16824 24546 16833
rect 24546 16768 24716 16776
rect 24490 16759 24492 16768
rect 24544 16748 24716 16768
rect 24492 16730 24544 16736
rect 24400 16652 24452 16658
rect 24044 16612 24164 16640
rect 24228 16612 24400 16640
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 24044 16250 24072 16612
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23846 16144 23902 16153
rect 23756 16108 23808 16114
rect 23846 16079 23902 16088
rect 23756 16050 23808 16056
rect 23768 13258 23796 16050
rect 23860 14822 23888 16079
rect 24044 16046 24072 16186
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 24136 15910 24164 16458
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24136 15337 24164 15846
rect 24228 15706 24256 16612
rect 24400 16594 24452 16600
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16250 24716 16748
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24596 15706 24624 16050
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24122 15328 24178 15337
rect 24122 15263 24178 15272
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24122 15192 24178 15201
rect 24289 15184 24585 15204
rect 24122 15127 24178 15136
rect 24780 15144 24808 17439
rect 24964 15638 24992 20975
rect 25042 19408 25098 19417
rect 25042 19343 25098 19352
rect 25056 19310 25084 19343
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 25148 18834 25176 23695
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25240 20913 25268 23462
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25424 22409 25452 23054
rect 25410 22400 25466 22409
rect 25410 22335 25466 22344
rect 25516 21593 25544 27520
rect 26160 25294 26188 27520
rect 26896 25430 26924 27520
rect 26884 25424 26936 25430
rect 26884 25366 26936 25372
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 27540 24585 27568 27520
rect 27526 24576 27582 24585
rect 27526 24511 27582 24520
rect 25686 23760 25742 23769
rect 25686 23695 25742 23704
rect 25502 21584 25558 21593
rect 25502 21519 25558 21528
rect 25226 20904 25282 20913
rect 25226 20839 25282 20848
rect 25228 19304 25280 19310
rect 25226 19272 25228 19281
rect 25280 19272 25282 19281
rect 25226 19207 25282 19216
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25516 19009 25544 19178
rect 25502 19000 25558 19009
rect 25502 18935 25558 18944
rect 25502 18864 25558 18873
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25412 18828 25464 18834
rect 25502 18799 25558 18808
rect 25412 18770 25464 18776
rect 25056 18068 25084 18770
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25240 18426 25268 18702
rect 25228 18420 25280 18426
rect 25228 18362 25280 18368
rect 25136 18080 25188 18086
rect 25056 18040 25136 18068
rect 25136 18022 25188 18028
rect 24952 15632 25004 15638
rect 24952 15574 25004 15580
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 24860 15156 24912 15162
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23846 14648 23902 14657
rect 23952 14618 23980 14962
rect 24136 14958 24164 15127
rect 24780 15116 24860 15144
rect 24860 15098 24912 15104
rect 25056 15094 25084 15506
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 23846 14583 23902 14592
rect 23940 14612 23992 14618
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23768 12442 23796 13194
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23768 11898 23796 12378
rect 23860 12345 23888 14583
rect 23940 14554 23992 14560
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 23952 13870 23980 14282
rect 24044 14278 24072 14758
rect 24320 14362 24348 14758
rect 25042 14512 25098 14521
rect 25042 14447 25044 14456
rect 25096 14447 25098 14456
rect 25044 14418 25096 14424
rect 24228 14334 24348 14362
rect 24032 14272 24084 14278
rect 24030 14240 24032 14249
rect 24084 14240 24086 14249
rect 24030 14175 24086 14184
rect 24228 14056 24256 14334
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24768 14068 24820 14074
rect 24228 14028 24348 14056
rect 23940 13864 23992 13870
rect 23992 13824 24072 13852
rect 23940 13806 23992 13812
rect 24044 13512 24072 13824
rect 24320 13530 24348 14028
rect 24768 14010 24820 14016
rect 24780 13802 24808 14010
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24768 13796 24820 13802
rect 24768 13738 24820 13744
rect 24308 13524 24360 13530
rect 24044 13484 24164 13512
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24044 12918 24072 13330
rect 24032 12912 24084 12918
rect 24030 12880 24032 12889
rect 24084 12880 24086 12889
rect 24136 12850 24164 13484
rect 24308 13466 24360 13472
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24030 12815 24086 12824
rect 24124 12844 24176 12850
rect 23846 12336 23902 12345
rect 23846 12271 23902 12280
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23768 11354 23796 11834
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23570 7304 23626 7313
rect 23570 7239 23626 7248
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23584 5710 23612 6598
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23492 2990 23520 5510
rect 23584 5370 23612 5646
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23584 4622 23612 5170
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23584 4146 23612 4558
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23492 2650 23520 2926
rect 23570 2680 23626 2689
rect 23480 2644 23532 2650
rect 23570 2615 23626 2624
rect 23480 2586 23532 2592
rect 22744 2508 22796 2514
rect 23400 2502 23520 2530
rect 22744 2450 22796 2456
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22742 1864 22798 1873
rect 22742 1799 22798 1808
rect 22756 480 22784 1799
rect 23492 480 23520 2502
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2318 0 2374 480
rect 2962 0 3018 480
rect 3698 0 3754 480
rect 4342 0 4398 480
rect 4986 0 5042 480
rect 5722 0 5778 480
rect 6366 0 6422 480
rect 7102 0 7158 480
rect 7746 0 7802 480
rect 8390 0 8446 480
rect 9126 0 9182 480
rect 9770 0 9826 480
rect 10506 0 10562 480
rect 11150 0 11206 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13174 0 13230 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15290 0 15346 480
rect 15934 0 15990 480
rect 16578 0 16634 480
rect 17314 0 17370 480
rect 17958 0 18014 480
rect 18694 0 18750 480
rect 19338 0 19394 480
rect 20074 0 20130 480
rect 20718 0 20774 480
rect 21362 0 21418 480
rect 22098 0 22154 480
rect 22742 0 22798 480
rect 23478 0 23534 480
rect 23584 377 23612 2615
rect 23676 2514 23704 10406
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23860 9722 23888 10202
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 23754 9480 23810 9489
rect 23754 9415 23810 9424
rect 23768 7857 23796 9415
rect 23952 9058 23980 10746
rect 24044 9178 24072 12815
rect 24124 12786 24176 12792
rect 24136 12374 24164 12786
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24214 12336 24270 12345
rect 24214 12271 24270 12280
rect 24228 11762 24256 12271
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24228 11642 24256 11698
rect 24136 11614 24256 11642
rect 24136 10305 24164 11614
rect 24596 11558 24624 11698
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24228 10606 24256 11494
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24122 10296 24178 10305
rect 24228 10266 24256 10406
rect 24320 10266 24348 10610
rect 24122 10231 24178 10240
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24122 9752 24178 9761
rect 24289 9744 24585 9764
rect 24122 9687 24178 9696
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 23860 9030 23980 9058
rect 23860 8945 23888 9030
rect 23846 8936 23902 8945
rect 23846 8871 23902 8880
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23754 7848 23810 7857
rect 23754 7783 23810 7792
rect 23860 7018 23888 8774
rect 23952 8090 23980 8842
rect 24044 8634 24072 9114
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 24136 8480 24164 9687
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 24044 8452 24164 8480
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23952 7342 23980 8026
rect 24044 7449 24072 8452
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 24136 7750 24164 8298
rect 24228 8265 24256 9318
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24214 8256 24270 8265
rect 24214 8191 24270 8200
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24030 7440 24086 7449
rect 24030 7375 24086 7384
rect 23940 7336 23992 7342
rect 23992 7296 24072 7324
rect 23940 7278 23992 7284
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 23768 6990 23888 7018
rect 23768 5914 23796 6990
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23860 6458 23888 6802
rect 23952 6662 23980 7142
rect 24044 6798 24072 7296
rect 24136 7206 24164 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23952 6338 23980 6598
rect 24044 6390 24072 6734
rect 23860 6310 23980 6338
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23860 5574 23888 6310
rect 24136 6202 24164 7142
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24044 6174 24164 6202
rect 23940 5840 23992 5846
rect 23940 5782 23992 5788
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 23860 5166 23888 5510
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 23860 4758 23888 5102
rect 23848 4752 23900 4758
rect 23848 4694 23900 4700
rect 23860 4162 23888 4694
rect 23768 4134 23888 4162
rect 23768 4078 23796 4134
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 2553 23796 3878
rect 23860 3738 23888 3946
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23952 3670 23980 5782
rect 24044 5710 24072 6174
rect 24596 5914 24624 6258
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24044 5370 24072 5646
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24124 5092 24176 5098
rect 24124 5034 24176 5040
rect 24136 4486 24164 5034
rect 24688 4826 24716 13330
rect 24780 13326 24808 13738
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24872 12986 24900 13806
rect 25056 13530 25084 14418
rect 25148 13734 25176 18022
rect 25240 17882 25268 18362
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25240 16726 25268 17818
rect 25424 17610 25452 18770
rect 25412 17604 25464 17610
rect 25412 17546 25464 17552
rect 25318 16824 25374 16833
rect 25318 16759 25374 16768
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 25240 16250 25268 16662
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25228 16040 25280 16046
rect 25226 16008 25228 16017
rect 25280 16008 25282 16017
rect 25226 15943 25282 15952
rect 25332 14618 25360 16759
rect 25320 14612 25372 14618
rect 25320 14554 25372 14560
rect 25226 13968 25282 13977
rect 25226 13903 25282 13912
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 24952 12708 25004 12714
rect 24952 12650 25004 12656
rect 24964 12442 24992 12650
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24860 11620 24912 11626
rect 24860 11562 24912 11568
rect 24872 10674 24900 11562
rect 24964 11354 24992 11698
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24964 10130 24992 11290
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24964 9722 24992 10066
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24964 9586 24992 9658
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24768 9036 24820 9042
rect 24820 8996 24900 9024
rect 24768 8978 24820 8984
rect 24766 8936 24822 8945
rect 24766 8871 24822 8880
rect 24780 6338 24808 8871
rect 24872 8090 24900 8996
rect 24964 8634 24992 9522
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 24780 6310 24900 6338
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24780 4826 24808 6190
rect 24872 6118 24900 6310
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24872 5522 24900 6054
rect 25056 5681 25084 6734
rect 25042 5672 25098 5681
rect 25042 5607 25098 5616
rect 24872 5494 24992 5522
rect 24860 5024 24912 5030
rect 24860 4966 24912 4972
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24872 4622 24900 4966
rect 24964 4758 24992 5494
rect 25042 4856 25098 4865
rect 25042 4791 25044 4800
rect 25096 4791 25098 4800
rect 25044 4762 25096 4768
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 23940 3664 23992 3670
rect 23940 3606 23992 3612
rect 24136 3466 24164 4422
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24964 4282 24992 4694
rect 24952 4276 25004 4282
rect 24952 4218 25004 4224
rect 24766 4176 24822 4185
rect 24766 4111 24822 4120
rect 24398 4040 24454 4049
rect 24398 3975 24454 3984
rect 24412 3738 24440 3975
rect 24674 3768 24730 3777
rect 24400 3732 24452 3738
rect 24228 3692 24400 3720
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 24136 3194 24164 3402
rect 24228 3194 24256 3692
rect 24674 3703 24730 3712
rect 24400 3674 24452 3680
rect 24688 3670 24716 3703
rect 24676 3664 24728 3670
rect 24676 3606 24728 3612
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3606
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 23846 3088 23902 3097
rect 23846 3023 23902 3032
rect 23754 2544 23810 2553
rect 23664 2508 23716 2514
rect 23754 2479 23810 2488
rect 23664 2450 23716 2456
rect 23860 2417 23888 3023
rect 23940 2916 23992 2922
rect 23940 2858 23992 2864
rect 23846 2408 23902 2417
rect 23846 2343 23902 2352
rect 23952 1601 23980 2858
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23938 1592 23994 1601
rect 23938 1527 23994 1536
rect 24124 604 24176 610
rect 24124 546 24176 552
rect 24136 480 24164 546
rect 24780 480 24808 4111
rect 25056 4026 25084 4762
rect 25148 4622 25176 12922
rect 25240 10810 25268 13903
rect 25320 12368 25372 12374
rect 25320 12310 25372 12316
rect 25332 11898 25360 12310
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25318 11248 25374 11257
rect 25318 11183 25320 11192
rect 25372 11183 25374 11192
rect 25320 11154 25372 11160
rect 25332 10810 25360 11154
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25424 9704 25452 17546
rect 25516 17218 25544 18799
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25608 17338 25636 17682
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25516 17190 25636 17218
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25516 16658 25544 17070
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25504 15972 25556 15978
rect 25504 15914 25556 15920
rect 25516 15473 25544 15914
rect 25502 15464 25558 15473
rect 25502 15399 25558 15408
rect 25424 9676 25544 9704
rect 25410 9616 25466 9625
rect 25410 9551 25412 9560
rect 25464 9551 25466 9560
rect 25412 9522 25464 9528
rect 25318 7032 25374 7041
rect 25318 6967 25374 6976
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 24964 3998 25084 4026
rect 24964 3738 24992 3998
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 25056 3534 25084 3878
rect 25148 3738 25176 4558
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25332 2514 25360 6967
rect 25516 5137 25544 9676
rect 25608 5778 25636 17190
rect 25700 11354 25728 23695
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 26160 15178 26188 16594
rect 26160 15162 26280 15178
rect 26160 15156 26292 15162
rect 26160 15150 26240 15156
rect 26240 15098 26292 15104
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 26068 14074 26096 14214
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25596 5772 25648 5778
rect 25596 5714 25648 5720
rect 25608 5370 25636 5714
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25502 5128 25558 5137
rect 25502 5063 25558 5072
rect 25516 4672 25544 5063
rect 25424 4644 25544 4672
rect 25424 3194 25452 4644
rect 25502 4584 25558 4593
rect 25502 4519 25558 4528
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 25424 2990 25452 3130
rect 25412 2984 25464 2990
rect 25412 2926 25464 2932
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25516 480 25544 4519
rect 25608 3641 25636 5306
rect 26068 4321 26096 13670
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26054 4312 26110 4321
rect 26054 4247 26110 4256
rect 25594 3632 25650 3641
rect 25594 3567 25650 3576
rect 26160 480 26188 5510
rect 26884 3120 26936 3126
rect 26884 3062 26936 3068
rect 26896 480 26924 3062
rect 27528 2372 27580 2378
rect 27528 2314 27580 2320
rect 27540 480 27568 2314
rect 23570 368 23626 377
rect 23570 303 23626 312
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25502 0 25558 480
rect 26146 0 26202 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 24582 27648 24638 27704
rect 938 23024 994 23080
rect 386 15408 442 15464
rect 294 7384 350 7440
rect 570 6976 626 7032
rect 2962 22480 3018 22536
rect 4066 20984 4122 21040
rect 3698 19896 3754 19952
rect 1582 19216 1638 19272
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 4986 22616 5042 22672
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 7746 24248 7802 24304
rect 7102 23568 7158 23624
rect 6366 23432 6422 23488
rect 7746 23432 7802 23488
rect 5998 20032 6054 20088
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 9126 24656 9182 24712
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10690 24248 10746 24304
rect 9770 23976 9826 24032
rect 9310 23568 9366 23624
rect 10782 24112 10838 24168
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 11886 24248 11942 24304
rect 12714 24792 12770 24848
rect 12622 23704 12678 23760
rect 10874 22208 10930 22264
rect 11242 23160 11298 23216
rect 12346 22616 12402 22672
rect 11886 22344 11942 22400
rect 9218 20984 9274 21040
rect 7838 20324 7894 20360
rect 7838 20304 7840 20324
rect 7840 20304 7892 20324
rect 7892 20304 7894 20324
rect 7838 20052 7894 20088
rect 7838 20032 7840 20052
rect 7840 20032 7892 20052
rect 7892 20032 7894 20052
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9310 19760 9366 19816
rect 4342 18944 4398 19000
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 9310 19080 9366 19136
rect 9586 19080 9642 19136
rect 10598 19236 10654 19272
rect 10598 19216 10600 19236
rect 10600 19216 10652 19236
rect 10652 19216 10654 19236
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18944 10194 19000
rect 9494 17060 9550 17096
rect 9494 17040 9496 17060
rect 9496 17040 9548 17060
rect 9548 17040 9550 17060
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 4066 13912 4122 13968
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 10046 15952 10102 16008
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 3698 8336 3754 8392
rect 2318 5616 2374 5672
rect 1398 3984 1454 4040
rect 1582 2488 1638 2544
rect 2962 5208 3018 5264
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 4342 6704 4398 6760
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 7746 11056 7802 11112
rect 7654 5072 7710 5128
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6366 3848 6422 3904
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 4986 3032 5042 3088
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5722 1400 5778 1456
rect 7102 3576 7158 3632
rect 9862 7792 9918 7848
rect 9586 4156 9588 4176
rect 9588 4156 9640 4176
rect 9640 4156 9642 4176
rect 9586 4120 9642 4156
rect 9770 5480 9826 5536
rect 8390 2896 8446 2952
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 11242 20440 11298 20496
rect 12346 21120 12402 21176
rect 12438 21004 12494 21040
rect 12438 20984 12440 21004
rect 12440 20984 12492 21004
rect 12492 20984 12494 21004
rect 12714 21528 12770 21584
rect 10966 18264 11022 18320
rect 11610 18128 11666 18184
rect 10874 15816 10930 15872
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10230 14356 10232 14376
rect 10232 14356 10284 14376
rect 10284 14356 10286 14376
rect 10230 14320 10286 14356
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10782 15428 10838 15464
rect 10782 15408 10784 15428
rect 10784 15408 10836 15428
rect 10836 15408 10838 15428
rect 10782 15136 10838 15192
rect 11242 15408 11298 15464
rect 11702 16652 11758 16688
rect 11702 16632 11704 16652
rect 11704 16632 11756 16652
rect 11756 16632 11758 16652
rect 11334 15136 11390 15192
rect 10782 12824 10838 12880
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10782 11600 10838 11656
rect 12254 18536 12310 18592
rect 12898 18128 12954 18184
rect 12898 17076 12900 17096
rect 12900 17076 12952 17096
rect 12952 17076 12954 17096
rect 12898 17040 12954 17076
rect 13266 24148 13268 24168
rect 13268 24148 13320 24168
rect 13320 24148 13322 24168
rect 13266 24112 13322 24148
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14554 24792 14610 24848
rect 13450 22480 13506 22536
rect 13634 22480 13690 22536
rect 14094 23024 14150 23080
rect 14002 20848 14058 20904
rect 13358 20032 13414 20088
rect 13634 18128 13690 18184
rect 13174 17040 13230 17096
rect 12990 16940 12992 16960
rect 12992 16940 13044 16960
rect 13044 16940 13046 16960
rect 12990 16904 13046 16940
rect 12622 16768 12678 16824
rect 13174 16632 13230 16688
rect 11978 12436 12034 12472
rect 11978 12416 11980 12436
rect 11980 12416 12032 12436
rect 12032 12416 12034 12436
rect 10966 10376 11022 10432
rect 10046 3848 10102 3904
rect 10782 9288 10838 9344
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10598 7384 10654 7440
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 11334 8372 11336 8392
rect 11336 8372 11388 8392
rect 11388 8372 11390 8392
rect 11334 8336 11390 8372
rect 10874 7384 10930 7440
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10782 5652 10784 5672
rect 10784 5652 10836 5672
rect 10836 5652 10838 5672
rect 10782 5616 10838 5652
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3576 10194 3632
rect 10782 3440 10838 3496
rect 10874 2760 10930 2816
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10874 2644 10930 2680
rect 10874 2624 10876 2644
rect 10876 2624 10928 2644
rect 10928 2624 10930 2644
rect 11334 7656 11390 7712
rect 11058 5616 11114 5672
rect 11150 3884 11152 3904
rect 11152 3884 11204 3904
rect 11204 3884 11206 3904
rect 11150 3848 11206 3884
rect 11150 3596 11206 3632
rect 11150 3576 11152 3596
rect 11152 3576 11204 3596
rect 11204 3576 11206 3596
rect 11058 3032 11114 3088
rect 11334 6024 11390 6080
rect 11610 4936 11666 4992
rect 11334 4020 11336 4040
rect 11336 4020 11388 4040
rect 11388 4020 11390 4040
rect 11334 3984 11390 4020
rect 11518 3984 11574 4040
rect 11426 3168 11482 3224
rect 11426 3068 11428 3088
rect 11428 3068 11480 3088
rect 11480 3068 11482 3088
rect 10782 1672 10838 1728
rect 11426 3032 11482 3068
rect 12254 12980 12310 13016
rect 12254 12960 12256 12980
rect 12256 12960 12308 12980
rect 12308 12960 12310 12980
rect 12438 12824 12494 12880
rect 12898 13388 12954 13424
rect 12898 13368 12900 13388
rect 12900 13368 12952 13388
rect 12952 13368 12954 13388
rect 13174 15408 13230 15464
rect 13082 13232 13138 13288
rect 12530 12280 12586 12336
rect 12438 11636 12440 11656
rect 12440 11636 12492 11656
rect 12492 11636 12494 11656
rect 12438 11600 12494 11636
rect 12438 10240 12494 10296
rect 12898 10648 12954 10704
rect 12438 7792 12494 7848
rect 12438 5752 12494 5808
rect 12346 5480 12402 5536
rect 12898 9324 12900 9344
rect 12900 9324 12952 9344
rect 12952 9324 12954 9344
rect 12898 9288 12954 9324
rect 12898 8880 12954 8936
rect 12806 6976 12862 7032
rect 12622 3712 12678 3768
rect 13174 12824 13230 12880
rect 14278 18572 14280 18592
rect 14280 18572 14332 18592
rect 14332 18572 14334 18592
rect 14278 18536 14334 18572
rect 14094 17740 14150 17776
rect 14094 17720 14096 17740
rect 14096 17720 14148 17740
rect 14148 17720 14150 17740
rect 13910 17584 13966 17640
rect 13634 16768 13690 16824
rect 13450 15544 13506 15600
rect 13266 11600 13322 11656
rect 12530 2896 12586 2952
rect 11610 1944 11666 2000
rect 13266 8472 13322 8528
rect 13450 6704 13506 6760
rect 13266 6196 13268 6216
rect 13268 6196 13320 6216
rect 13320 6196 13322 6216
rect 13266 6160 13322 6196
rect 13266 5072 13322 5128
rect 13818 14864 13874 14920
rect 13726 13776 13782 13832
rect 14278 16088 14334 16144
rect 14186 15680 14242 15736
rect 14922 24656 14978 24712
rect 15474 24792 15530 24848
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14554 23296 14610 23352
rect 14462 19352 14518 19408
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15290 22480 15346 22536
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15934 24656 15990 24712
rect 15842 24404 15898 24440
rect 15842 24384 15844 24404
rect 15844 24384 15896 24404
rect 15896 24384 15898 24404
rect 15658 23432 15714 23488
rect 15566 21972 15568 21992
rect 15568 21972 15620 21992
rect 15620 21972 15622 21992
rect 15566 21936 15622 21972
rect 14646 21120 14702 21176
rect 14002 13096 14058 13152
rect 13634 11328 13690 11384
rect 14002 10412 14004 10432
rect 14004 10412 14056 10432
rect 14056 10412 14058 10432
rect 14002 10376 14058 10412
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14738 19896 14794 19952
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14830 18828 14886 18864
rect 14830 18808 14832 18828
rect 14832 18808 14884 18828
rect 14884 18808 14886 18828
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14738 17584 14794 17640
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15382 17040 15438 17096
rect 15290 16904 15346 16960
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14646 13640 14702 13696
rect 14646 13504 14702 13560
rect 14462 12552 14518 12608
rect 14462 11056 14518 11112
rect 14462 10920 14518 10976
rect 13910 7656 13966 7712
rect 13726 7384 13782 7440
rect 13818 3576 13874 3632
rect 14370 7828 14372 7848
rect 14372 7828 14424 7848
rect 14424 7828 14426 7848
rect 14370 7792 14426 7828
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15474 15408 15530 15464
rect 15842 22208 15898 22264
rect 15842 19760 15898 19816
rect 15750 19352 15806 19408
rect 15750 16652 15806 16688
rect 15750 16632 15752 16652
rect 15752 16632 15804 16652
rect 15804 16632 15806 16652
rect 15750 16496 15806 16552
rect 15382 14048 15438 14104
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14830 12552 14886 12608
rect 15106 12180 15108 12200
rect 15108 12180 15160 12200
rect 15160 12180 15162 12200
rect 15106 12144 15162 12180
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14738 11192 14794 11248
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14830 10512 14886 10568
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15474 8608 15530 8664
rect 15382 7928 15438 7984
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14738 6060 14740 6080
rect 14740 6060 14792 6080
rect 14792 6060 14794 6080
rect 14738 6024 14794 6060
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14278 4548 14334 4584
rect 14278 4528 14280 4548
rect 14280 4528 14332 4548
rect 14332 4528 14334 4548
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15566 3848 15622 3904
rect 13634 2896 13690 2952
rect 13726 2372 13782 2408
rect 13726 2352 13728 2372
rect 13728 2352 13780 2372
rect 13780 2352 13782 2372
rect 15198 3576 15254 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14554 3168 14610 3224
rect 14462 1808 14518 1864
rect 15290 2760 15346 2816
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14830 1536 14886 1592
rect 15842 15272 15898 15328
rect 15750 15000 15806 15056
rect 15750 13812 15752 13832
rect 15752 13812 15804 13832
rect 15804 13812 15806 13832
rect 15750 13776 15806 13812
rect 15934 12280 15990 12336
rect 16210 20324 16266 20360
rect 16210 20304 16212 20324
rect 16212 20304 16264 20324
rect 16264 20304 16266 20324
rect 16394 23296 16450 23352
rect 16946 23468 16948 23488
rect 16948 23468 17000 23488
rect 17000 23468 17002 23488
rect 16946 23432 17002 23468
rect 16394 20168 16450 20224
rect 16578 20032 16634 20088
rect 17038 22072 17094 22128
rect 17038 20304 17094 20360
rect 16394 18164 16396 18184
rect 16396 18164 16448 18184
rect 16448 18164 16450 18184
rect 16394 18128 16450 18164
rect 16394 14864 16450 14920
rect 17222 19896 17278 19952
rect 17314 18808 17370 18864
rect 17038 14728 17094 14784
rect 16946 14456 17002 14512
rect 17130 14356 17132 14376
rect 17132 14356 17184 14376
rect 17184 14356 17186 14376
rect 17130 14320 17186 14356
rect 16486 13504 16542 13560
rect 16118 12688 16174 12744
rect 15934 11192 15990 11248
rect 16210 12316 16212 12336
rect 16212 12316 16264 12336
rect 16264 12316 16266 12336
rect 16210 12280 16266 12316
rect 16118 10104 16174 10160
rect 16026 9968 16082 10024
rect 15750 8064 15806 8120
rect 15934 7792 15990 7848
rect 15842 7112 15898 7168
rect 16210 8064 16266 8120
rect 16210 7520 16266 7576
rect 15842 5072 15898 5128
rect 16118 4256 16174 4312
rect 15934 3984 15990 4040
rect 16762 12164 16818 12200
rect 16762 12144 16764 12164
rect 16764 12144 16816 12164
rect 16816 12144 16818 12164
rect 17406 18028 17408 18048
rect 17408 18028 17460 18048
rect 17460 18028 17462 18048
rect 17406 17992 17462 18028
rect 17774 23160 17830 23216
rect 17130 12144 17186 12200
rect 16394 5344 16450 5400
rect 16854 9424 16910 9480
rect 16762 5616 16818 5672
rect 16578 3712 16634 3768
rect 16302 2760 16358 2816
rect 16118 1400 16174 1456
rect 16670 3440 16726 3496
rect 17038 5616 17094 5672
rect 17038 4664 17094 4720
rect 17038 2624 17094 2680
rect 16762 2216 16818 2272
rect 17314 11464 17370 11520
rect 17314 10240 17370 10296
rect 17682 15136 17738 15192
rect 17498 13368 17554 13424
rect 17498 12008 17554 12064
rect 17406 8880 17462 8936
rect 18142 20168 18198 20224
rect 18510 22380 18512 22400
rect 18512 22380 18564 22400
rect 18564 22380 18566 22400
rect 18510 22344 18566 22380
rect 18510 22208 18566 22264
rect 18510 20712 18566 20768
rect 18418 19896 18474 19952
rect 18326 19352 18382 19408
rect 18418 19252 18420 19272
rect 18420 19252 18472 19272
rect 18472 19252 18474 19272
rect 18418 19216 18474 19252
rect 18050 18808 18106 18864
rect 18602 17992 18658 18048
rect 17958 16632 18014 16688
rect 18510 15852 18512 15872
rect 18512 15852 18564 15872
rect 18564 15852 18566 15872
rect 18510 15816 18566 15852
rect 18418 15544 18474 15600
rect 18510 15272 18566 15328
rect 18326 15000 18382 15056
rect 18326 13776 18382 13832
rect 17866 12824 17922 12880
rect 17682 11600 17738 11656
rect 17682 10260 17738 10296
rect 17682 10240 17684 10260
rect 17684 10240 17736 10260
rect 17736 10240 17738 10260
rect 17958 11056 18014 11112
rect 17866 9560 17922 9616
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 21086 24556 21088 24576
rect 21088 24556 21140 24576
rect 21140 24556 21142 24576
rect 18878 24112 18934 24168
rect 18786 20204 18788 20224
rect 18788 20204 18840 20224
rect 18840 20204 18842 20224
rect 18786 20168 18842 20204
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19982 21528 20038 21584
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 18878 18808 18934 18864
rect 18694 17196 18750 17232
rect 18694 17176 18696 17196
rect 18696 17176 18748 17196
rect 18748 17176 18750 17196
rect 18786 15952 18842 16008
rect 18786 15000 18842 15056
rect 19338 17992 19394 18048
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19982 17584 20038 17640
rect 19246 15544 19302 15600
rect 18970 15272 19026 15328
rect 18694 12960 18750 13016
rect 18878 12844 18934 12880
rect 18878 12824 18880 12844
rect 18880 12824 18932 12844
rect 18932 12824 18934 12844
rect 18602 10648 18658 10704
rect 17958 9016 18014 9072
rect 17866 8744 17922 8800
rect 17498 8472 17554 8528
rect 18602 7792 18658 7848
rect 17958 7112 18014 7168
rect 17866 6976 17922 7032
rect 18142 6860 18198 6896
rect 18142 6840 18144 6860
rect 18144 6840 18196 6860
rect 18196 6840 18198 6860
rect 18878 11192 18934 11248
rect 19430 15680 19486 15736
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20074 15952 20130 16008
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19614 14884 19670 14920
rect 19614 14864 19616 14884
rect 19616 14864 19668 14884
rect 19668 14864 19670 14884
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19522 14320 19578 14376
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19338 11500 19340 11520
rect 19340 11500 19392 11520
rect 19392 11500 19394 11520
rect 19338 11464 19394 11500
rect 19154 10920 19210 10976
rect 19614 13232 19670 13288
rect 20074 13504 20130 13560
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19706 11056 19762 11112
rect 20626 22208 20682 22264
rect 20350 21004 20406 21040
rect 20350 20984 20352 21004
rect 20352 20984 20404 21004
rect 20404 20984 20406 21004
rect 20258 20712 20314 20768
rect 21086 24520 21142 24556
rect 20810 24248 20866 24304
rect 21178 23296 21234 23352
rect 21546 24384 21602 24440
rect 20810 22616 20866 22672
rect 20902 20848 20958 20904
rect 20810 20324 20866 20360
rect 20810 20304 20812 20324
rect 20812 20304 20864 20324
rect 20864 20304 20866 20324
rect 21086 20748 21088 20768
rect 21088 20748 21140 20768
rect 21140 20748 21142 20768
rect 21086 20712 21142 20748
rect 20994 20440 21050 20496
rect 20350 18284 20406 18320
rect 20350 18264 20352 18284
rect 20352 18264 20404 18284
rect 20404 18264 20406 18284
rect 18694 7248 18750 7304
rect 18694 5344 18750 5400
rect 18786 5092 18842 5128
rect 18786 5072 18788 5092
rect 18788 5072 18840 5092
rect 18840 5072 18842 5092
rect 18694 4972 18696 4992
rect 18696 4972 18748 4992
rect 18748 4972 18750 4992
rect 18694 4936 18750 4972
rect 18050 3188 18106 3224
rect 18050 3168 18052 3188
rect 18052 3168 18104 3188
rect 18104 3168 18106 3188
rect 17958 3032 18014 3088
rect 17314 1672 17370 1728
rect 17130 856 17186 912
rect 18694 2896 18750 2952
rect 18510 2796 18512 2816
rect 18512 2796 18564 2816
rect 18564 2796 18566 2816
rect 18510 2760 18566 2796
rect 19430 9596 19432 9616
rect 19432 9596 19484 9616
rect 19484 9596 19486 9616
rect 19430 9560 19486 9596
rect 19338 4528 19394 4584
rect 19246 3984 19302 4040
rect 19062 2352 19118 2408
rect 19062 1400 19118 1456
rect 20074 10376 20130 10432
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20166 10260 20222 10296
rect 20166 10240 20168 10260
rect 20168 10240 20220 10260
rect 20220 10240 20222 10260
rect 20074 9172 20130 9208
rect 20074 9152 20076 9172
rect 20076 9152 20128 9172
rect 20128 9152 20130 9172
rect 19982 8472 20038 8528
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20626 16904 20682 16960
rect 20534 16768 20590 16824
rect 20902 19624 20958 19680
rect 21270 22516 21272 22536
rect 21272 22516 21324 22536
rect 21324 22516 21326 22536
rect 21270 22480 21326 22516
rect 20994 19488 21050 19544
rect 21086 19352 21142 19408
rect 21454 22480 21510 22536
rect 21638 20848 21694 20904
rect 21362 19216 21418 19272
rect 21178 18808 21234 18864
rect 21086 18672 21142 18728
rect 21270 17992 21326 18048
rect 23386 26560 23442 26616
rect 23294 26016 23350 26072
rect 22282 24248 22338 24304
rect 21822 21140 21878 21176
rect 21822 21120 21824 21140
rect 21824 21120 21876 21140
rect 21876 21120 21878 21140
rect 22282 22208 22338 22264
rect 22742 22344 22798 22400
rect 22650 22072 22706 22128
rect 23662 25336 23718 25392
rect 23478 24384 23534 24440
rect 24766 27104 24822 27160
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24582 24792 24638 24848
rect 24766 24792 24822 24848
rect 22006 19216 22062 19272
rect 21546 17856 21602 17912
rect 20810 14048 20866 14104
rect 20902 13812 20904 13832
rect 20904 13812 20956 13832
rect 20956 13812 20958 13832
rect 20902 13776 20958 13812
rect 20626 12960 20682 13016
rect 20166 6840 20222 6896
rect 19982 6568 20038 6624
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 20074 5616 20130 5672
rect 19522 5480 19578 5536
rect 19614 5228 19670 5264
rect 19614 5208 19616 5228
rect 19616 5208 19668 5228
rect 19668 5208 19670 5228
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20258 4820 20314 4856
rect 20258 4800 20260 4820
rect 20260 4800 20312 4820
rect 20312 4800 20314 4820
rect 21270 16652 21326 16688
rect 21270 16632 21272 16652
rect 21272 16632 21324 16652
rect 21324 16632 21326 16652
rect 21086 13096 21142 13152
rect 21086 12824 21142 12880
rect 21362 15000 21418 15056
rect 20994 10512 21050 10568
rect 22466 19624 22522 19680
rect 22742 19352 22798 19408
rect 23478 22616 23534 22672
rect 23202 18944 23258 19000
rect 22466 17720 22522 17776
rect 21730 15544 21786 15600
rect 22006 14184 22062 14240
rect 22282 17176 22338 17232
rect 23018 17584 23074 17640
rect 22374 15408 22430 15464
rect 23202 15680 23258 15736
rect 23202 15000 23258 15056
rect 21086 9968 21142 10024
rect 20902 9036 20958 9072
rect 20902 9016 20904 9036
rect 20904 9016 20956 9036
rect 20956 9016 20958 9036
rect 20718 8744 20774 8800
rect 20718 5752 20774 5808
rect 20902 4256 20958 4312
rect 21362 5480 21418 5536
rect 21270 2624 21326 2680
rect 20902 2508 20958 2544
rect 20902 2488 20904 2508
rect 20904 2488 20956 2508
rect 20956 2488 20958 2508
rect 20718 1944 20774 2000
rect 21822 7540 21878 7576
rect 21822 7520 21824 7540
rect 21824 7520 21876 7540
rect 21876 7520 21878 7540
rect 22006 11736 22062 11792
rect 22558 12688 22614 12744
rect 22374 9560 22430 9616
rect 22098 7928 22154 7984
rect 21730 3984 21786 4040
rect 22006 6568 22062 6624
rect 21914 6296 21970 6352
rect 22374 6976 22430 7032
rect 22834 13232 22890 13288
rect 23202 13912 23258 13968
rect 23938 21684 23994 21720
rect 23938 21664 23940 21684
rect 23940 21664 23992 21684
rect 23992 21664 23994 21684
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 25134 23704 25190 23760
rect 24674 23160 24730 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 23662 17856 23718 17912
rect 23478 16088 23534 16144
rect 23478 14864 23534 14920
rect 23478 13368 23534 13424
rect 23018 10412 23020 10432
rect 23020 10412 23072 10432
rect 23072 10412 23074 10432
rect 23018 10376 23074 10412
rect 23018 9444 23074 9480
rect 23018 9424 23020 9444
rect 23020 9424 23072 9444
rect 23072 9424 23074 9444
rect 22650 6704 22706 6760
rect 22190 4664 22246 4720
rect 22098 4120 22154 4176
rect 21730 3168 21786 3224
rect 22650 4528 22706 4584
rect 21638 2388 21640 2408
rect 21640 2388 21692 2408
rect 21692 2388 21694 2408
rect 21638 2352 21694 2388
rect 23478 9152 23534 9208
rect 23478 7928 23534 7984
rect 23110 7248 23166 7304
rect 23018 6296 23074 6352
rect 22834 4800 22890 4856
rect 23294 5616 23350 5672
rect 24122 21392 24178 21448
rect 24030 19896 24086 19952
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24582 21120 24638 21176
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24398 19916 24454 19952
rect 24398 19896 24400 19916
rect 24400 19896 24452 19916
rect 24452 19896 24454 19916
rect 24214 19760 24270 19816
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24122 19488 24178 19544
rect 25042 23296 25098 23352
rect 25042 22208 25098 22264
rect 24950 20984 25006 21040
rect 24674 19080 24730 19136
rect 24214 18808 24270 18864
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 17448 24822 17504
rect 24398 16904 24454 16960
rect 24490 16788 24546 16824
rect 24490 16768 24492 16788
rect 24492 16768 24544 16788
rect 24544 16768 24546 16788
rect 23846 16088 23902 16144
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24122 15272 24178 15328
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24122 15136 24178 15192
rect 25042 19352 25098 19408
rect 25410 22344 25466 22400
rect 27526 24520 27582 24576
rect 25686 23704 25742 23760
rect 25502 21528 25558 21584
rect 25226 20848 25282 20904
rect 25226 19252 25228 19272
rect 25228 19252 25280 19272
rect 25280 19252 25282 19272
rect 25226 19216 25282 19252
rect 25502 18944 25558 19000
rect 25502 18808 25558 18864
rect 23846 14592 23902 14648
rect 25042 14476 25098 14512
rect 25042 14456 25044 14476
rect 25044 14456 25096 14476
rect 25096 14456 25098 14476
rect 24030 14220 24032 14240
rect 24032 14220 24084 14240
rect 24084 14220 24086 14240
rect 24030 14184 24086 14220
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24030 12860 24032 12880
rect 24032 12860 24084 12880
rect 24084 12860 24086 12880
rect 24030 12824 24086 12860
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 23846 12280 23902 12336
rect 23570 7248 23626 7304
rect 23570 2624 23626 2680
rect 22742 1808 22798 1864
rect 23754 9424 23810 9480
rect 24214 12280 24270 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24122 10240 24178 10296
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24122 9696 24178 9752
rect 23846 8880 23902 8936
rect 23754 7792 23810 7848
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24214 8200 24270 8256
rect 24030 7384 24086 7440
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25318 16768 25374 16824
rect 25226 15988 25228 16008
rect 25228 15988 25280 16008
rect 25280 15988 25282 16008
rect 25226 15952 25282 15988
rect 25226 13912 25282 13968
rect 24766 8880 24822 8936
rect 25042 5616 25098 5672
rect 25042 4820 25098 4856
rect 25042 4800 25044 4820
rect 25044 4800 25096 4820
rect 25096 4800 25098 4820
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24766 4120 24822 4176
rect 24398 3984 24454 4040
rect 24674 3712 24730 3768
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23846 3032 23902 3088
rect 23754 2488 23810 2544
rect 23846 2352 23902 2408
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23938 1536 23994 1592
rect 25318 11212 25374 11248
rect 25318 11192 25320 11212
rect 25320 11192 25372 11212
rect 25372 11192 25374 11212
rect 25502 15408 25558 15464
rect 25410 9580 25466 9616
rect 25410 9560 25412 9580
rect 25412 9560 25464 9580
rect 25464 9560 25466 9580
rect 25318 6976 25374 7032
rect 25502 5072 25558 5128
rect 25502 4528 25558 4584
rect 26054 4256 26110 4312
rect 25594 3576 25650 3632
rect 23570 312 23626 368
<< metal3 >>
rect 24577 27706 24643 27709
rect 27520 27706 28000 27736
rect 24577 27704 28000 27706
rect 24577 27648 24582 27704
rect 24638 27648 28000 27704
rect 24577 27646 28000 27648
rect 24577 27643 24643 27646
rect 27520 27616 28000 27646
rect 24761 27162 24827 27165
rect 27520 27162 28000 27192
rect 24761 27160 28000 27162
rect 24761 27104 24766 27160
rect 24822 27104 28000 27160
rect 24761 27102 28000 27104
rect 24761 27099 24827 27102
rect 27520 27072 28000 27102
rect 23381 26618 23447 26621
rect 27520 26618 28000 26648
rect 23381 26616 28000 26618
rect 23381 26560 23386 26616
rect 23442 26560 28000 26616
rect 23381 26558 28000 26560
rect 23381 26555 23447 26558
rect 27520 26528 28000 26558
rect 23289 26074 23355 26077
rect 27520 26074 28000 26104
rect 23289 26072 28000 26074
rect 23289 26016 23294 26072
rect 23350 26016 28000 26072
rect 23289 26014 28000 26016
rect 23289 26011 23355 26014
rect 27520 25984 28000 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 23657 25394 23723 25397
rect 27520 25394 28000 25424
rect 23657 25392 28000 25394
rect 23657 25336 23662 25392
rect 23718 25336 28000 25392
rect 23657 25334 28000 25336
rect 23657 25331 23723 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 12709 24850 12775 24853
rect 14549 24850 14615 24853
rect 12709 24848 14615 24850
rect 12709 24792 12714 24848
rect 12770 24792 14554 24848
rect 14610 24792 14615 24848
rect 12709 24790 14615 24792
rect 12709 24787 12775 24790
rect 14549 24787 14615 24790
rect 15469 24850 15535 24853
rect 24577 24850 24643 24853
rect 15469 24848 24643 24850
rect 15469 24792 15474 24848
rect 15530 24792 24582 24848
rect 24638 24792 24643 24848
rect 15469 24790 24643 24792
rect 15469 24787 15535 24790
rect 24577 24787 24643 24790
rect 24761 24850 24827 24853
rect 27520 24850 28000 24880
rect 24761 24848 28000 24850
rect 24761 24792 24766 24848
rect 24822 24792 28000 24848
rect 24761 24790 28000 24792
rect 24761 24787 24827 24790
rect 27520 24760 28000 24790
rect 9121 24714 9187 24717
rect 14917 24714 14983 24717
rect 15929 24714 15995 24717
rect 9121 24712 14842 24714
rect 9121 24656 9126 24712
rect 9182 24656 14842 24712
rect 9121 24654 14842 24656
rect 9121 24651 9187 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 14782 24442 14842 24654
rect 14917 24712 15995 24714
rect 14917 24656 14922 24712
rect 14978 24656 15934 24712
rect 15990 24656 15995 24712
rect 14917 24654 15995 24656
rect 14917 24651 14983 24654
rect 15929 24651 15995 24654
rect 21081 24578 21147 24581
rect 27521 24578 27587 24581
rect 21081 24576 27587 24578
rect 21081 24520 21086 24576
rect 21142 24520 27526 24576
rect 27582 24520 27587 24576
rect 21081 24518 27587 24520
rect 21081 24515 21147 24518
rect 27521 24515 27587 24518
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 15837 24442 15903 24445
rect 14782 24440 15903 24442
rect 14782 24384 15842 24440
rect 15898 24384 15903 24440
rect 14782 24382 15903 24384
rect 15837 24379 15903 24382
rect 21541 24442 21607 24445
rect 23473 24442 23539 24445
rect 21541 24440 23539 24442
rect 21541 24384 21546 24440
rect 21602 24384 23478 24440
rect 23534 24384 23539 24440
rect 21541 24382 23539 24384
rect 21541 24379 21607 24382
rect 23473 24379 23539 24382
rect 7741 24306 7807 24309
rect 10685 24306 10751 24309
rect 7741 24304 10751 24306
rect 7741 24248 7746 24304
rect 7802 24248 10690 24304
rect 10746 24248 10751 24304
rect 7741 24246 10751 24248
rect 7741 24243 7807 24246
rect 10685 24243 10751 24246
rect 11881 24306 11947 24309
rect 20805 24306 20871 24309
rect 11881 24304 20871 24306
rect 11881 24248 11886 24304
rect 11942 24248 20810 24304
rect 20866 24248 20871 24304
rect 11881 24246 20871 24248
rect 11881 24243 11947 24246
rect 20805 24243 20871 24246
rect 22277 24306 22343 24309
rect 27520 24306 28000 24336
rect 22277 24304 28000 24306
rect 22277 24248 22282 24304
rect 22338 24248 28000 24304
rect 22277 24246 28000 24248
rect 22277 24243 22343 24246
rect 27520 24216 28000 24246
rect 10777 24170 10843 24173
rect 13261 24170 13327 24173
rect 18873 24170 18939 24173
rect 10777 24168 13327 24170
rect 10777 24112 10782 24168
rect 10838 24112 13266 24168
rect 13322 24112 13327 24168
rect 10777 24110 13327 24112
rect 10777 24107 10843 24110
rect 13261 24107 13327 24110
rect 14782 24168 18939 24170
rect 14782 24112 18878 24168
rect 18934 24112 18939 24168
rect 14782 24110 18939 24112
rect 9765 24034 9831 24037
rect 14782 24034 14842 24110
rect 18873 24107 18939 24110
rect 9765 24032 14842 24034
rect 9765 23976 9770 24032
rect 9826 23976 14842 24032
rect 9765 23974 14842 23976
rect 9765 23971 9831 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 12617 23762 12683 23765
rect 25129 23762 25195 23765
rect 12617 23760 25195 23762
rect 12617 23704 12622 23760
rect 12678 23704 25134 23760
rect 25190 23704 25195 23760
rect 12617 23702 25195 23704
rect 12617 23699 12683 23702
rect 25129 23699 25195 23702
rect 25681 23762 25747 23765
rect 27520 23762 28000 23792
rect 25681 23760 28000 23762
rect 25681 23704 25686 23760
rect 25742 23704 28000 23760
rect 25681 23702 28000 23704
rect 25681 23699 25747 23702
rect 27520 23672 28000 23702
rect 7097 23626 7163 23629
rect 9305 23626 9371 23629
rect 7097 23624 9371 23626
rect 7097 23568 7102 23624
rect 7158 23568 9310 23624
rect 9366 23568 9371 23624
rect 7097 23566 9371 23568
rect 7097 23563 7163 23566
rect 9305 23563 9371 23566
rect 6361 23490 6427 23493
rect 7741 23490 7807 23493
rect 6361 23488 7807 23490
rect 6361 23432 6366 23488
rect 6422 23432 7746 23488
rect 7802 23432 7807 23488
rect 6361 23430 7807 23432
rect 6361 23427 6427 23430
rect 7741 23427 7807 23430
rect 15653 23490 15719 23493
rect 16941 23490 17007 23493
rect 15653 23488 17007 23490
rect 15653 23432 15658 23488
rect 15714 23432 16946 23488
rect 17002 23432 17007 23488
rect 15653 23430 17007 23432
rect 15653 23427 15719 23430
rect 16941 23427 17007 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 14549 23354 14615 23357
rect 16389 23354 16455 23357
rect 14549 23352 16455 23354
rect 14549 23296 14554 23352
rect 14610 23296 16394 23352
rect 16450 23296 16455 23352
rect 14549 23294 16455 23296
rect 14549 23291 14615 23294
rect 16389 23291 16455 23294
rect 21173 23354 21239 23357
rect 25037 23354 25103 23357
rect 21173 23352 25103 23354
rect 21173 23296 21178 23352
rect 21234 23296 25042 23352
rect 25098 23296 25103 23352
rect 21173 23294 25103 23296
rect 21173 23291 21239 23294
rect 25037 23291 25103 23294
rect 11237 23218 11303 23221
rect 17769 23218 17835 23221
rect 11237 23216 17835 23218
rect 11237 23160 11242 23216
rect 11298 23160 17774 23216
rect 17830 23160 17835 23216
rect 11237 23158 17835 23160
rect 11237 23155 11303 23158
rect 17769 23155 17835 23158
rect 24669 23218 24735 23221
rect 27520 23218 28000 23248
rect 24669 23216 28000 23218
rect 24669 23160 24674 23216
rect 24730 23160 28000 23216
rect 24669 23158 28000 23160
rect 24669 23155 24735 23158
rect 27520 23128 28000 23158
rect 933 23082 999 23085
rect 14089 23082 14155 23085
rect 933 23080 14155 23082
rect 933 23024 938 23080
rect 994 23024 14094 23080
rect 14150 23024 14155 23080
rect 933 23022 14155 23024
rect 933 23019 999 23022
rect 14089 23019 14155 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 4981 22674 5047 22677
rect 12341 22674 12407 22677
rect 4981 22672 12407 22674
rect 4981 22616 4986 22672
rect 5042 22616 12346 22672
rect 12402 22616 12407 22672
rect 4981 22614 12407 22616
rect 4981 22611 5047 22614
rect 12341 22611 12407 22614
rect 20805 22674 20871 22677
rect 23473 22674 23539 22677
rect 20805 22672 23539 22674
rect 20805 22616 20810 22672
rect 20866 22616 23478 22672
rect 23534 22616 23539 22672
rect 20805 22614 23539 22616
rect 20805 22611 20871 22614
rect 23473 22611 23539 22614
rect 2957 22538 3023 22541
rect 13445 22538 13511 22541
rect 2957 22536 13511 22538
rect 2957 22480 2962 22536
rect 3018 22480 13450 22536
rect 13506 22480 13511 22536
rect 2957 22478 13511 22480
rect 2957 22475 3023 22478
rect 13445 22475 13511 22478
rect 13629 22538 13695 22541
rect 15285 22538 15351 22541
rect 21265 22538 21331 22541
rect 13629 22536 15351 22538
rect 13629 22480 13634 22536
rect 13690 22480 15290 22536
rect 15346 22480 15351 22536
rect 13629 22478 15351 22480
rect 13629 22475 13695 22478
rect 15285 22475 15351 22478
rect 19382 22536 21331 22538
rect 19382 22480 21270 22536
rect 21326 22480 21331 22536
rect 19382 22478 21331 22480
rect 11881 22402 11947 22405
rect 18505 22402 18571 22405
rect 19382 22402 19442 22478
rect 21265 22475 21331 22478
rect 21449 22538 21515 22541
rect 27520 22538 28000 22568
rect 21449 22536 28000 22538
rect 21449 22480 21454 22536
rect 21510 22480 28000 22536
rect 21449 22478 28000 22480
rect 21449 22475 21515 22478
rect 27520 22448 28000 22478
rect 11881 22400 19442 22402
rect 11881 22344 11886 22400
rect 11942 22344 18510 22400
rect 18566 22344 19442 22400
rect 11881 22342 19442 22344
rect 22737 22402 22803 22405
rect 25405 22402 25471 22405
rect 22737 22400 25471 22402
rect 22737 22344 22742 22400
rect 22798 22344 25410 22400
rect 25466 22344 25471 22400
rect 22737 22342 25471 22344
rect 11881 22339 11947 22342
rect 18505 22339 18571 22342
rect 22737 22339 22803 22342
rect 25405 22339 25471 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 10869 22266 10935 22269
rect 15837 22266 15903 22269
rect 18505 22266 18571 22269
rect 10869 22264 14842 22266
rect 10869 22208 10874 22264
rect 10930 22208 14842 22264
rect 10869 22206 14842 22208
rect 10869 22203 10935 22206
rect 14782 22130 14842 22206
rect 15837 22264 18571 22266
rect 15837 22208 15842 22264
rect 15898 22208 18510 22264
rect 18566 22208 18571 22264
rect 15837 22206 18571 22208
rect 15837 22203 15903 22206
rect 18505 22203 18571 22206
rect 20621 22266 20687 22269
rect 22277 22266 22343 22269
rect 25037 22266 25103 22269
rect 20621 22264 22343 22266
rect 20621 22208 20626 22264
rect 20682 22208 22282 22264
rect 22338 22208 22343 22264
rect 20621 22206 22343 22208
rect 20621 22203 20687 22206
rect 22277 22203 22343 22206
rect 22510 22264 25103 22266
rect 22510 22208 25042 22264
rect 25098 22208 25103 22264
rect 22510 22206 25103 22208
rect 17033 22130 17099 22133
rect 22510 22130 22570 22206
rect 25037 22203 25103 22206
rect 14782 22128 17099 22130
rect 14782 22072 17038 22128
rect 17094 22072 17099 22128
rect 14782 22070 17099 22072
rect 17033 22067 17099 22070
rect 17726 22070 22570 22130
rect 22645 22130 22711 22133
rect 22645 22128 24410 22130
rect 22645 22072 22650 22128
rect 22706 22072 24410 22128
rect 22645 22070 24410 22072
rect 15561 21994 15627 21997
rect 17726 21994 17786 22070
rect 22645 22067 22711 22070
rect 15561 21992 17786 21994
rect 15561 21936 15566 21992
rect 15622 21936 17786 21992
rect 15561 21934 17786 21936
rect 24350 21994 24410 22070
rect 27520 21994 28000 22024
rect 24350 21934 28000 21994
rect 15561 21931 15627 21934
rect 27520 21904 28000 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 23933 21722 23999 21725
rect 15334 21720 23999 21722
rect 15334 21664 23938 21720
rect 23994 21664 23999 21720
rect 15334 21662 23999 21664
rect 12709 21586 12775 21589
rect 15334 21586 15394 21662
rect 23933 21659 23999 21662
rect 12709 21584 15394 21586
rect 12709 21528 12714 21584
rect 12770 21528 15394 21584
rect 12709 21526 15394 21528
rect 19977 21586 20043 21589
rect 25497 21586 25563 21589
rect 19977 21584 25563 21586
rect 19977 21528 19982 21584
rect 20038 21528 25502 21584
rect 25558 21528 25563 21584
rect 19977 21526 25563 21528
rect 12709 21523 12775 21526
rect 19977 21523 20043 21526
rect 25497 21523 25563 21526
rect 24117 21450 24183 21453
rect 27520 21450 28000 21480
rect 24117 21448 28000 21450
rect 24117 21392 24122 21448
rect 24178 21392 28000 21448
rect 24117 21390 28000 21392
rect 24117 21387 24183 21390
rect 27520 21360 28000 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 12341 21178 12407 21181
rect 14641 21178 14707 21181
rect 12341 21176 14707 21178
rect 12341 21120 12346 21176
rect 12402 21120 14646 21176
rect 14702 21120 14707 21176
rect 12341 21118 14707 21120
rect 12341 21115 12407 21118
rect 14641 21115 14707 21118
rect 21817 21178 21883 21181
rect 24577 21178 24643 21181
rect 21817 21176 24643 21178
rect 21817 21120 21822 21176
rect 21878 21120 24582 21176
rect 24638 21120 24643 21176
rect 21817 21118 24643 21120
rect 21817 21115 21883 21118
rect 24577 21115 24643 21118
rect 0 21042 480 21072
rect 4061 21042 4127 21045
rect 0 21040 4127 21042
rect 0 20984 4066 21040
rect 4122 20984 4127 21040
rect 0 20982 4127 20984
rect 0 20952 480 20982
rect 4061 20979 4127 20982
rect 9213 21042 9279 21045
rect 12433 21042 12499 21045
rect 9213 21040 12499 21042
rect 9213 20984 9218 21040
rect 9274 20984 12438 21040
rect 12494 20984 12499 21040
rect 9213 20982 12499 20984
rect 9213 20979 9279 20982
rect 12433 20979 12499 20982
rect 20345 21042 20411 21045
rect 24945 21042 25011 21045
rect 20345 21040 25011 21042
rect 20345 20984 20350 21040
rect 20406 20984 24950 21040
rect 25006 20984 25011 21040
rect 20345 20982 25011 20984
rect 20345 20979 20411 20982
rect 24945 20979 25011 20982
rect 13997 20906 14063 20909
rect 20897 20906 20963 20909
rect 21633 20906 21699 20909
rect 13997 20904 21699 20906
rect 13997 20848 14002 20904
rect 14058 20848 20902 20904
rect 20958 20848 21638 20904
rect 21694 20848 21699 20904
rect 13997 20846 21699 20848
rect 13997 20843 14063 20846
rect 20897 20843 20963 20846
rect 21633 20843 21699 20846
rect 25221 20906 25287 20909
rect 27520 20906 28000 20936
rect 25221 20904 28000 20906
rect 25221 20848 25226 20904
rect 25282 20848 28000 20904
rect 25221 20846 28000 20848
rect 25221 20843 25287 20846
rect 27520 20816 28000 20846
rect 18505 20770 18571 20773
rect 20253 20770 20319 20773
rect 18505 20768 20319 20770
rect 18505 20712 18510 20768
rect 18566 20712 20258 20768
rect 20314 20712 20319 20768
rect 18505 20710 20319 20712
rect 18505 20707 18571 20710
rect 20253 20707 20319 20710
rect 21081 20770 21147 20773
rect 21081 20768 24042 20770
rect 21081 20712 21086 20768
rect 21142 20712 24042 20768
rect 21081 20710 24042 20712
rect 21081 20707 21147 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 11237 20498 11303 20501
rect 20989 20498 21055 20501
rect 11237 20496 21055 20498
rect 11237 20440 11242 20496
rect 11298 20440 20994 20496
rect 21050 20440 21055 20496
rect 11237 20438 21055 20440
rect 11237 20435 11303 20438
rect 20989 20435 21055 20438
rect 7833 20362 7899 20365
rect 16205 20362 16271 20365
rect 7833 20360 16271 20362
rect 7833 20304 7838 20360
rect 7894 20304 16210 20360
rect 16266 20304 16271 20360
rect 7833 20302 16271 20304
rect 7833 20299 7899 20302
rect 16205 20299 16271 20302
rect 17033 20362 17099 20365
rect 20805 20362 20871 20365
rect 17033 20360 20871 20362
rect 17033 20304 17038 20360
rect 17094 20304 20810 20360
rect 20866 20304 20871 20360
rect 17033 20302 20871 20304
rect 23982 20362 24042 20710
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 27520 20362 28000 20392
rect 23982 20302 28000 20362
rect 17033 20299 17099 20302
rect 20805 20299 20871 20302
rect 27520 20272 28000 20302
rect 16389 20226 16455 20229
rect 18137 20226 18203 20229
rect 18781 20226 18847 20229
rect 16389 20224 18847 20226
rect 16389 20168 16394 20224
rect 16450 20168 18142 20224
rect 18198 20168 18786 20224
rect 18842 20168 18847 20224
rect 16389 20166 18847 20168
rect 16389 20163 16455 20166
rect 18137 20163 18203 20166
rect 18781 20163 18847 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 5993 20090 6059 20093
rect 7833 20090 7899 20093
rect 5993 20088 7899 20090
rect 5993 20032 5998 20088
rect 6054 20032 7838 20088
rect 7894 20032 7899 20088
rect 5993 20030 7899 20032
rect 5993 20027 6059 20030
rect 7833 20027 7899 20030
rect 13353 20090 13419 20093
rect 16573 20090 16639 20093
rect 13353 20088 16639 20090
rect 13353 20032 13358 20088
rect 13414 20032 16578 20088
rect 16634 20032 16639 20088
rect 13353 20030 16639 20032
rect 13353 20027 13419 20030
rect 16573 20027 16639 20030
rect 3693 19954 3759 19957
rect 14733 19954 14799 19957
rect 3693 19952 14799 19954
rect 3693 19896 3698 19952
rect 3754 19896 14738 19952
rect 14794 19896 14799 19952
rect 3693 19894 14799 19896
rect 3693 19891 3759 19894
rect 14733 19891 14799 19894
rect 17217 19954 17283 19957
rect 18413 19954 18479 19957
rect 24025 19954 24091 19957
rect 24393 19954 24459 19957
rect 17217 19952 24459 19954
rect 17217 19896 17222 19952
rect 17278 19896 18418 19952
rect 18474 19896 24030 19952
rect 24086 19896 24398 19952
rect 24454 19896 24459 19952
rect 17217 19894 24459 19896
rect 17217 19891 17283 19894
rect 18413 19891 18479 19894
rect 24025 19891 24091 19894
rect 24393 19891 24459 19894
rect 9305 19818 9371 19821
rect 15837 19818 15903 19821
rect 9305 19816 15903 19818
rect 9305 19760 9310 19816
rect 9366 19760 15842 19816
rect 15898 19760 15903 19816
rect 9305 19758 15903 19760
rect 9305 19755 9371 19758
rect 15837 19755 15903 19758
rect 24209 19818 24275 19821
rect 24209 19816 24824 19818
rect 24209 19760 24214 19816
rect 24270 19760 24824 19816
rect 24209 19758 24824 19760
rect 24209 19755 24275 19758
rect 20897 19682 20963 19685
rect 22461 19682 22527 19685
rect 20897 19680 22527 19682
rect 20897 19624 20902 19680
rect 20958 19624 22466 19680
rect 22522 19624 22527 19680
rect 20897 19622 22527 19624
rect 24764 19682 24824 19758
rect 27520 19682 28000 19712
rect 24764 19622 28000 19682
rect 20897 19619 20963 19622
rect 22461 19619 22527 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19622
rect 24277 19551 24597 19552
rect 20989 19546 21055 19549
rect 24117 19546 24183 19549
rect 20989 19544 24183 19546
rect 20989 19488 20994 19544
rect 21050 19488 24122 19544
rect 24178 19488 24183 19544
rect 20989 19486 24183 19488
rect 20989 19483 21055 19486
rect 24117 19483 24183 19486
rect 14457 19410 14523 19413
rect 15745 19410 15811 19413
rect 14457 19408 15811 19410
rect 14457 19352 14462 19408
rect 14518 19352 15750 19408
rect 15806 19352 15811 19408
rect 14457 19350 15811 19352
rect 14457 19347 14523 19350
rect 15745 19347 15811 19350
rect 18321 19410 18387 19413
rect 21081 19410 21147 19413
rect 18321 19408 21147 19410
rect 18321 19352 18326 19408
rect 18382 19352 21086 19408
rect 21142 19352 21147 19408
rect 18321 19350 21147 19352
rect 18321 19347 18387 19350
rect 21081 19347 21147 19350
rect 22737 19410 22803 19413
rect 25037 19410 25103 19413
rect 22737 19408 25103 19410
rect 22737 19352 22742 19408
rect 22798 19352 25042 19408
rect 25098 19352 25103 19408
rect 22737 19350 25103 19352
rect 22737 19347 22803 19350
rect 25037 19347 25103 19350
rect 1577 19274 1643 19277
rect 10593 19274 10659 19277
rect 1577 19272 10659 19274
rect 1577 19216 1582 19272
rect 1638 19216 10598 19272
rect 10654 19216 10659 19272
rect 1577 19214 10659 19216
rect 1577 19211 1643 19214
rect 10593 19211 10659 19214
rect 18413 19274 18479 19277
rect 21357 19274 21423 19277
rect 18413 19272 21423 19274
rect 18413 19216 18418 19272
rect 18474 19216 21362 19272
rect 21418 19216 21423 19272
rect 18413 19214 21423 19216
rect 18413 19211 18479 19214
rect 21357 19211 21423 19214
rect 22001 19274 22067 19277
rect 25221 19274 25287 19277
rect 22001 19272 25287 19274
rect 22001 19216 22006 19272
rect 22062 19216 25226 19272
rect 25282 19216 25287 19272
rect 22001 19214 25287 19216
rect 22001 19211 22067 19214
rect 25221 19211 25287 19214
rect 9305 19138 9371 19141
rect 9581 19138 9647 19141
rect 9305 19136 9647 19138
rect 9305 19080 9310 19136
rect 9366 19080 9586 19136
rect 9642 19080 9647 19136
rect 9305 19078 9647 19080
rect 9305 19075 9371 19078
rect 9581 19075 9647 19078
rect 24669 19138 24735 19141
rect 27520 19138 28000 19168
rect 24669 19136 28000 19138
rect 24669 19080 24674 19136
rect 24730 19080 28000 19136
rect 24669 19078 28000 19080
rect 24669 19075 24735 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 4337 19002 4403 19005
rect 10133 19002 10199 19005
rect 4337 19000 10199 19002
rect 4337 18944 4342 19000
rect 4398 18944 10138 19000
rect 10194 18944 10199 19000
rect 4337 18942 10199 18944
rect 4337 18939 4403 18942
rect 10133 18939 10199 18942
rect 23197 19002 23263 19005
rect 25497 19002 25563 19005
rect 23197 19000 25563 19002
rect 23197 18944 23202 19000
rect 23258 18944 25502 19000
rect 25558 18944 25563 19000
rect 23197 18942 25563 18944
rect 23197 18939 23263 18942
rect 25497 18939 25563 18942
rect 14825 18866 14891 18869
rect 17309 18866 17375 18869
rect 18045 18866 18111 18869
rect 14825 18864 18111 18866
rect 14825 18808 14830 18864
rect 14886 18808 17314 18864
rect 17370 18808 18050 18864
rect 18106 18808 18111 18864
rect 14825 18806 18111 18808
rect 14825 18803 14891 18806
rect 17309 18803 17375 18806
rect 18045 18803 18111 18806
rect 18873 18866 18939 18869
rect 21173 18866 21239 18869
rect 18873 18864 21239 18866
rect 18873 18808 18878 18864
rect 18934 18808 21178 18864
rect 21234 18808 21239 18864
rect 18873 18806 21239 18808
rect 18873 18803 18939 18806
rect 21173 18803 21239 18806
rect 24209 18866 24275 18869
rect 25497 18866 25563 18869
rect 24209 18864 25563 18866
rect 24209 18808 24214 18864
rect 24270 18808 25502 18864
rect 25558 18808 25563 18864
rect 24209 18806 25563 18808
rect 24209 18803 24275 18806
rect 25497 18803 25563 18806
rect 21081 18730 21147 18733
rect 21081 18728 24962 18730
rect 21081 18672 21086 18728
rect 21142 18672 24962 18728
rect 21081 18670 24962 18672
rect 21081 18667 21147 18670
rect 12249 18594 12315 18597
rect 14273 18594 14339 18597
rect 12249 18592 14339 18594
rect 12249 18536 12254 18592
rect 12310 18536 14278 18592
rect 14334 18536 14339 18592
rect 12249 18534 14339 18536
rect 24902 18594 24962 18670
rect 27520 18594 28000 18624
rect 24902 18534 28000 18594
rect 12249 18531 12315 18534
rect 14273 18531 14339 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 27520 18504 28000 18534
rect 24277 18463 24597 18464
rect 10961 18322 11027 18325
rect 20345 18322 20411 18325
rect 10961 18320 20411 18322
rect 10961 18264 10966 18320
rect 11022 18264 20350 18320
rect 20406 18264 20411 18320
rect 10961 18262 20411 18264
rect 10961 18259 11027 18262
rect 20345 18259 20411 18262
rect 11605 18186 11671 18189
rect 12893 18186 12959 18189
rect 11605 18184 12959 18186
rect 11605 18128 11610 18184
rect 11666 18128 12898 18184
rect 12954 18128 12959 18184
rect 11605 18126 12959 18128
rect 11605 18123 11671 18126
rect 12893 18123 12959 18126
rect 13629 18186 13695 18189
rect 16389 18186 16455 18189
rect 13629 18184 16455 18186
rect 13629 18128 13634 18184
rect 13690 18128 16394 18184
rect 16450 18128 16455 18184
rect 13629 18126 16455 18128
rect 13629 18123 13695 18126
rect 16389 18123 16455 18126
rect 17166 17988 17172 18052
rect 17236 18050 17242 18052
rect 17401 18050 17467 18053
rect 17236 18048 17467 18050
rect 17236 17992 17406 18048
rect 17462 17992 17467 18048
rect 17236 17990 17467 17992
rect 17236 17988 17242 17990
rect 17401 17987 17467 17990
rect 18597 18050 18663 18053
rect 19333 18050 19399 18053
rect 18597 18048 19399 18050
rect 18597 17992 18602 18048
rect 18658 17992 19338 18048
rect 19394 17992 19399 18048
rect 18597 17990 19399 17992
rect 18597 17987 18663 17990
rect 19333 17987 19399 17990
rect 21265 18050 21331 18053
rect 27520 18050 28000 18080
rect 21265 18048 28000 18050
rect 21265 17992 21270 18048
rect 21326 17992 28000 18048
rect 21265 17990 28000 17992
rect 21265 17987 21331 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 21541 17914 21607 17917
rect 23657 17914 23723 17917
rect 21541 17912 23723 17914
rect 21541 17856 21546 17912
rect 21602 17856 23662 17912
rect 23718 17856 23723 17912
rect 21541 17854 23723 17856
rect 21541 17851 21607 17854
rect 23657 17851 23723 17854
rect 14089 17778 14155 17781
rect 22461 17778 22527 17781
rect 14089 17776 22527 17778
rect 14089 17720 14094 17776
rect 14150 17720 22466 17776
rect 22522 17720 22527 17776
rect 14089 17718 22527 17720
rect 14089 17715 14155 17718
rect 22461 17715 22527 17718
rect 13905 17642 13971 17645
rect 14733 17642 14799 17645
rect 19977 17642 20043 17645
rect 23013 17642 23079 17645
rect 13905 17640 23079 17642
rect 13905 17584 13910 17640
rect 13966 17584 14738 17640
rect 14794 17584 19982 17640
rect 20038 17584 23018 17640
rect 23074 17584 23079 17640
rect 13905 17582 23079 17584
rect 13905 17579 13971 17582
rect 14733 17579 14799 17582
rect 19977 17579 20043 17582
rect 23013 17579 23079 17582
rect 24761 17506 24827 17509
rect 27520 17506 28000 17536
rect 24761 17504 28000 17506
rect 24761 17448 24766 17504
rect 24822 17448 28000 17504
rect 24761 17446 28000 17448
rect 24761 17443 24827 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 18689 17234 18755 17237
rect 22277 17234 22343 17237
rect 18689 17232 22343 17234
rect 18689 17176 18694 17232
rect 18750 17176 22282 17232
rect 22338 17176 22343 17232
rect 18689 17174 22343 17176
rect 18689 17171 18755 17174
rect 22277 17171 22343 17174
rect 9489 17098 9555 17101
rect 12893 17098 12959 17101
rect 9489 17096 12959 17098
rect 9489 17040 9494 17096
rect 9550 17040 12898 17096
rect 12954 17040 12959 17096
rect 9489 17038 12959 17040
rect 9489 17035 9555 17038
rect 12893 17035 12959 17038
rect 13169 17098 13235 17101
rect 15377 17098 15443 17101
rect 13169 17096 15443 17098
rect 13169 17040 13174 17096
rect 13230 17040 15382 17096
rect 15438 17040 15443 17096
rect 13169 17038 15443 17040
rect 13169 17035 13235 17038
rect 15377 17035 15443 17038
rect 12985 16962 13051 16965
rect 15285 16962 15351 16965
rect 12985 16960 15351 16962
rect 12985 16904 12990 16960
rect 13046 16904 15290 16960
rect 15346 16904 15351 16960
rect 12985 16902 15351 16904
rect 12985 16899 13051 16902
rect 15285 16899 15351 16902
rect 20621 16962 20687 16965
rect 24393 16962 24459 16965
rect 20621 16960 24459 16962
rect 20621 16904 20626 16960
rect 20682 16904 24398 16960
rect 24454 16904 24459 16960
rect 20621 16902 24459 16904
rect 20621 16899 20687 16902
rect 24393 16899 24459 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 12617 16826 12683 16829
rect 13629 16826 13695 16829
rect 20529 16826 20595 16829
rect 24485 16826 24551 16829
rect 12617 16824 13554 16826
rect 12617 16768 12622 16824
rect 12678 16768 13554 16824
rect 12617 16766 13554 16768
rect 12617 16763 12683 16766
rect 11697 16690 11763 16693
rect 13169 16690 13235 16693
rect 11697 16688 13235 16690
rect 11697 16632 11702 16688
rect 11758 16632 13174 16688
rect 13230 16632 13235 16688
rect 11697 16630 13235 16632
rect 13494 16690 13554 16766
rect 13629 16824 18154 16826
rect 13629 16768 13634 16824
rect 13690 16768 18154 16824
rect 13629 16766 18154 16768
rect 13629 16763 13695 16766
rect 15745 16690 15811 16693
rect 17953 16690 18019 16693
rect 13494 16630 15578 16690
rect 11697 16627 11763 16630
rect 13169 16627 13235 16630
rect 15518 16554 15578 16630
rect 15745 16688 18019 16690
rect 15745 16632 15750 16688
rect 15806 16632 17958 16688
rect 18014 16632 18019 16688
rect 15745 16630 18019 16632
rect 18094 16690 18154 16766
rect 20529 16824 24551 16826
rect 20529 16768 20534 16824
rect 20590 16768 24490 16824
rect 24546 16768 24551 16824
rect 20529 16766 24551 16768
rect 20529 16763 20595 16766
rect 24485 16763 24551 16766
rect 25313 16826 25379 16829
rect 27520 16826 28000 16856
rect 25313 16824 28000 16826
rect 25313 16768 25318 16824
rect 25374 16768 28000 16824
rect 25313 16766 28000 16768
rect 25313 16763 25379 16766
rect 27520 16736 28000 16766
rect 21265 16690 21331 16693
rect 18094 16688 21331 16690
rect 18094 16632 21270 16688
rect 21326 16632 21331 16688
rect 18094 16630 21331 16632
rect 15745 16627 15811 16630
rect 17953 16627 18019 16630
rect 21265 16627 21331 16630
rect 15745 16554 15811 16557
rect 15518 16552 15811 16554
rect 15518 16496 15750 16552
rect 15806 16496 15811 16552
rect 15518 16494 15811 16496
rect 15745 16491 15811 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 27520 16282 28000 16312
rect 24764 16222 28000 16282
rect 14273 16146 14339 16149
rect 23473 16146 23539 16149
rect 14273 16144 23539 16146
rect 14273 16088 14278 16144
rect 14334 16088 23478 16144
rect 23534 16088 23539 16144
rect 14273 16086 23539 16088
rect 14273 16083 14339 16086
rect 23473 16083 23539 16086
rect 23841 16146 23907 16149
rect 24764 16146 24824 16222
rect 27520 16192 28000 16222
rect 23841 16144 24824 16146
rect 23841 16088 23846 16144
rect 23902 16088 24824 16144
rect 23841 16086 24824 16088
rect 23841 16083 23907 16086
rect 10041 16010 10107 16013
rect 18781 16010 18847 16013
rect 10041 16008 18847 16010
rect 10041 15952 10046 16008
rect 10102 15952 18786 16008
rect 18842 15952 18847 16008
rect 10041 15950 18847 15952
rect 10041 15947 10107 15950
rect 18781 15947 18847 15950
rect 20069 16010 20135 16013
rect 25221 16010 25287 16013
rect 20069 16008 25287 16010
rect 20069 15952 20074 16008
rect 20130 15952 25226 16008
rect 25282 15952 25287 16008
rect 20069 15950 25287 15952
rect 20069 15947 20135 15950
rect 25221 15947 25287 15950
rect 10869 15874 10935 15877
rect 18505 15874 18571 15877
rect 10869 15872 18571 15874
rect 10869 15816 10874 15872
rect 10930 15816 18510 15872
rect 18566 15816 18571 15872
rect 10869 15814 18571 15816
rect 10869 15811 10935 15814
rect 18505 15811 18571 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 14181 15738 14247 15741
rect 19425 15738 19491 15741
rect 14181 15736 19491 15738
rect 14181 15680 14186 15736
rect 14242 15680 19430 15736
rect 19486 15680 19491 15736
rect 14181 15678 19491 15680
rect 14181 15675 14247 15678
rect 19425 15675 19491 15678
rect 23197 15738 23263 15741
rect 27520 15738 28000 15768
rect 23197 15736 28000 15738
rect 23197 15680 23202 15736
rect 23258 15680 28000 15736
rect 23197 15678 28000 15680
rect 23197 15675 23263 15678
rect 27520 15648 28000 15678
rect 13445 15602 13511 15605
rect 18413 15602 18479 15605
rect 13445 15600 18479 15602
rect 13445 15544 13450 15600
rect 13506 15544 18418 15600
rect 18474 15544 18479 15600
rect 13445 15542 18479 15544
rect 13445 15539 13511 15542
rect 18413 15539 18479 15542
rect 19241 15602 19307 15605
rect 21725 15602 21791 15605
rect 19241 15600 21791 15602
rect 19241 15544 19246 15600
rect 19302 15544 21730 15600
rect 21786 15544 21791 15600
rect 19241 15542 21791 15544
rect 19241 15539 19307 15542
rect 21725 15539 21791 15542
rect 381 15466 447 15469
rect 10777 15466 10843 15469
rect 11237 15466 11303 15469
rect 381 15464 11303 15466
rect 381 15408 386 15464
rect 442 15408 10782 15464
rect 10838 15408 11242 15464
rect 11298 15408 11303 15464
rect 381 15406 11303 15408
rect 381 15403 447 15406
rect 10777 15403 10843 15406
rect 11237 15403 11303 15406
rect 13169 15466 13235 15469
rect 15469 15466 15535 15469
rect 13169 15464 15535 15466
rect 13169 15408 13174 15464
rect 13230 15408 15474 15464
rect 15530 15408 15535 15464
rect 13169 15406 15535 15408
rect 13169 15403 13235 15406
rect 15469 15403 15535 15406
rect 22369 15466 22435 15469
rect 25497 15466 25563 15469
rect 22369 15464 25563 15466
rect 22369 15408 22374 15464
rect 22430 15408 25502 15464
rect 25558 15408 25563 15464
rect 22369 15406 25563 15408
rect 22369 15403 22435 15406
rect 25497 15403 25563 15406
rect 15837 15330 15903 15333
rect 18505 15330 18571 15333
rect 15837 15328 18571 15330
rect 15837 15272 15842 15328
rect 15898 15272 18510 15328
rect 18566 15272 18571 15328
rect 15837 15270 18571 15272
rect 15837 15267 15903 15270
rect 18505 15267 18571 15270
rect 18965 15330 19031 15333
rect 24117 15330 24183 15333
rect 18965 15328 24183 15330
rect 18965 15272 18970 15328
rect 19026 15272 24122 15328
rect 24178 15272 24183 15328
rect 18965 15270 24183 15272
rect 18965 15267 19031 15270
rect 24117 15267 24183 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10777 15194 10843 15197
rect 11329 15194 11395 15197
rect 10777 15192 11395 15194
rect 10777 15136 10782 15192
rect 10838 15136 11334 15192
rect 11390 15136 11395 15192
rect 10777 15134 11395 15136
rect 10777 15131 10843 15134
rect 11329 15131 11395 15134
rect 17677 15194 17743 15197
rect 24117 15194 24183 15197
rect 27520 15194 28000 15224
rect 17677 15192 24183 15194
rect 17677 15136 17682 15192
rect 17738 15136 24122 15192
rect 24178 15136 24183 15192
rect 17677 15134 24183 15136
rect 17677 15131 17743 15134
rect 24117 15131 24183 15134
rect 24902 15134 28000 15194
rect 15745 15058 15811 15061
rect 18321 15058 18387 15061
rect 15745 15056 18387 15058
rect 15745 15000 15750 15056
rect 15806 15000 18326 15056
rect 18382 15000 18387 15056
rect 15745 14998 18387 15000
rect 15745 14995 15811 14998
rect 18321 14995 18387 14998
rect 18781 15058 18847 15061
rect 21357 15058 21423 15061
rect 23197 15058 23263 15061
rect 18781 15056 23263 15058
rect 18781 15000 18786 15056
rect 18842 15000 21362 15056
rect 21418 15000 23202 15056
rect 23258 15000 23263 15056
rect 18781 14998 23263 15000
rect 18781 14995 18847 14998
rect 21357 14995 21423 14998
rect 23197 14995 23263 14998
rect 13813 14922 13879 14925
rect 16389 14922 16455 14925
rect 19609 14922 19675 14925
rect 13813 14920 19675 14922
rect 13813 14864 13818 14920
rect 13874 14864 16394 14920
rect 16450 14864 19614 14920
rect 19670 14864 19675 14920
rect 13813 14862 19675 14864
rect 13813 14859 13879 14862
rect 16389 14859 16455 14862
rect 19609 14859 19675 14862
rect 23473 14922 23539 14925
rect 24902 14922 24962 15134
rect 27520 15104 28000 15134
rect 23473 14920 24962 14922
rect 23473 14864 23478 14920
rect 23534 14864 24962 14920
rect 23473 14862 24962 14864
rect 23473 14859 23539 14862
rect 17033 14786 17099 14789
rect 17350 14786 17356 14788
rect 17033 14784 17356 14786
rect 17033 14728 17038 14784
rect 17094 14728 17356 14784
rect 17033 14726 17356 14728
rect 17033 14723 17099 14726
rect 17350 14724 17356 14726
rect 17420 14724 17426 14788
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 23841 14650 23907 14653
rect 27520 14650 28000 14680
rect 23841 14648 28000 14650
rect 23841 14592 23846 14648
rect 23902 14592 28000 14648
rect 23841 14590 28000 14592
rect 23841 14587 23907 14590
rect 27520 14560 28000 14590
rect 16941 14514 17007 14517
rect 25037 14514 25103 14517
rect 16941 14512 25103 14514
rect 16941 14456 16946 14512
rect 17002 14456 25042 14512
rect 25098 14456 25103 14512
rect 16941 14454 25103 14456
rect 16941 14451 17007 14454
rect 25037 14451 25103 14454
rect 10225 14378 10291 14381
rect 17125 14378 17191 14381
rect 19517 14378 19583 14381
rect 10225 14376 19583 14378
rect 10225 14320 10230 14376
rect 10286 14320 17130 14376
rect 17186 14320 19522 14376
rect 19578 14320 19583 14376
rect 10225 14318 19583 14320
rect 10225 14315 10291 14318
rect 17125 14315 17191 14318
rect 19517 14315 19583 14318
rect 22001 14242 22067 14245
rect 24025 14242 24091 14245
rect 22001 14240 24091 14242
rect 22001 14184 22006 14240
rect 22062 14184 24030 14240
rect 24086 14184 24091 14240
rect 22001 14182 24091 14184
rect 22001 14179 22067 14182
rect 24025 14179 24091 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 15377 14106 15443 14109
rect 20805 14106 20871 14109
rect 15377 14104 20871 14106
rect 15377 14048 15382 14104
rect 15438 14048 20810 14104
rect 20866 14048 20871 14104
rect 15377 14046 20871 14048
rect 15377 14043 15443 14046
rect 20805 14043 20871 14046
rect 4061 13970 4127 13973
rect 23197 13970 23263 13973
rect 4061 13968 23263 13970
rect 4061 13912 4066 13968
rect 4122 13912 23202 13968
rect 23258 13912 23263 13968
rect 4061 13910 23263 13912
rect 4061 13907 4127 13910
rect 23197 13907 23263 13910
rect 25221 13970 25287 13973
rect 27520 13970 28000 14000
rect 25221 13968 28000 13970
rect 25221 13912 25226 13968
rect 25282 13912 28000 13968
rect 25221 13910 28000 13912
rect 25221 13907 25287 13910
rect 27520 13880 28000 13910
rect 13721 13834 13787 13837
rect 15745 13834 15811 13837
rect 13721 13832 15811 13834
rect 13721 13776 13726 13832
rect 13782 13776 15750 13832
rect 15806 13776 15811 13832
rect 13721 13774 15811 13776
rect 13721 13771 13787 13774
rect 15745 13771 15811 13774
rect 18321 13834 18387 13837
rect 20897 13834 20963 13837
rect 18321 13832 20963 13834
rect 18321 13776 18326 13832
rect 18382 13776 20902 13832
rect 20958 13776 20963 13832
rect 18321 13774 20963 13776
rect 18321 13771 18387 13774
rect 20897 13771 20963 13774
rect 14641 13700 14707 13701
rect 14590 13698 14596 13700
rect 14550 13638 14596 13698
rect 14660 13696 14707 13700
rect 14702 13640 14707 13696
rect 14590 13636 14596 13638
rect 14660 13636 14707 13640
rect 14641 13635 14707 13636
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 14641 13562 14707 13565
rect 16481 13562 16547 13565
rect 14641 13560 16547 13562
rect 14641 13504 14646 13560
rect 14702 13504 16486 13560
rect 16542 13504 16547 13560
rect 14641 13502 16547 13504
rect 14641 13499 14707 13502
rect 16481 13499 16547 13502
rect 20069 13562 20135 13565
rect 20069 13560 24962 13562
rect 20069 13504 20074 13560
rect 20130 13504 24962 13560
rect 20069 13502 24962 13504
rect 20069 13499 20135 13502
rect 12893 13426 12959 13429
rect 17493 13426 17559 13429
rect 23473 13426 23539 13429
rect 12893 13424 23539 13426
rect 12893 13368 12898 13424
rect 12954 13368 17498 13424
rect 17554 13368 23478 13424
rect 23534 13368 23539 13424
rect 12893 13366 23539 13368
rect 24902 13426 24962 13502
rect 27520 13426 28000 13456
rect 24902 13366 28000 13426
rect 12893 13363 12959 13366
rect 17493 13363 17559 13366
rect 23473 13363 23539 13366
rect 27520 13336 28000 13366
rect 13077 13290 13143 13293
rect 19609 13290 19675 13293
rect 22829 13290 22895 13293
rect 13077 13288 15394 13290
rect 13077 13232 13082 13288
rect 13138 13232 15394 13288
rect 13077 13230 15394 13232
rect 13077 13227 13143 13230
rect 13997 13154 14063 13157
rect 13862 13152 14063 13154
rect 13862 13096 14002 13152
rect 14058 13096 14063 13152
rect 13862 13094 14063 13096
rect 15334 13154 15394 13230
rect 19609 13288 22895 13290
rect 19609 13232 19614 13288
rect 19670 13232 22834 13288
rect 22890 13232 22895 13288
rect 19609 13230 22895 13232
rect 19609 13227 19675 13230
rect 22829 13227 22895 13230
rect 21081 13154 21147 13157
rect 15334 13152 21147 13154
rect 15334 13096 21086 13152
rect 21142 13096 21147 13152
rect 15334 13094 21147 13096
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 12249 13018 12315 13021
rect 13862 13018 13922 13094
rect 13997 13091 14063 13094
rect 21081 13091 21147 13094
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 12249 13016 13922 13018
rect 12249 12960 12254 13016
rect 12310 12960 13922 13016
rect 12249 12958 13922 12960
rect 18689 13018 18755 13021
rect 20621 13018 20687 13021
rect 18689 13016 20687 13018
rect 18689 12960 18694 13016
rect 18750 12960 20626 13016
rect 20682 12960 20687 13016
rect 18689 12958 20687 12960
rect 12249 12955 12315 12958
rect 18689 12955 18755 12958
rect 20621 12955 20687 12958
rect 10777 12882 10843 12885
rect 12433 12882 12499 12885
rect 10777 12880 12499 12882
rect 10777 12824 10782 12880
rect 10838 12824 12438 12880
rect 12494 12824 12499 12880
rect 10777 12822 12499 12824
rect 10777 12819 10843 12822
rect 12433 12819 12499 12822
rect 13169 12882 13235 12885
rect 17861 12882 17927 12885
rect 13169 12880 17927 12882
rect 13169 12824 13174 12880
rect 13230 12824 17866 12880
rect 17922 12824 17927 12880
rect 13169 12822 17927 12824
rect 13169 12819 13235 12822
rect 17861 12819 17927 12822
rect 18873 12882 18939 12885
rect 21081 12882 21147 12885
rect 18873 12880 21147 12882
rect 18873 12824 18878 12880
rect 18934 12824 21086 12880
rect 21142 12824 21147 12880
rect 18873 12822 21147 12824
rect 18873 12819 18939 12822
rect 21081 12819 21147 12822
rect 24025 12882 24091 12885
rect 27520 12882 28000 12912
rect 24025 12880 28000 12882
rect 24025 12824 24030 12880
rect 24086 12824 28000 12880
rect 24025 12822 28000 12824
rect 24025 12819 24091 12822
rect 27520 12792 28000 12822
rect 16113 12746 16179 12749
rect 22553 12746 22619 12749
rect 16113 12744 22619 12746
rect 16113 12688 16118 12744
rect 16174 12688 22558 12744
rect 22614 12688 22619 12744
rect 16113 12686 22619 12688
rect 16113 12683 16179 12686
rect 22553 12683 22619 12686
rect 14457 12610 14523 12613
rect 14825 12610 14891 12613
rect 14457 12608 14891 12610
rect 14457 12552 14462 12608
rect 14518 12552 14830 12608
rect 14886 12552 14891 12608
rect 14457 12550 14891 12552
rect 14457 12547 14523 12550
rect 14825 12547 14891 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 11973 12474 12039 12477
rect 17166 12474 17172 12476
rect 11973 12472 17172 12474
rect 11973 12416 11978 12472
rect 12034 12416 17172 12472
rect 11973 12414 17172 12416
rect 11973 12411 12039 12414
rect 17166 12412 17172 12414
rect 17236 12412 17242 12476
rect 12525 12338 12591 12341
rect 15929 12338 15995 12341
rect 12525 12336 15995 12338
rect 12525 12280 12530 12336
rect 12586 12280 15934 12336
rect 15990 12280 15995 12336
rect 12525 12278 15995 12280
rect 12525 12275 12591 12278
rect 15929 12275 15995 12278
rect 16205 12338 16271 12341
rect 23841 12338 23907 12341
rect 16205 12336 23907 12338
rect 16205 12280 16210 12336
rect 16266 12280 23846 12336
rect 23902 12280 23907 12336
rect 16205 12278 23907 12280
rect 16205 12275 16271 12278
rect 23841 12275 23907 12278
rect 24209 12338 24275 12341
rect 27520 12338 28000 12368
rect 24209 12336 28000 12338
rect 24209 12280 24214 12336
rect 24270 12280 28000 12336
rect 24209 12278 28000 12280
rect 24209 12275 24275 12278
rect 27520 12248 28000 12278
rect 15101 12202 15167 12205
rect 16757 12202 16823 12205
rect 15101 12200 16823 12202
rect 15101 12144 15106 12200
rect 15162 12144 16762 12200
rect 16818 12144 16823 12200
rect 15101 12142 16823 12144
rect 15101 12139 15167 12142
rect 16757 12139 16823 12142
rect 17125 12204 17191 12205
rect 17125 12200 17172 12204
rect 17236 12202 17242 12204
rect 17125 12144 17130 12200
rect 17125 12140 17172 12144
rect 17236 12142 17282 12202
rect 17236 12140 17242 12142
rect 17125 12139 17191 12140
rect 17350 12004 17356 12068
rect 17420 12066 17426 12068
rect 17493 12066 17559 12069
rect 17420 12064 17559 12066
rect 17420 12008 17498 12064
rect 17554 12008 17559 12064
rect 17420 12006 17559 12008
rect 17420 12004 17426 12006
rect 17493 12003 17559 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 22001 11794 22067 11797
rect 27520 11794 28000 11824
rect 22001 11792 28000 11794
rect 22001 11736 22006 11792
rect 22062 11736 28000 11792
rect 22001 11734 28000 11736
rect 22001 11731 22067 11734
rect 27520 11704 28000 11734
rect 10777 11658 10843 11661
rect 12433 11658 12499 11661
rect 10777 11656 12499 11658
rect 10777 11600 10782 11656
rect 10838 11600 12438 11656
rect 12494 11600 12499 11656
rect 10777 11598 12499 11600
rect 10777 11595 10843 11598
rect 12433 11595 12499 11598
rect 13261 11658 13327 11661
rect 17677 11658 17743 11661
rect 13261 11656 17743 11658
rect 13261 11600 13266 11656
rect 13322 11600 17682 11656
rect 17738 11600 17743 11656
rect 13261 11598 17743 11600
rect 13261 11595 13327 11598
rect 17677 11595 17743 11598
rect 17309 11522 17375 11525
rect 19333 11522 19399 11525
rect 17309 11520 19399 11522
rect 17309 11464 17314 11520
rect 17370 11464 19338 11520
rect 19394 11464 19399 11520
rect 17309 11462 19399 11464
rect 17309 11459 17375 11462
rect 19333 11459 19399 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 13629 11386 13695 11389
rect 13629 11384 19074 11386
rect 13629 11328 13634 11384
rect 13690 11328 19074 11384
rect 13629 11326 19074 11328
rect 13629 11323 13695 11326
rect 14733 11250 14799 11253
rect 15929 11250 15995 11253
rect 18873 11250 18939 11253
rect 14733 11248 18939 11250
rect 14733 11192 14738 11248
rect 14794 11192 15934 11248
rect 15990 11192 18878 11248
rect 18934 11192 18939 11248
rect 14733 11190 18939 11192
rect 19014 11250 19074 11326
rect 25313 11250 25379 11253
rect 19014 11248 25379 11250
rect 19014 11192 25318 11248
rect 25374 11192 25379 11248
rect 19014 11190 25379 11192
rect 14733 11187 14799 11190
rect 15929 11187 15995 11190
rect 18873 11187 18939 11190
rect 25313 11187 25379 11190
rect 7741 11114 7807 11117
rect 14457 11114 14523 11117
rect 7741 11112 14523 11114
rect 7741 11056 7746 11112
rect 7802 11056 14462 11112
rect 14518 11056 14523 11112
rect 7741 11054 14523 11056
rect 7741 11051 7807 11054
rect 14457 11051 14523 11054
rect 17953 11114 18019 11117
rect 19701 11114 19767 11117
rect 27520 11114 28000 11144
rect 17953 11112 19767 11114
rect 17953 11056 17958 11112
rect 18014 11056 19706 11112
rect 19762 11056 19767 11112
rect 17953 11054 19767 11056
rect 17953 11051 18019 11054
rect 19701 11051 19767 11054
rect 19934 11054 28000 11114
rect 14457 10978 14523 10981
rect 14590 10978 14596 10980
rect 14457 10976 14596 10978
rect 14457 10920 14462 10976
rect 14518 10920 14596 10976
rect 14457 10918 14596 10920
rect 14457 10915 14523 10918
rect 14590 10916 14596 10918
rect 14660 10916 14666 10980
rect 19149 10978 19215 10981
rect 19934 10978 19994 11054
rect 27520 11024 28000 11054
rect 19149 10976 19994 10978
rect 19149 10920 19154 10976
rect 19210 10920 19994 10976
rect 19149 10918 19994 10920
rect 19149 10915 19215 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 12893 10706 12959 10709
rect 18597 10706 18663 10709
rect 12893 10704 18663 10706
rect 12893 10648 12898 10704
rect 12954 10648 18602 10704
rect 18658 10648 18663 10704
rect 12893 10646 18663 10648
rect 12893 10643 12959 10646
rect 18597 10643 18663 10646
rect 14825 10570 14891 10573
rect 20989 10570 21055 10573
rect 27520 10570 28000 10600
rect 14825 10568 21055 10570
rect 14825 10512 14830 10568
rect 14886 10512 20994 10568
rect 21050 10512 21055 10568
rect 14825 10510 21055 10512
rect 14825 10507 14891 10510
rect 20989 10507 21055 10510
rect 24902 10510 28000 10570
rect 10961 10434 11027 10437
rect 13997 10434 14063 10437
rect 10961 10432 14063 10434
rect 10961 10376 10966 10432
rect 11022 10376 14002 10432
rect 14058 10376 14063 10432
rect 10961 10374 14063 10376
rect 10961 10371 11027 10374
rect 13997 10371 14063 10374
rect 20069 10434 20135 10437
rect 23013 10434 23079 10437
rect 20069 10432 23079 10434
rect 20069 10376 20074 10432
rect 20130 10376 23018 10432
rect 23074 10376 23079 10432
rect 20069 10374 23079 10376
rect 20069 10371 20135 10374
rect 23013 10371 23079 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 12433 10298 12499 10301
rect 17309 10298 17375 10301
rect 17677 10298 17743 10301
rect 12433 10296 17743 10298
rect 12433 10240 12438 10296
rect 12494 10240 17314 10296
rect 17370 10240 17682 10296
rect 17738 10240 17743 10296
rect 12433 10238 17743 10240
rect 12433 10235 12499 10238
rect 17309 10235 17375 10238
rect 17677 10235 17743 10238
rect 20161 10298 20227 10301
rect 24117 10298 24183 10301
rect 20161 10296 24183 10298
rect 20161 10240 20166 10296
rect 20222 10240 24122 10296
rect 24178 10240 24183 10296
rect 20161 10238 24183 10240
rect 20161 10235 20227 10238
rect 24117 10235 24183 10238
rect 16113 10162 16179 10165
rect 24902 10162 24962 10510
rect 27520 10480 28000 10510
rect 16113 10160 24962 10162
rect 16113 10104 16118 10160
rect 16174 10104 24962 10160
rect 16113 10102 24962 10104
rect 16113 10099 16179 10102
rect 16021 10026 16087 10029
rect 21081 10026 21147 10029
rect 27520 10026 28000 10056
rect 16021 10024 21147 10026
rect 16021 9968 16026 10024
rect 16082 9968 21086 10024
rect 21142 9968 21147 10024
rect 16021 9966 21147 9968
rect 16021 9963 16087 9966
rect 21081 9963 21147 9966
rect 24166 9966 28000 10026
rect 24166 9924 24226 9966
rect 27520 9936 28000 9966
rect 24120 9864 24226 9924
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24120 9757 24180 9864
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 24117 9752 24183 9757
rect 24117 9696 24122 9752
rect 24178 9696 24183 9752
rect 24117 9691 24183 9696
rect 17861 9618 17927 9621
rect 19425 9618 19491 9621
rect 17861 9616 19491 9618
rect 17861 9560 17866 9616
rect 17922 9560 19430 9616
rect 19486 9560 19491 9616
rect 17861 9558 19491 9560
rect 17861 9555 17927 9558
rect 19425 9555 19491 9558
rect 22369 9618 22435 9621
rect 25405 9618 25471 9621
rect 22369 9616 25471 9618
rect 22369 9560 22374 9616
rect 22430 9560 25410 9616
rect 25466 9560 25471 9616
rect 22369 9558 25471 9560
rect 22369 9555 22435 9558
rect 25405 9555 25471 9558
rect 16849 9482 16915 9485
rect 23013 9482 23079 9485
rect 16849 9480 23079 9482
rect 16849 9424 16854 9480
rect 16910 9424 23018 9480
rect 23074 9424 23079 9480
rect 16849 9422 23079 9424
rect 16849 9419 16915 9422
rect 23013 9419 23079 9422
rect 23749 9482 23815 9485
rect 27520 9482 28000 9512
rect 23749 9480 28000 9482
rect 23749 9424 23754 9480
rect 23810 9424 28000 9480
rect 23749 9422 28000 9424
rect 23749 9419 23815 9422
rect 27520 9392 28000 9422
rect 10777 9346 10843 9349
rect 12893 9346 12959 9349
rect 10777 9344 12959 9346
rect 10777 9288 10782 9344
rect 10838 9288 12898 9344
rect 12954 9288 12959 9344
rect 10777 9286 12959 9288
rect 10777 9283 10843 9286
rect 12893 9283 12959 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 20069 9210 20135 9213
rect 23473 9210 23539 9213
rect 20069 9208 23539 9210
rect 20069 9152 20074 9208
rect 20130 9152 23478 9208
rect 23534 9152 23539 9208
rect 20069 9150 23539 9152
rect 20069 9147 20135 9150
rect 23473 9147 23539 9150
rect 17953 9074 18019 9077
rect 20897 9074 20963 9077
rect 17953 9072 20963 9074
rect 17953 9016 17958 9072
rect 18014 9016 20902 9072
rect 20958 9016 20963 9072
rect 17953 9014 20963 9016
rect 17953 9011 18019 9014
rect 20897 9011 20963 9014
rect 12893 8938 12959 8941
rect 17401 8938 17467 8941
rect 12893 8936 17467 8938
rect 12893 8880 12898 8936
rect 12954 8880 17406 8936
rect 17462 8880 17467 8936
rect 12893 8878 17467 8880
rect 12893 8875 12959 8878
rect 17401 8875 17467 8878
rect 23841 8936 23907 8941
rect 23841 8880 23846 8936
rect 23902 8880 23907 8936
rect 23841 8875 23907 8880
rect 24761 8938 24827 8941
rect 27520 8938 28000 8968
rect 24761 8936 28000 8938
rect 24761 8880 24766 8936
rect 24822 8880 28000 8936
rect 24761 8878 28000 8880
rect 24761 8875 24827 8878
rect 17861 8802 17927 8805
rect 20713 8802 20779 8805
rect 23844 8802 23904 8875
rect 27520 8848 28000 8878
rect 17861 8800 20779 8802
rect 17861 8744 17866 8800
rect 17922 8744 20718 8800
rect 20774 8744 20779 8800
rect 17861 8742 20779 8744
rect 17861 8739 17927 8742
rect 20713 8739 20779 8742
rect 21590 8742 23904 8802
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 15469 8666 15535 8669
rect 21590 8666 21650 8742
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 15334 8664 21650 8666
rect 15334 8608 15474 8664
rect 15530 8608 21650 8664
rect 15334 8606 21650 8608
rect 13261 8530 13327 8533
rect 15334 8530 15394 8606
rect 15469 8603 15535 8606
rect 13261 8528 15394 8530
rect 13261 8472 13266 8528
rect 13322 8472 15394 8528
rect 13261 8470 15394 8472
rect 17493 8530 17559 8533
rect 19977 8530 20043 8533
rect 17493 8528 20043 8530
rect 17493 8472 17498 8528
rect 17554 8472 19982 8528
rect 20038 8472 20043 8528
rect 17493 8470 20043 8472
rect 13261 8467 13327 8470
rect 17493 8467 17559 8470
rect 19977 8467 20043 8470
rect 3693 8394 3759 8397
rect 11329 8394 11395 8397
rect 3693 8392 11395 8394
rect 3693 8336 3698 8392
rect 3754 8336 11334 8392
rect 11390 8336 11395 8392
rect 3693 8334 11395 8336
rect 3693 8331 3759 8334
rect 11329 8331 11395 8334
rect 24209 8258 24275 8261
rect 27520 8258 28000 8288
rect 24209 8256 28000 8258
rect 24209 8200 24214 8256
rect 24270 8200 28000 8256
rect 24209 8198 28000 8200
rect 24209 8195 24275 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 15745 8122 15811 8125
rect 16205 8122 16271 8125
rect 15745 8120 16271 8122
rect 15745 8064 15750 8120
rect 15806 8064 16210 8120
rect 16266 8064 16271 8120
rect 15745 8062 16271 8064
rect 15745 8059 15811 8062
rect 16205 8059 16271 8062
rect 15377 7986 15443 7989
rect 22093 7986 22159 7989
rect 15377 7984 22159 7986
rect 15377 7928 15382 7984
rect 15438 7928 22098 7984
rect 22154 7928 22159 7984
rect 15377 7926 22159 7928
rect 15377 7923 15443 7926
rect 22093 7923 22159 7926
rect 23473 7986 23539 7989
rect 23473 7984 24778 7986
rect 23473 7928 23478 7984
rect 23534 7928 24778 7984
rect 23473 7926 24778 7928
rect 23473 7923 23539 7926
rect 9857 7850 9923 7853
rect 12433 7850 12499 7853
rect 9857 7848 12499 7850
rect 9857 7792 9862 7848
rect 9918 7792 12438 7848
rect 12494 7792 12499 7848
rect 9857 7790 12499 7792
rect 9857 7787 9923 7790
rect 12433 7787 12499 7790
rect 14365 7850 14431 7853
rect 15929 7850 15995 7853
rect 14365 7848 15995 7850
rect 14365 7792 14370 7848
rect 14426 7792 15934 7848
rect 15990 7792 15995 7848
rect 14365 7790 15995 7792
rect 14365 7787 14431 7790
rect 15929 7787 15995 7790
rect 18597 7850 18663 7853
rect 23749 7850 23815 7853
rect 18597 7848 23815 7850
rect 18597 7792 18602 7848
rect 18658 7792 23754 7848
rect 23810 7792 23815 7848
rect 18597 7790 23815 7792
rect 18597 7787 18663 7790
rect 23749 7787 23815 7790
rect 11329 7714 11395 7717
rect 13905 7714 13971 7717
rect 11329 7712 13971 7714
rect 11329 7656 11334 7712
rect 11390 7656 13910 7712
rect 13966 7656 13971 7712
rect 11329 7654 13971 7656
rect 24718 7714 24778 7926
rect 27520 7714 28000 7744
rect 24718 7654 28000 7714
rect 11329 7651 11395 7654
rect 13905 7651 13971 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 16205 7578 16271 7581
rect 21817 7578 21883 7581
rect 16205 7576 21883 7578
rect 16205 7520 16210 7576
rect 16266 7520 21822 7576
rect 21878 7520 21883 7576
rect 16205 7518 21883 7520
rect 16205 7515 16271 7518
rect 21817 7515 21883 7518
rect 289 7442 355 7445
rect 10593 7442 10659 7445
rect 289 7440 10659 7442
rect 289 7384 294 7440
rect 350 7384 10598 7440
rect 10654 7384 10659 7440
rect 289 7382 10659 7384
rect 289 7379 355 7382
rect 10593 7379 10659 7382
rect 10869 7442 10935 7445
rect 13721 7442 13787 7445
rect 24025 7442 24091 7445
rect 10869 7440 24091 7442
rect 10869 7384 10874 7440
rect 10930 7384 13726 7440
rect 13782 7384 24030 7440
rect 24086 7384 24091 7440
rect 10869 7382 24091 7384
rect 10869 7379 10935 7382
rect 13721 7379 13787 7382
rect 24025 7379 24091 7382
rect 18689 7306 18755 7309
rect 23105 7306 23171 7309
rect 23565 7306 23631 7309
rect 18689 7304 22018 7306
rect 18689 7248 18694 7304
rect 18750 7272 22018 7304
rect 23105 7304 23631 7306
rect 18750 7248 22202 7272
rect 18689 7246 22202 7248
rect 18689 7243 18755 7246
rect 21958 7212 22202 7246
rect 23105 7248 23110 7304
rect 23166 7248 23570 7304
rect 23626 7248 23631 7304
rect 23105 7246 23631 7248
rect 23105 7243 23171 7246
rect 23565 7243 23631 7246
rect 15837 7170 15903 7173
rect 17953 7170 18019 7173
rect 15837 7168 18019 7170
rect 15837 7112 15842 7168
rect 15898 7112 17958 7168
rect 18014 7112 18019 7168
rect 15837 7110 18019 7112
rect 22142 7170 22202 7212
rect 27520 7170 28000 7200
rect 22142 7110 28000 7170
rect 15837 7107 15903 7110
rect 17953 7107 18019 7110
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 27520 7080 28000 7110
rect 19610 7039 19930 7040
rect 565 7034 631 7037
rect 0 7032 631 7034
rect 0 6976 570 7032
rect 626 6976 631 7032
rect 0 6974 631 6976
rect 0 6944 480 6974
rect 565 6971 631 6974
rect 12801 7034 12867 7037
rect 17861 7034 17927 7037
rect 12801 7032 17927 7034
rect 12801 6976 12806 7032
rect 12862 6976 17866 7032
rect 17922 6976 17927 7032
rect 12801 6974 17927 6976
rect 12801 6971 12867 6974
rect 17861 6971 17927 6974
rect 22369 7034 22435 7037
rect 25313 7034 25379 7037
rect 22369 7032 25379 7034
rect 22369 6976 22374 7032
rect 22430 6976 25318 7032
rect 25374 6976 25379 7032
rect 22369 6974 25379 6976
rect 22369 6971 22435 6974
rect 25313 6971 25379 6974
rect 18137 6898 18203 6901
rect 20161 6898 20227 6901
rect 18137 6896 20227 6898
rect 18137 6840 18142 6896
rect 18198 6840 20166 6896
rect 20222 6840 20227 6896
rect 18137 6838 20227 6840
rect 18137 6835 18203 6838
rect 20161 6835 20227 6838
rect 4337 6762 4403 6765
rect 13445 6762 13511 6765
rect 4337 6760 13511 6762
rect 4337 6704 4342 6760
rect 4398 6704 13450 6760
rect 13506 6704 13511 6760
rect 4337 6702 13511 6704
rect 4337 6699 4403 6702
rect 13445 6699 13511 6702
rect 22645 6762 22711 6765
rect 22645 6760 24778 6762
rect 22645 6704 22650 6760
rect 22706 6704 24778 6760
rect 22645 6702 24778 6704
rect 22645 6699 22711 6702
rect 19977 6626 20043 6629
rect 22001 6626 22067 6629
rect 19977 6624 22067 6626
rect 19977 6568 19982 6624
rect 20038 6568 22006 6624
rect 22062 6568 22067 6624
rect 19977 6566 22067 6568
rect 24718 6626 24778 6702
rect 27520 6626 28000 6656
rect 24718 6566 28000 6626
rect 19977 6563 20043 6566
rect 22001 6563 22067 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 21909 6354 21975 6357
rect 23013 6354 23079 6357
rect 21909 6352 23079 6354
rect 21909 6296 21914 6352
rect 21970 6296 23018 6352
rect 23074 6296 23079 6352
rect 21909 6294 23079 6296
rect 21909 6291 21975 6294
rect 23013 6291 23079 6294
rect 13261 6218 13327 6221
rect 13261 6216 20132 6218
rect 13261 6160 13266 6216
rect 13322 6160 20132 6216
rect 13261 6158 20132 6160
rect 13261 6155 13327 6158
rect 11329 6082 11395 6085
rect 14733 6082 14799 6085
rect 11329 6080 14799 6082
rect 11329 6024 11334 6080
rect 11390 6024 14738 6080
rect 14794 6024 14799 6080
rect 11329 6022 14799 6024
rect 20072 6082 20132 6158
rect 27520 6082 28000 6112
rect 20072 6022 28000 6082
rect 11329 6019 11395 6022
rect 14733 6019 14799 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 12433 5810 12499 5813
rect 20713 5810 20779 5813
rect 12433 5808 20779 5810
rect 12433 5752 12438 5808
rect 12494 5752 20718 5808
rect 20774 5752 20779 5808
rect 12433 5750 20779 5752
rect 12433 5747 12499 5750
rect 20713 5747 20779 5750
rect 2313 5674 2379 5677
rect 10777 5674 10843 5677
rect 2313 5672 10843 5674
rect 2313 5616 2318 5672
rect 2374 5616 10782 5672
rect 10838 5616 10843 5672
rect 2313 5614 10843 5616
rect 2313 5611 2379 5614
rect 10777 5611 10843 5614
rect 11053 5674 11119 5677
rect 16757 5674 16823 5677
rect 11053 5672 16823 5674
rect 11053 5616 11058 5672
rect 11114 5616 16762 5672
rect 16818 5616 16823 5672
rect 11053 5614 16823 5616
rect 11053 5611 11119 5614
rect 16757 5611 16823 5614
rect 17033 5674 17099 5677
rect 20069 5674 20135 5677
rect 17033 5672 20135 5674
rect 17033 5616 17038 5672
rect 17094 5616 20074 5672
rect 20130 5616 20135 5672
rect 17033 5614 20135 5616
rect 17033 5611 17099 5614
rect 20069 5611 20135 5614
rect 23289 5674 23355 5677
rect 25037 5674 25103 5677
rect 23289 5672 25103 5674
rect 23289 5616 23294 5672
rect 23350 5616 25042 5672
rect 25098 5616 25103 5672
rect 23289 5614 25103 5616
rect 23289 5611 23355 5614
rect 25037 5611 25103 5614
rect 9765 5538 9831 5541
rect 12341 5538 12407 5541
rect 9765 5536 12407 5538
rect 9765 5480 9770 5536
rect 9826 5480 12346 5536
rect 12402 5480 12407 5536
rect 9765 5478 12407 5480
rect 9765 5475 9831 5478
rect 12341 5475 12407 5478
rect 19517 5538 19583 5541
rect 21357 5538 21423 5541
rect 19517 5536 21423 5538
rect 19517 5480 19522 5536
rect 19578 5480 21362 5536
rect 21418 5480 21423 5536
rect 19517 5478 21423 5480
rect 19517 5475 19583 5478
rect 21357 5475 21423 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 16389 5402 16455 5405
rect 18689 5402 18755 5405
rect 27520 5402 28000 5432
rect 16389 5400 23536 5402
rect 16389 5344 16394 5400
rect 16450 5344 18694 5400
rect 18750 5344 23536 5400
rect 16389 5342 23536 5344
rect 16389 5339 16455 5342
rect 18689 5339 18755 5342
rect 2957 5266 3023 5269
rect 19609 5266 19675 5269
rect 2957 5264 19675 5266
rect 2957 5208 2962 5264
rect 3018 5208 19614 5264
rect 19670 5208 19675 5264
rect 2957 5206 19675 5208
rect 23476 5266 23536 5342
rect 24672 5342 28000 5402
rect 24672 5266 24732 5342
rect 27520 5312 28000 5342
rect 23476 5206 24732 5266
rect 2957 5203 3023 5206
rect 19609 5203 19675 5206
rect 7649 5130 7715 5133
rect 13261 5130 13327 5133
rect 15837 5130 15903 5133
rect 7649 5128 10794 5130
rect 7649 5072 7654 5128
rect 7710 5072 10794 5128
rect 7649 5070 10794 5072
rect 7649 5067 7715 5070
rect 10734 4994 10794 5070
rect 13261 5128 15903 5130
rect 13261 5072 13266 5128
rect 13322 5072 15842 5128
rect 15898 5072 15903 5128
rect 13261 5070 15903 5072
rect 13261 5067 13327 5070
rect 15837 5067 15903 5070
rect 18781 5130 18847 5133
rect 25497 5130 25563 5133
rect 18781 5128 25563 5130
rect 18781 5072 18786 5128
rect 18842 5072 25502 5128
rect 25558 5072 25563 5128
rect 18781 5070 25563 5072
rect 18781 5067 18847 5070
rect 25497 5067 25563 5070
rect 11605 4994 11671 4997
rect 18689 4994 18755 4997
rect 10734 4992 18755 4994
rect 10734 4936 11610 4992
rect 11666 4936 18694 4992
rect 18750 4936 18755 4992
rect 10734 4934 18755 4936
rect 11605 4931 11671 4934
rect 18689 4931 18755 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 20253 4858 20319 4861
rect 22829 4858 22895 4861
rect 20253 4856 22895 4858
rect 20253 4800 20258 4856
rect 20314 4800 22834 4856
rect 22890 4800 22895 4856
rect 20253 4798 22895 4800
rect 20253 4795 20319 4798
rect 22829 4795 22895 4798
rect 25037 4858 25103 4861
rect 27520 4858 28000 4888
rect 25037 4856 28000 4858
rect 25037 4800 25042 4856
rect 25098 4800 28000 4856
rect 25037 4798 28000 4800
rect 25037 4795 25103 4798
rect 27520 4768 28000 4798
rect 17033 4722 17099 4725
rect 22185 4722 22251 4725
rect 17033 4720 22251 4722
rect 17033 4664 17038 4720
rect 17094 4664 22190 4720
rect 22246 4664 22251 4720
rect 17033 4662 22251 4664
rect 17033 4659 17099 4662
rect 22185 4659 22251 4662
rect 14273 4586 14339 4589
rect 19333 4586 19399 4589
rect 14273 4584 19399 4586
rect 14273 4528 14278 4584
rect 14334 4528 19338 4584
rect 19394 4528 19399 4584
rect 14273 4526 19399 4528
rect 14273 4523 14339 4526
rect 19333 4523 19399 4526
rect 22645 4586 22711 4589
rect 25497 4586 25563 4589
rect 22645 4584 25563 4586
rect 22645 4528 22650 4584
rect 22706 4528 25502 4584
rect 25558 4528 25563 4584
rect 22645 4526 25563 4528
rect 22645 4523 22711 4526
rect 25497 4523 25563 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 16113 4314 16179 4317
rect 20897 4314 20963 4317
rect 16113 4312 20963 4314
rect 16113 4256 16118 4312
rect 16174 4256 20902 4312
rect 20958 4256 20963 4312
rect 16113 4254 20963 4256
rect 16113 4251 16179 4254
rect 20897 4251 20963 4254
rect 26049 4314 26115 4317
rect 27520 4314 28000 4344
rect 26049 4312 28000 4314
rect 26049 4256 26054 4312
rect 26110 4256 28000 4312
rect 26049 4254 28000 4256
rect 26049 4251 26115 4254
rect 27520 4224 28000 4254
rect 9581 4178 9647 4181
rect 22093 4178 22159 4181
rect 24761 4178 24827 4181
rect 9581 4176 22018 4178
rect 9581 4120 9586 4176
rect 9642 4120 22018 4176
rect 9581 4118 22018 4120
rect 9581 4115 9647 4118
rect 1393 4042 1459 4045
rect 11329 4042 11395 4045
rect 1393 4040 11395 4042
rect 1393 3984 1398 4040
rect 1454 3984 11334 4040
rect 11390 3984 11395 4040
rect 1393 3982 11395 3984
rect 1393 3979 1459 3982
rect 11329 3979 11395 3982
rect 11513 4042 11579 4045
rect 15929 4042 15995 4045
rect 11513 4040 15995 4042
rect 11513 3984 11518 4040
rect 11574 3984 15934 4040
rect 15990 3984 15995 4040
rect 11513 3982 15995 3984
rect 11513 3979 11579 3982
rect 15929 3979 15995 3982
rect 19241 4042 19307 4045
rect 21725 4042 21791 4045
rect 19241 4040 21791 4042
rect 19241 3984 19246 4040
rect 19302 3984 21730 4040
rect 21786 3984 21791 4040
rect 19241 3982 21791 3984
rect 21958 4042 22018 4118
rect 22093 4176 24827 4178
rect 22093 4120 22098 4176
rect 22154 4120 24766 4176
rect 24822 4120 24827 4176
rect 22093 4118 24827 4120
rect 22093 4115 22159 4118
rect 24761 4115 24827 4118
rect 24393 4042 24459 4045
rect 21958 4040 24459 4042
rect 21958 3984 24398 4040
rect 24454 3984 24459 4040
rect 21958 3982 24459 3984
rect 19241 3979 19307 3982
rect 21725 3979 21791 3982
rect 24393 3979 24459 3982
rect 6361 3906 6427 3909
rect 10041 3906 10107 3909
rect 6361 3904 10107 3906
rect 6361 3848 6366 3904
rect 6422 3848 10046 3904
rect 10102 3848 10107 3904
rect 6361 3846 10107 3848
rect 6361 3843 6427 3846
rect 10041 3843 10107 3846
rect 11145 3906 11211 3909
rect 15561 3906 15627 3909
rect 11145 3904 15627 3906
rect 11145 3848 11150 3904
rect 11206 3848 15566 3904
rect 15622 3848 15627 3904
rect 11145 3846 15627 3848
rect 11145 3843 11211 3846
rect 15561 3843 15627 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 12617 3770 12683 3773
rect 16573 3770 16639 3773
rect 12617 3768 16639 3770
rect 12617 3712 12622 3768
rect 12678 3712 16578 3768
rect 16634 3712 16639 3768
rect 12617 3710 16639 3712
rect 12617 3707 12683 3710
rect 16573 3707 16639 3710
rect 24669 3770 24735 3773
rect 27520 3770 28000 3800
rect 24669 3768 28000 3770
rect 24669 3712 24674 3768
rect 24730 3712 28000 3768
rect 24669 3710 28000 3712
rect 24669 3707 24735 3710
rect 27520 3680 28000 3710
rect 7097 3634 7163 3637
rect 10133 3634 10199 3637
rect 7097 3632 10199 3634
rect 7097 3576 7102 3632
rect 7158 3576 10138 3632
rect 10194 3576 10199 3632
rect 7097 3574 10199 3576
rect 7097 3571 7163 3574
rect 10133 3571 10199 3574
rect 11145 3634 11211 3637
rect 13813 3634 13879 3637
rect 11145 3632 13879 3634
rect 11145 3576 11150 3632
rect 11206 3576 13818 3632
rect 13874 3576 13879 3632
rect 11145 3574 13879 3576
rect 11145 3571 11211 3574
rect 13813 3571 13879 3574
rect 15193 3634 15259 3637
rect 25589 3634 25655 3637
rect 15193 3632 25655 3634
rect 15193 3576 15198 3632
rect 15254 3576 25594 3632
rect 25650 3576 25655 3632
rect 15193 3574 25655 3576
rect 15193 3571 15259 3574
rect 25589 3571 25655 3574
rect 10777 3498 10843 3501
rect 16665 3498 16731 3501
rect 10777 3496 16731 3498
rect 10777 3440 10782 3496
rect 10838 3440 16670 3496
rect 16726 3440 16731 3496
rect 10777 3438 16731 3440
rect 10777 3435 10843 3438
rect 16665 3435 16731 3438
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 11421 3226 11487 3229
rect 14549 3226 14615 3229
rect 11421 3224 14615 3226
rect 11421 3168 11426 3224
rect 11482 3168 14554 3224
rect 14610 3168 14615 3224
rect 11421 3166 14615 3168
rect 11421 3163 11487 3166
rect 14549 3163 14615 3166
rect 18045 3226 18111 3229
rect 21725 3226 21791 3229
rect 27520 3226 28000 3256
rect 18045 3224 21791 3226
rect 18045 3168 18050 3224
rect 18106 3168 21730 3224
rect 21786 3168 21791 3224
rect 18045 3166 21791 3168
rect 18045 3163 18111 3166
rect 21725 3163 21791 3166
rect 24718 3166 28000 3226
rect 4981 3090 5047 3093
rect 11053 3090 11119 3093
rect 4981 3088 11119 3090
rect 4981 3032 4986 3088
rect 5042 3032 11058 3088
rect 11114 3032 11119 3088
rect 4981 3030 11119 3032
rect 4981 3027 5047 3030
rect 11053 3027 11119 3030
rect 11421 3090 11487 3093
rect 17953 3090 18019 3093
rect 11421 3088 18019 3090
rect 11421 3032 11426 3088
rect 11482 3032 17958 3088
rect 18014 3032 18019 3088
rect 11421 3030 18019 3032
rect 11421 3027 11487 3030
rect 17953 3027 18019 3030
rect 23841 3090 23907 3093
rect 24718 3090 24778 3166
rect 27520 3136 28000 3166
rect 23841 3088 24778 3090
rect 23841 3032 23846 3088
rect 23902 3032 24778 3088
rect 23841 3030 24778 3032
rect 23841 3027 23907 3030
rect 8385 2954 8451 2957
rect 12525 2954 12591 2957
rect 8385 2952 12591 2954
rect 8385 2896 8390 2952
rect 8446 2896 12530 2952
rect 12586 2896 12591 2952
rect 8385 2894 12591 2896
rect 8385 2891 8451 2894
rect 12525 2891 12591 2894
rect 13629 2954 13695 2957
rect 18689 2954 18755 2957
rect 13629 2952 18755 2954
rect 13629 2896 13634 2952
rect 13690 2896 18694 2952
rect 18750 2896 18755 2952
rect 13629 2894 18755 2896
rect 13629 2891 13695 2894
rect 18689 2891 18755 2894
rect 10869 2818 10935 2821
rect 15285 2818 15351 2821
rect 10869 2816 15351 2818
rect 10869 2760 10874 2816
rect 10930 2760 15290 2816
rect 15346 2760 15351 2816
rect 10869 2758 15351 2760
rect 10869 2755 10935 2758
rect 15285 2755 15351 2758
rect 16297 2818 16363 2821
rect 18505 2818 18571 2821
rect 16297 2816 18571 2818
rect 16297 2760 16302 2816
rect 16358 2760 18510 2816
rect 18566 2760 18571 2816
rect 16297 2758 18571 2760
rect 16297 2755 16363 2758
rect 18505 2755 18571 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 10869 2682 10935 2685
rect 17033 2682 17099 2685
rect 10869 2680 17099 2682
rect 10869 2624 10874 2680
rect 10930 2624 17038 2680
rect 17094 2624 17099 2680
rect 10869 2622 17099 2624
rect 10869 2619 10935 2622
rect 17033 2619 17099 2622
rect 21265 2682 21331 2685
rect 23565 2682 23631 2685
rect 21265 2680 23631 2682
rect 21265 2624 21270 2680
rect 21326 2624 23570 2680
rect 23626 2624 23631 2680
rect 21265 2622 23631 2624
rect 21265 2619 21331 2622
rect 23565 2619 23631 2622
rect 1577 2546 1643 2549
rect 20897 2546 20963 2549
rect 1577 2544 20963 2546
rect 1577 2488 1582 2544
rect 1638 2488 20902 2544
rect 20958 2488 20963 2544
rect 1577 2486 20963 2488
rect 1577 2483 1643 2486
rect 20897 2483 20963 2486
rect 23749 2546 23815 2549
rect 27520 2546 28000 2576
rect 23749 2544 28000 2546
rect 23749 2488 23754 2544
rect 23810 2488 28000 2544
rect 23749 2486 28000 2488
rect 23749 2483 23815 2486
rect 27520 2456 28000 2486
rect 13721 2410 13787 2413
rect 19057 2410 19123 2413
rect 13721 2408 19123 2410
rect 13721 2352 13726 2408
rect 13782 2352 19062 2408
rect 19118 2352 19123 2408
rect 13721 2350 19123 2352
rect 13721 2347 13787 2350
rect 19057 2347 19123 2350
rect 21633 2410 21699 2413
rect 23841 2410 23907 2413
rect 21633 2408 23907 2410
rect 21633 2352 21638 2408
rect 21694 2352 23846 2408
rect 23902 2352 23907 2408
rect 21633 2350 23907 2352
rect 21633 2347 21699 2350
rect 23841 2347 23907 2350
rect 16757 2274 16823 2277
rect 16757 2272 20914 2274
rect 16757 2216 16762 2272
rect 16818 2216 20914 2272
rect 16757 2214 20914 2216
rect 16757 2211 16823 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 11605 2002 11671 2005
rect 20713 2002 20779 2005
rect 11605 2000 20779 2002
rect 11605 1944 11610 2000
rect 11666 1944 20718 2000
rect 20774 1944 20779 2000
rect 11605 1942 20779 1944
rect 20854 2002 20914 2214
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 27520 2002 28000 2032
rect 20854 1942 28000 2002
rect 11605 1939 11671 1942
rect 20713 1939 20779 1942
rect 27520 1912 28000 1942
rect 14457 1866 14523 1869
rect 22737 1866 22803 1869
rect 14457 1864 22803 1866
rect 14457 1808 14462 1864
rect 14518 1808 22742 1864
rect 22798 1808 22803 1864
rect 14457 1806 22803 1808
rect 14457 1803 14523 1806
rect 22737 1803 22803 1806
rect 10777 1730 10843 1733
rect 17309 1730 17375 1733
rect 10777 1728 17375 1730
rect 10777 1672 10782 1728
rect 10838 1672 17314 1728
rect 17370 1672 17375 1728
rect 10777 1670 17375 1672
rect 10777 1667 10843 1670
rect 17309 1667 17375 1670
rect 14825 1594 14891 1597
rect 23933 1594 23999 1597
rect 14825 1592 23999 1594
rect 14825 1536 14830 1592
rect 14886 1536 23938 1592
rect 23994 1536 23999 1592
rect 14825 1534 23999 1536
rect 14825 1531 14891 1534
rect 23933 1531 23999 1534
rect 5717 1458 5783 1461
rect 16113 1458 16179 1461
rect 5717 1456 16179 1458
rect 5717 1400 5722 1456
rect 5778 1400 16118 1456
rect 16174 1400 16179 1456
rect 5717 1398 16179 1400
rect 5717 1395 5783 1398
rect 16113 1395 16179 1398
rect 19057 1458 19123 1461
rect 27520 1458 28000 1488
rect 19057 1456 28000 1458
rect 19057 1400 19062 1456
rect 19118 1400 28000 1456
rect 19057 1398 28000 1400
rect 19057 1395 19123 1398
rect 27520 1368 28000 1398
rect 17125 914 17191 917
rect 27520 914 28000 944
rect 17125 912 28000 914
rect 17125 856 17130 912
rect 17186 856 28000 912
rect 17125 854 28000 856
rect 17125 851 17191 854
rect 27520 824 28000 854
rect 23565 370 23631 373
rect 27520 370 28000 400
rect 23565 368 28000 370
rect 23565 312 23570 368
rect 23626 312 28000 368
rect 23565 310 28000 312
rect 23565 307 23631 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 17172 17988 17236 18052
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 17356 14724 17420 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 14596 13696 14660 13700
rect 14596 13640 14646 13696
rect 14646 13640 14660 13696
rect 14596 13636 14660 13640
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 17172 12412 17236 12476
rect 17172 12200 17236 12204
rect 17172 12144 17186 12200
rect 17186 12144 17236 12200
rect 17172 12140 17236 12144
rect 17356 12004 17420 12068
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 14596 10916 14660 10980
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 17171 18052 17237 18053
rect 17171 17988 17172 18052
rect 17236 17988 17237 18052
rect 17171 17987 17237 17988
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14595 13700 14661 13701
rect 14595 13636 14596 13700
rect 14660 13636 14661 13700
rect 14595 13635 14661 13636
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 14598 10981 14658 13635
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 17174 12477 17234 17987
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 17355 14788 17421 14789
rect 17355 14724 17356 14788
rect 17420 14724 17421 14788
rect 17355 14723 17421 14724
rect 17171 12476 17237 12477
rect 17171 12412 17172 12476
rect 17236 12412 17237 12476
rect 17171 12411 17237 12412
rect 17174 12205 17234 12411
rect 17171 12204 17237 12205
rect 17171 12140 17172 12204
rect 17236 12140 17237 12204
rect 17171 12139 17237 12140
rect 17358 12069 17418 14723
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 17355 12068 17421 12069
rect 17355 12004 17356 12068
rect 17420 12004 17421 12068
rect 17355 12003 17421 12004
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14595 10980 14661 10981
rect 14595 10916 14596 10980
rect 14660 10916 14661 10980
rect 14595 10915 14661 10916
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _101_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_108
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12880 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1604681595
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1604681595
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15364 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_174
timestamp 1604681595
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_174
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_178
timestamp 1604681595
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1604681595
transform 1 0 20056 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_203
timestamp 1604681595
transform 1 0 19780 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp 1604681595
transform 1 0 20424 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_229
timestamp 1604681595
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1604681595
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1604681595
transform 1 0 22540 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604681595
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_237
timestamp 1604681595
transform 1 0 22908 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_239
timestamp 1604681595
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1604681595
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_243
timestamp 1604681595
transform 1 0 23460 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_255
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_251
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_255
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_267
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_263
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_267
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 24932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_275
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _038_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10120 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_97
timestamp 1604681595
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_101
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_113
timestamp 1604681595
transform 1 0 11500 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp 1604681595
transform 1 0 13064 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_142
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1604681595
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1604681595
transform 1 0 16192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_189
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1604681595
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21528 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21344 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1604681595
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_262
timestamp 1604681595
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_266
timestamp 1604681595
transform 1 0 25576 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1604681595
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1604681595
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1604681595
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1604681595
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18124 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1604681595
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_176
timestamp 1604681595
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_191
timestamp 1604681595
transform 1 0 18676 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_218
timestamp 1604681595
transform 1 0 21160 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_223
timestamp 1604681595
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1604681595
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1604681595
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_268
timestamp 1604681595
transform 1 0 25760 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1604681595
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_132
timestamp 1604681595
transform 1 0 13248 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1604681595
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16836 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1604681595
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 1604681595
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1604681595
transform 1 0 17756 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_196
timestamp 1604681595
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_200
timestamp 1604681595
transform 1 0 19504 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1604681595
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1604681595
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604681595
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1604681595
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_222
timestamp 1604681595
transform 1 0 21528 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23000 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22448 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_230
timestamp 1604681595
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_234
timestamp 1604681595
transform 1 0 22632 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_247
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24564 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_264
timestamp 1604681595
transform 1 0 25392 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_272
timestamp 1604681595
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_106
timestamp 1604681595
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1604681595
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_161
timestamp 1604681595
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1604681595
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18216 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19780 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_195
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1604681595
transform 1 0 20608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 1604681595
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_224
timestamp 1604681595
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_228
timestamp 1604681595
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23828 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_266
timestamp 1604681595
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_270
timestamp 1604681595
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_77
timestamp 1604681595
transform 1 0 8188 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_70
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1604681595
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1604681595
transform 1 0 9752 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1604681595
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 1604681595
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_107
timestamp 1604681595
transform 1 0 10948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1604681595
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_132
timestamp 1604681595
transform 1 0 13248 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1604681595
transform 1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13340 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1604681595
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1604681595
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1604681595
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_149
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_163
timestamp 1604681595
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1604681595
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15732 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_167
timestamp 1604681595
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_182
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18124 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18216 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 19688 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_205
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_194
timestamp 1604681595
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1604681595
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 1604681595
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1604681595
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1604681595
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20976 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1604681595
transform 1 0 22908 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_233
timestamp 1604681595
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_235
timestamp 1604681595
transform 1 0 22724 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_241
timestamp 1604681595
transform 1 0 23276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23276 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23460 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp 1604681595
transform 1 0 24012 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 25024 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24380 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24472 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_252
timestamp 1604681595
transform 1 0 24288 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_256
timestamp 1604681595
transform 1 0 24656 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_264
timestamp 1604681595
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_262
timestamp 1604681595
transform 1 0 25208 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_272
timestamp 1604681595
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_274
timestamp 1604681595
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_140
timestamp 1604681595
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1604681595
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_148
timestamp 1604681595
transform 1 0 14720 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18216 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17940 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1604681595
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20976 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23460 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_235
timestamp 1604681595
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 25024 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_252
timestamp 1604681595
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_256
timestamp 1604681595
transform 1 0 24656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_82
timestamp 1604681595
transform 1 0 8648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 14352 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_138
timestamp 1604681595
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_142
timestamp 1604681595
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_160
timestamp 1604681595
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_164
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_168
timestamp 1604681595
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1604681595
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1604681595
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_219
timestamp 1604681595
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_264
timestamp 1604681595
transform 1 0 25392 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604681595
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1604681595
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_132
timestamp 1604681595
transform 1 0 13248 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 17204 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_167
timestamp 1604681595
transform 1 0 16468 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_182
timestamp 1604681595
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 19780 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_195
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_199
timestamp 1604681595
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_206
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_224
timestamp 1604681595
transform 1 0 21712 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_229
timestamp 1604681595
transform 1 0 22172 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22540 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22356 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 25024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_252
timestamp 1604681595
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_256
timestamp 1604681595
transform 1 0 24656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12512 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14076 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1604681595
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_137
timestamp 1604681595
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1604681595
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_164
timestamp 1604681595
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18952 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21436 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1604681595
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1604681595
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23828 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_230
timestamp 1604681595
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_234
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_266
timestamp 1604681595
transform 1 0 25576 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_274
timestamp 1604681595
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1604681595
transform 1 0 10948 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_132
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15548 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_176
timestamp 1604681595
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_180
timestamp 1604681595
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1604681595
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1604681595
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20332 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23828 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22816 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_234
timestamp 1604681595
transform 1 0 22632 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_238
timestamp 1604681595
transform 1 0 23000 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_243
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_256
timestamp 1604681595
transform 1 0 24656 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_268
timestamp 1604681595
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1604681595
transform 1 0 10948 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_106
timestamp 1604681595
transform 1 0 10856 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11316 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_134
timestamp 1604681595
transform 1 0 13432 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_138
timestamp 1604681595
transform 1 0 13800 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604681595
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_140
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_145
timestamp 1604681595
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_149
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1604681595
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1604681595
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_170
timestamp 1604681595
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1604681595
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_171
timestamp 1604681595
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17204 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1604681595
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_207
timestamp 1604681595
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_188
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20516 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20516 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604681595
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604681595
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_224
timestamp 1604681595
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 22080 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_232
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_235
timestamp 1604681595
transform 1 0 22724 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_231
timestamp 1604681595
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22724 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 22908 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_244
timestamp 1604681595
transform 1 0 23552 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_240
timestamp 1604681595
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23828 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23920 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_256
timestamp 1604681595
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_260
timestamp 1604681595
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_267
timestamp 1604681595
transform 1 0 25668 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_267
timestamp 1604681595
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_275
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1604681595
transform 1 0 10488 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_138
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15732 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 1604681595
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_168
timestamp 1604681595
transform 1 0 16560 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_172
timestamp 1604681595
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 19964 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 19688 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1604681595
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_201
timestamp 1604681595
transform 1 0 19596 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20976 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1604681595
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1604681595
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_229
timestamp 1604681595
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23736 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_255
timestamp 1604681595
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_259
timestamp 1604681595
transform 1 0 24932 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_270
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_107
timestamp 1604681595
transform 1 0 10948 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_115
timestamp 1604681595
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_119
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_150
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_169
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_192
timestamp 1604681595
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_196
timestamp 1604681595
transform 1 0 19136 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1604681595
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_228
timestamp 1604681595
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22816 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_232
timestamp 1604681595
transform 1 0 22448 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_255
timestamp 1604681595
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_259
timestamp 1604681595
transform 1 0 24932 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1604681595
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1604681595
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1604681595
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp 1604681595
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_133
timestamp 1604681595
transform 1 0 13340 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1604681595
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1604681595
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_165
timestamp 1604681595
transform 1 0 16284 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1604681595
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_207
timestamp 1604681595
transform 1 0 20148 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1604681595
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1604681595
transform 1 0 24012 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24288 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_261
timestamp 1604681595
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1604681595
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11500 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_136
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_139
timestamp 1604681595
transform 1 0 13892 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_171
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1604681595
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1604681595
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_209
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23552 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23184 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_234
timestamp 1604681595
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1604681595
transform 1 0 23000 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_242
timestamp 1604681595
transform 1 0 23368 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_94
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_97
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1604681595
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_124
timestamp 1604681595
transform 1 0 12512 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_133
timestamp 1604681595
transform 1 0 13340 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp 1604681595
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13708 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1604681595
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_159
timestamp 1604681595
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16008 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17848 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18216 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_173
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_195
timestamp 1604681595
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_191
timestamp 1604681595
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_195
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1604681595
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19780 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604681595
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_226
timestamp 1604681595
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_229
timestamp 1604681595
transform 1 0 22172 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_241
timestamp 1604681595
transform 1 0 23276 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_245
timestamp 1604681595
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 24104 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 25024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_258
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_262
timestamp 1604681595
transform 1 0 25208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_266
timestamp 1604681595
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1604681595
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1604681595
transform 1 0 9752 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12788 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_140
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16100 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 16928 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_211
timestamp 1604681595
transform 1 0 20516 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 24104 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_273
timestamp 1604681595
transform 1 0 26220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_100
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_123
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_127
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15548 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 17112 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16744 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_172
timestamp 1604681595
transform 1 0 16928 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_193
timestamp 1604681595
transform 1 0 18860 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_199
timestamp 1604681595
transform 1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_224
timestamp 1604681595
transform 1 0 21712 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_229
timestamp 1604681595
transform 1 0 22172 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 22540 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22356 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 25024 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24472 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_252
timestamp 1604681595
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_256
timestamp 1604681595
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_264
timestamp 1604681595
transform 1 0 25392 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_272
timestamp 1604681595
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_94
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15364 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_146
timestamp 1604681595
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_150
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18216 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_174
timestamp 1604681595
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_178
timestamp 1604681595
transform 1 0 17480 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19780 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1604681595
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_199
timestamp 1604681595
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_226
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1604681595
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_270
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_274
timestamp 1604681595
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 10304 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_99
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1604681595
transform 1 0 10580 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_107
timestamp 1604681595
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1604681595
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_134
timestamp 1604681595
transform 1 0 13432 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1604681595
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_162
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16744 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_179
timestamp 1604681595
transform 1 0 17572 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18952 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1604681595
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1604681595
transform 1 0 18768 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_196
timestamp 1604681595
transform 1 0 19136 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_224
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_228
timestamp 1604681595
transform 1 0 22080 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 22540 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22356 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24472 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_252
timestamp 1604681595
transform 1 0 24288 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_256
timestamp 1604681595
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_266
timestamp 1604681595
transform 1 0 25576 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604681595
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_94
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1604681595
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_165
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20056 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_197
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_202
timestamp 1604681595
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1604681595
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_219
timestamp 1604681595
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_268
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_272
timestamp 1604681595
transform 1 0 26128 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_82
timestamp 1604681595
transform 1 0 8648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_89
timestamp 1604681595
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_100
timestamp 1604681595
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10672 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1604681595
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11408 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_133
timestamp 1604681595
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_131
timestamp 1604681595
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_138
timestamp 1604681595
transform 1 0 13800 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_135
timestamp 1604681595
transform 1 0 13524 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_150
timestamp 1604681595
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_158
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_176
timestamp 1604681595
transform 1 0 17296 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1604681595
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1604681595
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1604681595
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1604681595
transform 1 0 17664 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_197
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18400 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1604681595
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_205
timestamp 1604681595
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_201
timestamp 1604681595
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20148 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20148 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604681595
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1604681595
transform 1 0 20332 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20516 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_226
timestamp 1604681595
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1604681595
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_234
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_230
timestamp 1604681595
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22448 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_247
timestamp 1604681595
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1604681595
transform 1 0 23276 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_258
timestamp 1604681595
transform 1 0 24840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_262
timestamp 1604681595
transform 1 0 25208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1604681595
transform 1 0 25576 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1604681595
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_268
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604681595
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604681595
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_89
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_106
timestamp 1604681595
transform 1 0 10856 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_112
timestamp 1604681595
transform 1 0 11408 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_115
timestamp 1604681595
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1604681595
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14904 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 17756 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1604681595
transform 1 0 17020 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_177
timestamp 1604681595
transform 1 0 17388 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_200
timestamp 1604681595
transform 1 0 19504 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_205
timestamp 1604681595
transform 1 0 19964 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1604681595
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23920 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_234
timestamp 1604681595
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_238
timestamp 1604681595
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_242
timestamp 1604681595
transform 1 0 23368 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_247
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_257
timestamp 1604681595
transform 1 0 24748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_261
timestamp 1604681595
transform 1 0 25116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1604681595
transform 1 0 25484 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 1604681595
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8740 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_80
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_102
timestamp 1604681595
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1604681595
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1604681595
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_145
timestamp 1604681595
transform 1 0 14444 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_163
timestamp 1604681595
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18308 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1604681595
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_177
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_206
timestamp 1604681595
transform 1 0 20056 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_211
timestamp 1604681595
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1604681595
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_223
timestamp 1604681595
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1604681595
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_268
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_74
timestamp 1604681595
transform 1 0 7912 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1604681595
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_81
timestamp 1604681595
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1604681595
transform 1 0 8924 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1604681595
transform 1 0 9292 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11776 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_107
timestamp 1604681595
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_111
timestamp 1604681595
transform 1 0 11316 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 14260 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1604681595
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_146
timestamp 1604681595
transform 1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1604681595
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_157
timestamp 1604681595
transform 1 0 15548 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_162
timestamp 1604681595
transform 1 0 16008 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16192 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16468 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1604681595
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1604681595
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19228 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_193
timestamp 1604681595
transform 1 0 18860 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1604681595
transform 1 0 19412 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 21068 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_225
timestamp 1604681595
transform 1 0 21804 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1604681595
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21620 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22172 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_248
timestamp 1604681595
transform 1 0 23920 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24472 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_252
timestamp 1604681595
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1604681595
transform 1 0 25484 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_273
timestamp 1604681595
transform 1 0 26220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1604681595
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1604681595
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_102
timestamp 1604681595
transform 1 0 10488 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12604 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_31_150
timestamp 1604681595
transform 1 0 14904 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1604681595
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1604681595
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1604681595
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19688 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1604681595
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21252 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1604681595
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_228
timestamp 1604681595
transform 1 0 22080 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_233
timestamp 1604681595
transform 1 0 22540 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1604681595
transform 1 0 22908 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1604681595
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_268
timestamp 1604681595
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_272
timestamp 1604681595
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_276
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_77
timestamp 1604681595
transform 1 0 8188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12144 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_112
timestamp 1604681595
transform 1 0 11408 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_131
timestamp 1604681595
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_135
timestamp 1604681595
transform 1 0 13524 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_142
timestamp 1604681595
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15824 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_146
timestamp 1604681595
transform 1 0 14536 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 18308 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1604681595
transform 1 0 17572 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1604681595
transform 1 0 17940 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_186
timestamp 1604681595
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21620 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_210
timestamp 1604681595
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1604681595
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_225
timestamp 1604681595
transform 1 0 21804 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_229
timestamp 1604681595
transform 1 0 22172 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22356 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23920 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_240
timestamp 1604681595
transform 1 0 23184 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_244
timestamp 1604681595
transform 1 0 23552 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_247
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_257
timestamp 1604681595
transform 1 0 24748 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_261
timestamp 1604681595
transform 1 0 25116 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1604681595
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7544 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_72
timestamp 1604681595
transform 1 0 7728 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_89
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_97
timestamp 1604681595
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_34_116
timestamp 1604681595
transform 1 0 11776 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12328 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12512 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_133
timestamp 1604681595
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1604681595
transform 1 0 13340 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_137
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13892 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_158
timestamp 1604681595
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_162
timestamp 1604681595
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_147
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1604681595
transform 1 0 17020 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_177
timestamp 1604681595
transform 1 0 17388 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17572 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1604681595
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_194
timestamp 1604681595
transform 1 0 18952 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_190
timestamp 1604681595
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 19136 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_206
timestamp 1604681595
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_201
timestamp 1604681595
transform 1 0 19596 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 19320 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19504 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_34_210
timestamp 1604681595
transform 1 0 20424 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_223
timestamp 1604681595
transform 1 0 21620 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_219
timestamp 1604681595
transform 1 0 21252 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_223
timestamp 1604681595
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_219
timestamp 1604681595
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 21804 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 21436 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21804 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23920 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_246
timestamp 1604681595
transform 1 0 23736 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_250
timestamp 1604681595
transform 1 0 24104 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24472 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_264
timestamp 1604681595
transform 1 0 25392 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_260
timestamp 1604681595
transform 1 0 25024 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_272
timestamp 1604681595
transform 1 0 26128 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_97
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_101
timestamp 1604681595
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604681595
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14444 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_126
timestamp 1604681595
transform 1 0 12696 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_141
timestamp 1604681595
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_154
timestamp 1604681595
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_158
timestamp 1604681595
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_171
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1604681595
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1604681595
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1604681595
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_201
timestamp 1604681595
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1604681595
transform 1 0 19964 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_234
timestamp 1604681595
transform 1 0 22632 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_238
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24104 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 25576 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24288 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_258
timestamp 1604681595
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1604681595
transform 1 0 25208 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_90
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11040 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_107
timestamp 1604681595
transform 1 0 10948 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13524 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13340 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_127
timestamp 1604681595
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_131
timestamp 1604681595
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_144
timestamp 1604681595
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_148
timestamp 1604681595
transform 1 0 14720 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_160
timestamp 1604681595
transform 1 0 15824 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_164
timestamp 1604681595
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 16560 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17572 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_171
timestamp 1604681595
transform 1 0 16836 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_175
timestamp 1604681595
transform 1 0 17204 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19136 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18768 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_188
timestamp 1604681595
transform 1 0 18400 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1604681595
transform 1 0 18952 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 21252 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_210
timestamp 1604681595
transform 1 0 20424 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1604681595
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1604681595
transform 1 0 21620 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_229
timestamp 1604681595
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 22356 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_36_240
timestamp 1604681595
transform 1 0 23184 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 24564 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_252
timestamp 1604681595
transform 1 0 24288 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_259
timestamp 1604681595
transform 1 0 24932 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1604681595
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_106
timestamp 1604681595
transform 1 0 10856 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_111
timestamp 1604681595
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_115
timestamp 1604681595
transform 1 0 11684 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1604681595
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13340 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_129
timestamp 1604681595
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_152
timestamp 1604681595
transform 1 0 15088 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1604681595
transform 1 0 15456 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_162
timestamp 1604681595
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18768 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18584 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_188
timestamp 1604681595
transform 1 0 18400 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 21896 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_211
timestamp 1604681595
transform 1 0 20516 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_217
timestamp 1604681595
transform 1 0 21068 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_224
timestamp 1604681595
transform 1 0 21712 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_228
timestamp 1604681595
transform 1 0 22080 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23736 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1604681595
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 25024 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_252
timestamp 1604681595
transform 1 0 24288 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_256
timestamp 1604681595
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1604681595
transform 1 0 25392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_268
timestamp 1604681595
transform 1 0 25760 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604681595
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11132 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_107
timestamp 1604681595
transform 1 0 10948 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_128
timestamp 1604681595
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_132
timestamp 1604681595
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1604681595
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_149
timestamp 1604681595
transform 1 0 14812 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14904 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_162
timestamp 1604681595
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_158
timestamp 1604681595
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16100 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_182
timestamp 1604681595
transform 1 0 17848 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1604681595
transform 1 0 18216 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19596 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_199
timestamp 1604681595
transform 1 0 19412 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_203
timestamp 1604681595
transform 1 0 19780 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1604681595
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_219
timestamp 1604681595
transform 1 0 21252 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22816 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24104 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23736 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_231
timestamp 1604681595
transform 1 0 22356 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_235
timestamp 1604681595
transform 1 0 22724 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_242
timestamp 1604681595
transform 1 0 23368 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_248
timestamp 1604681595
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 25392 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_256
timestamp 1604681595
transform 1 0 24656 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_267
timestamp 1604681595
transform 1 0 25668 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_102
timestamp 1604681595
transform 1 0 10488 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_125
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_119
timestamp 1604681595
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_107
timestamp 1604681595
transform 1 0 10948 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_39_142
timestamp 1604681595
transform 1 0 14168 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_136
timestamp 1604681595
transform 1 0 13616 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15364 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_148
timestamp 1604681595
transform 1 0 14720 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1604681595
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_164
timestamp 1604681595
transform 1 0 16192 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_176
timestamp 1604681595
transform 1 0 17296 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_174
timestamp 1604681595
transform 1 0 17112 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1604681595
transform 1 0 16652 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604681595
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 16928 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 18032 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 19228 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_203
timestamp 1604681595
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_207
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1604681595
transform 1 0 18400 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_196
timestamp 1604681595
transform 1 0 19136 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1604681595
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1604681595
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_215
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_220
timestamp 1604681595
transform 1 0 21344 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_218
timestamp 1604681595
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 20976 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_226
timestamp 1604681595
transform 1 0 21896 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_229
timestamp 1604681595
transform 1 0 22172 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_235
timestamp 1604681595
transform 1 0 22724 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23736 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_247
timestamp 1604681595
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 25024 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_252
timestamp 1604681595
transform 1 0 24288 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1604681595
transform 1 0 25392 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_268
timestamp 1604681595
transform 1 0 25760 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_259
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_276
timestamp 1604681595
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1604681595
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 12512 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 13616 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604681595
transform 1 0 13064 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_128
timestamp 1604681595
transform 1 0 12880 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_140
timestamp 1604681595
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 15824 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 14720 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604681595
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604681595
transform 1 0 15272 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_152
timestamp 1604681595
transform 1 0 15088 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_156
timestamp 1604681595
transform 1 0 15456 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_164
timestamp 1604681595
transform 1 0 16192 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 16928 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604681595
transform 1 0 16744 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_168
timestamp 1604681595
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_175
timestamp 1604681595
transform 1 0 17204 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 19504 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 20056 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_188
timestamp 1604681595
transform 1 0 18400 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_192
timestamp 1604681595
transform 1 0 18768 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_195
timestamp 1604681595
transform 1 0 19044 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_204
timestamp 1604681595
transform 1 0 19872 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 20884 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 21988 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 21712 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 20700 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_212
timestamp 1604681595
transform 1 0 20608 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_219
timestamp 1604681595
transform 1 0 21252 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1604681595
transform 1 0 21620 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_226
timestamp 1604681595
transform 1 0 21896 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_231
timestamp 1604681595
transform 1 0 22356 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_235
timestamp 1604681595
transform 1 0 22724 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_238
timestamp 1604681595
transform 1 0 23000 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_259
timestamp 1604681595
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_275
timestamp 1604681595
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 16192 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 18860 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1604681595
transform 1 0 19228 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 21712 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1604681595
transform 1 0 20332 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_228
timestamp 1604681595
transform 1 0 22080 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 22816 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_240
timestamp 1604681595
transform 1 0 23184 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 6944 480 7064 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 20952 480 21072 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27520 23672 28000 23792 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26882 0 26938 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 938 27520 994 28000 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 7746 27520 7802 28000 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 9126 27520 9182 28000 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1582 27520 1638 28000 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2962 27520 3018 28000 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4986 27520 5042 28000 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 5722 27520 5778 28000 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 23478 27520 23534 28000 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 25502 27520 25558 28000 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 26146 27520 26202 28000 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 26882 27520 26938 28000 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 27526 27520 27582 28000 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 15290 27520 15346 28000 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 17314 27520 17370 28000 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 20718 27520 20774 28000 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 prog_clk
port 123 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 124 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 125 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 126 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 127 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_bottom_grid_pin_38_
port 128 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 129 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 130 nsew default input
rlabel metal3 s 27520 4224 28000 4344 6 right_bottom_grid_pin_41_
port 131 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
