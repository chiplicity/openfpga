* NGSPICE file created from sb_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

.subckt sb_0__1_ bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk right_top_grid_pin_42_ right_top_grid_pin_43_ right_top_grid_pin_44_
+ right_top_grid_pin_45_ right_top_grid_pin_46_ right_top_grid_pin_47_ right_top_grid_pin_48_
+ right_top_grid_pin_49_ top_left_grid_pin_1_ vpwr vgnd
XFILLER_22_133 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_25.scs8hd_buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X _083_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_9_115 vpwr vgnd scs8hd_fill_2
XFILLER_9_148 vpwr vgnd scs8hd_fill_2
XFILLER_13_144 vgnd vpwr scs8hd_fill_1
XFILLER_13_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_18.mux_l1_in_0__S mux_right_track_18.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_181 vgnd vpwr scs8hd_decap_6
XFILLER_27_214 vgnd vpwr scs8hd_fill_1
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_236 vgnd vpwr scs8hd_decap_8
XFILLER_18_247 vpwr vgnd scs8hd_fill_2
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_18.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_16.mux_l2_in_0_/S mux_right_track_18.mux_l1_in_1_/S
+ mem_right_track_18.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_217 vpwr vgnd scs8hd_fill_2
X_062_ _062_/A chanx_right_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_23_86 vgnd vpwr scs8hd_decap_12
XFILLER_2_165 vgnd vpwr scs8hd_fill_1
XFILLER_2_132 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_231 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_2__A1 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
X_114_ _114_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
X_045_ _045_/HI _045_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__S mux_bottom_track_25.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_238 vpwr vgnd scs8hd_fill_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
X_028_ _028_/HI _028_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_161 vpwr vgnd scs8hd_fill_2
XFILLER_19_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 mux_right_track_2.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_33.scs8hd_buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X _079_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_15_98 vgnd vpwr scs8hd_decap_6
XFILLER_31_86 vgnd vpwr scs8hd_decap_3
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_31_112 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vpwr vgnd scs8hd_fill_2
XFILLER_22_145 vgnd vpwr scs8hd_decap_6
Xmem_right_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_127 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_215 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D mux_top_track_8.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_126 vpwr vgnd scs8hd_fill_2
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_33_207 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XFILLER_18_259 vgnd vpwr scs8hd_decap_12
XFILLER_17_270 vgnd vpwr scs8hd_decap_6
XFILLER_24_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_23_240 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__D mux_right_track_18.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
X_061_ chany_bottom_in[11] chanx_right_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_23_98 vgnd vpwr scs8hd_decap_12
XFILLER_14_262 vpwr vgnd scs8hd_fill_2
XFILLER_20_243 vpwr vgnd scs8hd_fill_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
X_113_ _113_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
X_044_ _044_/HI _044_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l3_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D mux_top_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_86 vgnd vpwr scs8hd_decap_8
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_132 vpwr vgnd scs8hd_fill_2
XFILLER_34_143 vgnd vpwr scs8hd_decap_4
XFILLER_1_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D mux_bottom_track_25.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_143 vpwr vgnd scs8hd_fill_2
XFILLER_15_22 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D mux_bottom_track_5.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_132 vpwr vgnd scs8hd_fill_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_224 vpwr vgnd scs8hd_fill_2
XFILLER_39_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1__A0 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_1_/S
+ mem_right_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.scs8hd_buf_4_0__A mux_right_track_12.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XFILLER_12_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_20.mux_l2_in_0__S mux_right_track_20.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_227 vpwr vgnd scs8hd_fill_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_149 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_3__A0 _033_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0__A1 mux_right_track_10.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_5_164 vgnd vpwr scs8hd_decap_4
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0__A0 mux_right_track_6.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0__S mux_right_track_14.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l3_in_0_ mux_right_track_10.mux_l2_in_1_/X mux_right_track_10.mux_l2_in_0_/X
+ mux_right_track_10.mux_l3_in_0_/S mux_right_track_10.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_263 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
X_060_ chany_bottom_in[7] chanx_right_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_3
XFILLER_0_26 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__061__A chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
X_112_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_043_ _043_/HI _043_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_10.mux_l2_in_1_ _051_/HI chany_bottom_in[9] mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l2_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_163 vpwr vgnd scs8hd_fill_2
XFILLER_1_91 vpwr vgnd scs8hd_fill_2
XFILLER_4_207 vgnd vpwr scs8hd_decap_4
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_26.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_26.mux_l1_in_0_/S mux_right_track_26.mux_l2_in_0_/S
+ mem_right_track_26.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_34_188 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D mux_right_track_0.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_158 vpwr vgnd scs8hd_fill_2
XFILLER_25_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2__S mux_bottom_track_9.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_34 vgnd vpwr scs8hd_decap_12
XFILLER_40_169 vgnd vpwr scs8hd_decap_6
XFILLER_0_232 vpwr vgnd scs8hd_fill_2
XFILLER_31_169 vgnd vpwr scs8hd_decap_3
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l3_in_0__S mux_right_track_12.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_158 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l1_in_1__A1 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ mem_right_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XFILLER_21_180 vgnd vpwr scs8hd_fill_1
XFILLER_36_206 vgnd vpwr scs8hd_fill_1
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_140 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.scs8hd_buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _093_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_27_239 vgnd vpwr scs8hd_decap_3
XFILLER_27_217 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.scs8hd_buf_4_0_ mux_right_track_12.mux_l3_in_0_/X _069_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__064__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XFILLER_37_98 vgnd vpwr scs8hd_decap_6
XFILLER_26_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.mux_l1_in_0__S mux_right_track_6.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l2_in_0__A1 mux_right_track_6.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_209 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 mux_top_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XANTENNA__059__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0__A0 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_2_135 vgnd vpwr scs8hd_fill_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D mux_right_track_2.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_201 vgnd vpwr scs8hd_fill_1
XFILLER_11_223 vpwr vgnd scs8hd_fill_2
X_111_ _111_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 bottom_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_11_234 vpwr vgnd scs8hd_fill_2
XFILLER_11_245 vgnd vpwr scs8hd_decap_3
X_042_ _042_/HI _042_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_10.mux_l2_in_0_ right_top_grid_pin_43_ mux_right_track_10.mux_l1_in_0_/X
+ mux_right_track_10.mux_l2_in_0_/S mux_right_track_10.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D mux_top_track_16.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_3.mux_l1_in_1_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_142 vpwr vgnd scs8hd_fill_2
XFILLER_37_197 vpwr vgnd scs8hd_fill_2
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__072__A _072_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XFILLER_28_197 vgnd vpwr scs8hd_decap_6
XFILLER_3_241 vgnd vpwr scs8hd_fill_1
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
Xmem_right_track_26.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_24.mux_l3_in_0_/S mux_right_track_26.mux_l1_in_0_/S
+ mem_right_track_26.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_34_167 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__D mux_right_track_20.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 _048_/HI vgnd vpwr scs8hd_diode_2
XFILLER_40_126 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_156 vpwr vgnd scs8hd_fill_2
XFILLER_15_46 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_1__A0 _052_/HI vgnd vpwr scs8hd_diode_2
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
XFILLER_0_222 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_3__S mux_right_track_6.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_1_ _035_/HI chany_bottom_in[8] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_145 vpwr vgnd scs8hd_fill_2
XFILLER_16_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_20.scs8hd_buf_4_0_ mux_right_track_20.mux_l2_in_0_/X _065_/A vgnd
+ vpwr scs8hd_buf_1
Xmux_top_track_0.mux_l2_in_1_ _036_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_192 vpwr vgnd scs8hd_fill_2
XFILLER_30_170 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_38_270 vgnd vpwr scs8hd_decap_4
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l3_in_0__A0 mux_right_track_12.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D mux_right_track_2.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_22.mux_l1_in_0__A0 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XANTENNA__080__A chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_41_243 vgnd vpwr scs8hd_fill_1
XFILLER_41_221 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_2_ chany_bottom_in[12] chany_bottom_in[2] mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_133 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.scs8hd_buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _114_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_232 vgnd vpwr scs8hd_fill_1
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_2_158 vgnd vpwr scs8hd_decap_4
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_22.mux_l1_in_1__S mux_right_track_22.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__D mux_right_track_20.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_224 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l1_in_0__S mux_right_track_10.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
X_110_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
X_041_ _041_/HI _041_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_24.mux_l2_in_1__S mux_top_track_24.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_132 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_264 vgnd vpwr scs8hd_decap_12
XFILLER_3_220 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XFILLER_19_165 vpwr vgnd scs8hd_fill_2
XFILLER_42_190 vgnd vpwr scs8hd_decap_8
XFILLER_19_176 vgnd vpwr scs8hd_decap_4
XFILLER_19_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 mux_bottom_track_5.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_149 vgnd vpwr scs8hd_fill_1
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_1__A1 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_ chany_top_in[11] chany_top_in[9] mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_8.mux_l2_in_0_ right_top_grid_pin_42_ mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_138 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 _035_/HI vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_249 vgnd vpwr scs8hd_decap_4
Xmux_right_track_22.mux_l2_in_0_ mux_right_track_22.mux_l1_in_1_/X mux_right_track_22.mux_l1_in_0_/X
+ mux_right_track_22.mux_l2_in_0_/S mux_right_track_22.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_105 vgnd vpwr scs8hd_decap_12
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XANTENNA__078__A chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_164 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l3_in_0__A1 mux_right_track_12.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_22.mux_l1_in_0__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_233 vpwr vgnd scs8hd_fill_2
XFILLER_26_252 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_ chanx_right_in[15] chanx_right_in[8] mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_22.mux_l1_in_1_ _030_/HI chany_bottom_in[17] mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_17_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_1__S mux_right_track_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_2_104 vgnd vpwr scs8hd_decap_8
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_20.scs8hd_buf_4_0__A mux_right_track_20.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_247 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__D mux_right_track_6.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_040_ _040_/HI _040_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_6_240 vgnd vpwr scs8hd_decap_3
XFILLER_6_273 vpwr vgnd scs8hd_fill_2
XFILLER_37_111 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1__S mux_top_track_8.mux_l1_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_136 vpwr vgnd scs8hd_fill_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D mux_right_track_24.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_228 vgnd vpwr scs8hd_decap_4
XFILLER_39_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 _041_/HI vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_117 vgnd vpwr scs8hd_decap_12
XFILLER_38_250 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A0 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 _054_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_21_172 vpwr vgnd scs8hd_fill_2
XFILLER_36_209 vgnd vpwr scs8hd_decap_3
XFILLER_8_154 vgnd vpwr scs8hd_fill_1
XFILLER_12_194 vgnd vpwr scs8hd_decap_6
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_3__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_198 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A mux_bottom_track_17.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D mux_right_track_8.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_264 vgnd vpwr scs8hd_decap_8
XFILLER_26_242 vgnd vpwr scs8hd_fill_1
XANTENNA__089__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_41_201 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_ chanx_right_in[1] top_left_grid_pin_1_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_1__S mux_right_track_6.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_22.mux_l1_in_0_ right_top_grid_pin_49_ chany_top_in[17] mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_5_168 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_32_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 mux_bottom_track_9.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_223 vgnd vpwr scs8hd_decap_3
XFILLER_23_245 vgnd vpwr scs8hd_decap_8
XFILLER_2_116 vgnd vpwr scs8hd_decap_8
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.scs8hd_buf_4_0__A mux_right_track_6.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_201 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_25.mux_l2_in_1_ _045_/HI chanx_right_in[14] mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S mux_bottom_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__D mux_right_track_26.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_219 vpwr vgnd scs8hd_fill_2
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
X_099_ _099_/A chany_top_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_167 vgnd vpwr scs8hd_decap_4
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__097__A chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_28_167 vpwr vgnd scs8hd_fill_2
XFILLER_3_233 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_1_ _049_/HI mux_bottom_track_9.mux_l1_in_2_/X mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_19_123 vgnd vpwr scs8hd_decap_6
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XFILLER_42_181 vgnd vpwr scs8hd_decap_3
XFILLER_33_170 vpwr vgnd scs8hd_fill_2
XFILLER_25_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_115 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 mux_top_track_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_129 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[16] mux_bottom_track_9.mux_l1_in_1_/S
+ mux_bottom_track_9.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_144 vgnd vpwr scs8hd_decap_6
XFILLER_12_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_41_213 vgnd vpwr scs8hd_decap_4
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A mux_bottom_track_5.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 mux_top_track_16.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_114 vgnd vpwr scs8hd_decap_4
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_254 vpwr vgnd scs8hd_fill_2
XFILLER_17_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_4.scs8hd_buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _073_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_2_128 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
XFILLER_14_235 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S mux_bottom_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l2_in_1__S mux_right_track_10.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_227 vpwr vgnd scs8hd_fill_2
XFILLER_11_238 vgnd vpwr scs8hd_decap_4
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_098_ chany_bottom_in[16] chany_top_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_37_179 vpwr vgnd scs8hd_fill_2
XFILLER_37_146 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_135 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_25.mux_l1_in_1_ chanx_right_in[7] chanx_right_in[0] mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_0_/S mux_bottom_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_149 vpwr vgnd scs8hd_fill_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_8
XFILLER_42_160 vpwr vgnd scs8hd_fill_2
XFILLER_25_138 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_16.mux_l1_in_1_/S mux_right_track_16.mux_l2_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XFILLER_0_215 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_16_105 vgnd vpwr scs8hd_decap_8
XFILLER_16_149 vpwr vgnd scs8hd_fill_2
XFILLER_31_108 vpwr vgnd scs8hd_fill_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_30_130 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vgnd vpwr scs8hd_fill_1
XFILLER_15_182 vgnd vpwr scs8hd_fill_1
XFILLER_30_196 vpwr vgnd scs8hd_fill_2
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_1_ chanx_right_in[9] chanx_right_in[2] mux_bottom_track_9.mux_l1_in_1_/S
+ mux_bottom_track_9.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1__A0 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_225 vpwr vgnd scs8hd_fill_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D mux_bottom_track_9.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.scs8hd_buf_4_0__A mux_top_track_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_18.scs8hd_buf_4_0_ mux_right_track_18.mux_l2_in_0_/X _066_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_4_181 vgnd vpwr scs8hd_decap_3
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S mux_top_track_16.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 mux_top_track_8.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_184 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_6
XFILLER_20_228 vgnd vpwr scs8hd_fill_1
XFILLER_6_210 vpwr vgnd scs8hd_fill_2
XFILLER_10_261 vgnd vpwr scs8hd_decap_12
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
X_097_ chany_bottom_in[17] chany_top_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_6_254 vpwr vgnd scs8hd_fill_2
XFILLER_6_265 vgnd vpwr scs8hd_decap_8
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_86 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_1_ _037_/HI chany_bottom_in[17] mux_top_track_16.mux_l2_in_1_/S
+ mux_top_track_16.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D mux_top_track_24.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A0 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_25_106 vgnd vpwr scs8hd_decap_3
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_14.mux_l3_in_0_/S mux_right_track_16.mux_l1_in_1_/S
+ mem_right_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_128 vpwr vgnd scs8hd_fill_2
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_30_164 vgnd vpwr scs8hd_decap_6
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_150 vpwr vgnd scs8hd_fill_2
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_1_/S
+ mux_bottom_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_197 vpwr vgnd scs8hd_fill_2
Xmux_right_track_26.scs8hd_buf_4_0_ mux_right_track_26.mux_l2_in_0_/X _062_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_29_231 vpwr vgnd scs8hd_fill_2
XFILLER_29_220 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1__A1 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l3_in_0__S mux_top_track_32.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_3
XFILLER_35_223 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_41_237 vgnd vpwr scs8hd_decap_6
XFILLER_26_256 vgnd vpwr scs8hd_decap_4
XFILLER_26_234 vpwr vgnd scs8hd_fill_2
XFILLER_32_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D mux_top_track_0.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_234 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.scs8hd_buf_4_0_ mux_top_track_8.mux_l3_in_0_/X _111_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_130 vpwr vgnd scs8hd_fill_2
XFILLER_1_174 vgnd vpwr scs8hd_decap_3
XANTENNA__100__A chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__D mux_right_track_8.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A mux_bottom_track_25.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_273 vpwr vgnd scs8hd_fill_2
X_096_ chany_bottom_in[18] chany_top_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_159 vpwr vgnd scs8hd_fill_2
XFILLER_37_104 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S mux_top_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XFILLER_36_181 vgnd vpwr scs8hd_decap_6
XFILLER_42_173 vgnd vpwr scs8hd_decap_8
X_079_ _079_/A chany_bottom_out[16] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A1 mux_top_track_32.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_18_181 vpwr vgnd scs8hd_fill_2
XFILLER_18_192 vgnd vpwr scs8hd_decap_3
XFILLER_33_140 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_228 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_3_ _033_/HI chany_bottom_in[5] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_1_ chany_bottom_in[8] chanx_right_in[19] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D mux_top_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_154 vgnd vpwr scs8hd_fill_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vgnd vpwr scs8hd_decap_12
XFILLER_21_132 vgnd vpwr scs8hd_decap_8
XFILLER_21_176 vgnd vpwr scs8hd_decap_4
XFILLER_29_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_213 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l3_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_8.scs8hd_buf_4_0__A mux_top_track_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_191 vpwr vgnd scs8hd_fill_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_202 vgnd vpwr scs8hd_fill_1
XFILLER_5_106 vgnd vpwr scs8hd_decap_3
XFILLER_32_238 vgnd vpwr scs8hd_decap_8
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
Xmem_right_track_24.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l3_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l3_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XFILLER_1_142 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_0.mux_l1_in_2_/S mux_right_track_0.mux_l2_in_1_/S
+ mem_right_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_10.scs8hd_buf_4_0__A mux_right_track_10.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
X_095_ _095_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_230 vgnd vpwr scs8hd_fill_1
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__S mux_bottom_track_17.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_237 vgnd vpwr scs8hd_decap_4
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
XANTENNA__106__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
X_078_ chany_top_in[16] chany_bottom_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_174 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_218 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_2_ right_top_grid_pin_48_ right_top_grid_pin_46_ mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_2__D mux_right_track_12.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_141 vgnd vpwr scs8hd_fill_1
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[5] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_122 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_174 vpwr vgnd scs8hd_fill_2
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l3_in_0__S mux_top_track_8.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_21_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_266 vpwr vgnd scs8hd_fill_2
XFILLER_12_133 vgnd vpwr scs8hd_decap_8
XFILLER_12_144 vgnd vpwr scs8hd_decap_3
XFILLER_12_177 vpwr vgnd scs8hd_fill_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_35_236 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_1.mux_l1_in_1_/S mux_bottom_track_1.mux_l2_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_118 vgnd vpwr scs8hd_fill_1
XFILLER_17_203 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_258 vgnd vpwr scs8hd_decap_12
Xmem_right_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_24.mux_l1_in_0_/S mux_right_track_24.mux_l2_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D mux_top_track_4.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_4.mux_l1_in_0_/S mux_top_track_4.mux_l2_in_1_/S
+ mem_top_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_261 vpwr vgnd scs8hd_fill_2
XFILLER_23_228 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_20.mux_l1_in_0__S mux_right_track_20.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_228 vgnd vpwr scs8hd_decap_4
XFILLER_14_239 vgnd vpwr scs8hd_decap_4
XFILLER_13_86 vgnd vpwr scs8hd_decap_6
XFILLER_1_165 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_265 vgnd vpwr scs8hd_decap_12
XFILLER_34_19 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_32.mux_l3_in_0_/S mux_right_track_0.mux_l1_in_2_/S
+ mem_right_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__D mux_right_track_14.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
X_094_ _094_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_128 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.scs8hd_buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _095_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_164 vgnd vpwr scs8hd_decap_4
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_077_ chany_top_in[17] chany_bottom_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_ _054_/HI chany_bottom_in[13] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_4.mux_l1_in_1_ right_top_grid_pin_44_ right_top_grid_pin_42_ mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_197 vgnd vpwr scs8hd_decap_4
XFILLER_21_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_30_101 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0__A0 chany_top_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_30_145 vpwr vgnd scs8hd_fill_2
XFILLER_30_134 vpwr vgnd scs8hd_fill_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_123 vgnd vpwr scs8hd_decap_6
XFILLER_21_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D mux_bottom_track_3.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_9.mux_l2_in_0_/S mux_bottom_track_9.mux_l3_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_8_127 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_26.mux_l2_in_0_/S mux_bottom_track_1.mux_l1_in_1_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 bottom_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0__S mux_right_track_12.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D mux_right_track_14.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_18.mux_l1_in_1__S mux_right_track_18.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_22.mux_l2_in_0_/S mux_right_track_24.mux_l1_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
Xmem_top_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_273 vgnd vpwr scs8hd_decap_4
XFILLER_31_240 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 _043_/HI vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_222 vgnd vpwr scs8hd_decap_3
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_18.scs8hd_buf_4_0__A mux_right_track_18.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_093_ _093_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_236 vpwr vgnd scs8hd_fill_2
XFILLER_6_258 vpwr vgnd scs8hd_fill_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D mux_top_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_228 vgnd vpwr scs8hd_fill_1
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_4
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
XFILLER_42_198 vgnd vpwr scs8hd_fill_1
XFILLER_32_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_250 vpwr vgnd scs8hd_fill_2
X_076_ chany_top_in[18] chany_bottom_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_33_132 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_0_ right_top_grid_pin_46_ chany_top_in[13] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[5] chany_top_in[1] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_209 vgnd vpwr scs8hd_decap_4
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_3
XFILLER_21_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vgnd vpwr scs8hd_decap_3
XFILLER_15_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A mux_bottom_track_33.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
X_059_ chany_bottom_in[3] chanx_right_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_246 vpwr vgnd scs8hd_fill_2
XFILLER_38_224 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_21_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_235 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_9.mux_l1_in_1_/S mux_bottom_track_9.mux_l2_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_190 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_238 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_32_208 vgnd vpwr scs8hd_decap_3
XFILLER_4_164 vpwr vgnd scs8hd_fill_2
XFILLER_4_186 vgnd vpwr scs8hd_decap_3
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_23_208 vgnd vpwr scs8hd_decap_6
XFILLER_23_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D mux_bottom_track_17.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_1_ _048_/HI mux_bottom_track_5.mux_l1_in_2_/X mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_6.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 mux_right_track_4.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_233 vgnd vpwr scs8hd_fill_1
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
X_092_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_37_119 vgnd vpwr scs8hd_fill_1
XFILLER_5_270 vgnd vpwr scs8hd_decap_6
XFILLER_36_152 vgnd vpwr scs8hd_fill_1
XFILLER_36_141 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[17] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
X_075_ _075_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_33_166 vpwr vgnd scs8hd_fill_2
XFILLER_33_144 vgnd vpwr scs8hd_fill_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D mux_top_track_32.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_188 vgnd vpwr scs8hd_decap_4
X_058_ chany_bottom_in[1] chanx_right_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_38_236 vgnd vpwr scs8hd_fill_1
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XFILLER_38_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_29_258 vpwr vgnd scs8hd_fill_2
XFILLER_29_214 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_9.mux_l1_in_1_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_195 vgnd vpwr scs8hd_decap_3
XFILLER_26_206 vpwr vgnd scs8hd_fill_2
XFILLER_41_209 vpwr vgnd scs8hd_fill_2
XFILLER_34_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XFILLER_27_98 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_4_198 vgnd vpwr scs8hd_decap_3
XFILLER_4_154 vpwr vgnd scs8hd_fill_2
XFILLER_4_143 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D mux_top_track_32.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_231 vgnd vpwr scs8hd_decap_4
XFILLER_1_102 vpwr vgnd scs8hd_fill_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 _036_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_091_ _091_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_10_201 vpwr vgnd scs8hd_fill_2
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__S mux_top_track_16.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_36_164 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_1_ chanx_right_in[10] chanx_right_in[3] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XANTENNA__062__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_142 vpwr vgnd scs8hd_fill_2
XFILLER_35_98 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
X_074_ _074_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 mux_bottom_track_5.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__057__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.scs8hd_buf_4_0__A mux_right_track_4.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0__A0 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_30_126 vpwr vgnd scs8hd_fill_2
XFILLER_15_167 vgnd vpwr scs8hd_decap_4
XFILLER_15_178 vgnd vpwr scs8hd_decap_4
X_057_ chany_bottom_in[0] chanx_right_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_119 vgnd vpwr scs8hd_decap_6
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_35_218 vgnd vpwr scs8hd_decap_3
XFILLER_7_152 vpwr vgnd scs8hd_fill_2
X_109_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_34_273 vpwr vgnd scs8hd_fill_2
XANTENNA__070__A _070_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_207 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_232 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_14.mux_l2_in_0_/S mux_right_track_14.mux_l3_in_0_/S
+ mem_right_track_14.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__065__A _065_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_254 vgnd vpwr scs8hd_decap_8
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_20.mux_l1_in_1__A0 _029_/HI vgnd vpwr scs8hd_diode_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_169 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.mux_l1_in_1__S mux_right_track_6.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ ccff_tail mux_bottom_track_33.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_236 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 mux_top_track_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_4
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
X_090_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_206 vpwr vgnd scs8hd_fill_2
XFILLER_6_228 vpwr vgnd scs8hd_fill_2
XFILLER_10_257 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D mux_right_track_2.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_fill_1
XFILLER_36_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_20.mux_l2_in_0__A0 mux_right_track_20.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A mux_bottom_track_3.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_33.mux_l1_in_1_ _047_/HI chanx_right_in[13] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_168 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_073_ _073_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D mux_top_track_16.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_132 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_3__A0 _034_/HI vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.scs8hd_buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _075_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_right_track_26.scs8hd_buf_4_0__A mux_right_track_26.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0__A1 mux_right_track_12.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_30_149 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
X_056_ _056_/A chanx_right_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_21_149 vgnd vpwr scs8hd_decap_4
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_3
XFILLER_12_149 vpwr vgnd scs8hd_fill_2
XFILLER_20_182 vpwr vgnd scs8hd_fill_2
XFILLER_20_193 vpwr vgnd scs8hd_fill_2
X_108_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
X_039_ _039_/HI _039_/LO vgnd vpwr scs8hd_conb_1
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XFILLER_40_200 vgnd vpwr scs8hd_fill_1
XFILLER_25_263 vpwr vgnd scs8hd_fill_2
XFILLER_25_241 vgnd vpwr scs8hd_fill_1
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_211 vgnd vpwr scs8hd_decap_4
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D mux_right_track_4.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_14.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_14.mux_l1_in_0_/S mux_right_track_14.mux_l2_in_0_/S
+ mem_right_track_14.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_20.mux_l1_in_1__A1 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA__081__A chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_1_126 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S mux_top_track_24.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_222 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_192 vpwr vgnd scs8hd_fill_2
XFILLER_39_163 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_20.mux_l2_in_0__A1 mux_right_track_20.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
Xmux_top_track_24.mux_l2_in_1_ _039_/HI chany_bottom_in[18] mux_top_track_24.mux_l2_in_1_/S
+ mux_top_track_24.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__D mux_right_track_22.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_27_188 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_33.mux_l1_in_0_ chanx_right_in[6] chany_top_in[10] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_147 vgnd vpwr scs8hd_decap_8
XFILLER_2_254 vgnd vpwr scs8hd_decap_4
XFILLER_2_210 vpwr vgnd scs8hd_fill_2
X_072_ _072_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_136 vpwr vgnd scs8hd_fill_2
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_33_103 vgnd vpwr scs8hd_decap_6
XFILLER_18_177 vpwr vgnd scs8hd_fill_2
XFILLER_18_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_26.mux_l2_in_0__S mux_right_track_26.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.scs8hd_buf_4_0_ mux_right_track_14.mux_l3_in_0_/X _068_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_2_93 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l1_in_3__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
X_055_ _055_/HI _055_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l3_in_0_ mux_right_track_12.mux_l2_in_1_/X mux_right_track_12.mux_l2_in_0_/X
+ mux_right_track_12.mux_l3_in_0_/S mux_right_track_12.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 mux_top_track_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_206 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_180 vgnd vpwr scs8hd_decap_4
XFILLER_29_239 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__D mux_right_track_4.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA__084__A chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_28_261 vgnd vpwr scs8hd_decap_12
X_107_ _107_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_8
XFILLER_7_143 vgnd vpwr scs8hd_decap_3
XFILLER_7_187 vpwr vgnd scs8hd_fill_2
X_038_ _038_/HI _038_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_275 vpwr vgnd scs8hd_fill_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XFILLER_25_220 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_1_ _052_/HI chany_bottom_in[10] mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_12.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_0.mux_l2_in_1_ _050_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_253 vgnd vpwr scs8hd_decap_4
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_12.mux_l3_in_0_/S mux_right_track_14.mux_l1_in_0_/S
+ mem_right_track_14.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D mux_right_track_22.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_201 vpwr vgnd scs8hd_fill_2
XFILLER_13_234 vgnd vpwr scs8hd_decap_4
XFILLER_13_245 vgnd vpwr scs8hd_decap_3
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XFILLER_0_171 vpwr vgnd scs8hd_fill_2
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_1__A0 _053_/HI vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[2] right_top_grid_pin_48_ mux_right_track_0.mux_l1_in_2_/S
+ mux_right_track_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_226 vgnd vpwr scs8hd_decap_4
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_right_track_22.scs8hd_buf_4_0_ mux_right_track_22.mux_l2_in_0_/X _064_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_17.mux_l2_in_1_/S
+ mux_bottom_track_17.mux_l3_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
Xmux_top_track_24.mux_l2_in_0_ chany_bottom_in[9] mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_1_/S mux_top_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_6
XFILLER_27_178 vgnd vpwr scs8hd_decap_4
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_071_ _071_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_2_233 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l3_in_0__A0 mux_right_track_14.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2__S mux_top_track_8.mux_l1_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XFILLER_15_104 vgnd vpwr scs8hd_fill_1
XFILLER_15_137 vpwr vgnd scs8hd_fill_2
XFILLER_23_181 vpwr vgnd scs8hd_fill_2
X_054_ _054_/HI _054_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.scs8hd_buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _113_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vgnd vpwr scs8hd_decap_12
XFILLER_21_129 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vpwr vgnd scs8hd_fill_2
XFILLER_28_273 vpwr vgnd scs8hd_fill_2
X_106_ chany_bottom_in[8] chany_top_out[9] vgnd vpwr scs8hd_buf_2
X_037_ _037_/HI _037_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_80 vgnd vpwr scs8hd_decap_12
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_40_235 vgnd vpwr scs8hd_decap_8
XFILLER_40_224 vgnd vpwr scs8hd_decap_8
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.mux_l2_in_0_ right_top_grid_pin_44_ mux_right_track_12.mux_l1_in_0_/X
+ mux_right_track_12.mux_l2_in_0_/S mux_right_track_12.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_158 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_32.mux_l2_in_0__S mux_top_track_32.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_fill_1
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vpwr vgnd scs8hd_fill_2
XFILLER_3_180 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_1_106 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D mux_right_track_8.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D mux_bottom_track_25.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_1__A1 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_1_ right_top_grid_pin_46_ right_top_grid_pin_44_ mux_right_track_0.mux_l1_in_2_/S
+ mux_right_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_2.mux_l2_in_1_ _038_/HI chany_bottom_in[13] mux_top_track_2.mux_l2_in_0_/S
+ mux_top_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l2_in_1_ _031_/HI chany_bottom_in[19] mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XFILLER_36_168 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l2_in_1_/S mem_bottom_track_17.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_35_190 vpwr vgnd scs8hd_fill_2
XFILLER_27_146 vpwr vgnd scs8hd_fill_2
X_070_ _070_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_41_193 vgnd vpwr scs8hd_decap_6
XFILLER_41_171 vgnd vpwr scs8hd_decap_6
XPHY_80 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_14.mux_l3_in_0__A1 mux_right_track_14.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_190 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l3_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XFILLER_24_149 vpwr vgnd scs8hd_fill_2
XFILLER_32_182 vpwr vgnd scs8hd_fill_2
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XANTENNA__098__A chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_23_160 vpwr vgnd scs8hd_fill_2
X_053_ _053_/HI _053_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[6] mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_22.mux_l2_in_0__S mux_right_track_22.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_274 vgnd vpwr scs8hd_decap_3
XFILLER_37_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
X_105_ chany_bottom_in[9] chany_top_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_24.mux_l3_in_0__S mux_top_track_24.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_036_ _036_/HI _036_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XFILLER_34_244 vpwr vgnd scs8hd_fill_2
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_233 vpwr vgnd scs8hd_fill_2
XFILLER_40_247 vgnd vpwr scs8hd_decap_8
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_200 vgnd vpwr scs8hd_decap_3
XFILLER_16_222 vpwr vgnd scs8hd_fill_2
XFILLER_16_266 vgnd vpwr scs8hd_decap_8
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vpwr vgnd scs8hd_fill_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A0 _044_/HI vgnd vpwr scs8hd_diode_2
XFILLER_9_218 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_ chany_top_in[15] chany_top_in[10] mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_8_273 vpwr vgnd scs8hd_fill_2
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_ right_top_grid_pin_42_ chany_top_in[2] mux_right_track_0.mux_l1_in_2_/S
+ mux_right_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_10_206 vgnd vpwr scs8hd_decap_6
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l2_in_0_ chany_bottom_in[18] mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_276 vgnd vpwr scs8hd_fill_1
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_36_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A0 mux_bottom_track_17.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_9.mux_l3_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_18.mux_l1_in_1__A0 _055_/HI vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_169 vgnd vpwr scs8hd_decap_3
XFILLER_2_202 vpwr vgnd scs8hd_fill_2
XFILLER_2_224 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
Xmem_right_track_22.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_22.mux_l1_in_0_/S mux_right_track_22.mux_l2_in_0_/S
+ mem_right_track_22.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_14.mux_l3_in_0__S mux_right_track_14.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_2.mux_l1_in_1_ chany_bottom_in[4] chanx_right_in[16] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_180 vgnd vpwr scs8hd_fill_1
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
X_052_ _052_/HI _052_/LO vgnd vpwr scs8hd_conb_1
Xmem_right_track_6.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l3_in_0_/S
+ mem_right_track_6.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_18.mux_l2_in_0__A0 mux_right_track_18.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_20_186 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_253 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
X_104_ chany_bottom_in[10] chany_top_out[11] vgnd vpwr scs8hd_buf_2
X_035_ _035_/HI _035_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_1_ _043_/HI mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_142 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vgnd vpwr scs8hd_decap_4
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_34_201 vpwr vgnd scs8hd_fill_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A0 _045_/HI vgnd vpwr scs8hd_diode_2
XFILLER_25_267 vgnd vpwr scs8hd_decap_8
XFILLER_25_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A1 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[19] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_226 vpwr vgnd scs8hd_fill_2
XFILLER_21_270 vgnd vpwr scs8hd_decap_6
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A0 mux_bottom_track_25.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.scs8hd_buf_4_0__A mux_top_track_16.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_167 vpwr vgnd scs8hd_fill_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_6
XFILLER_5_222 vgnd vpwr scs8hd_decap_3
XFILLER_5_266 vpwr vgnd scs8hd_fill_2
XFILLER_36_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A1 mux_bottom_track_17.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_18.mux_l1_in_1__A1 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_35_170 vpwr vgnd scs8hd_fill_2
Xmem_right_track_22.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_20.mux_l2_in_0_/S mux_right_track_22.mux_l1_in_0_/S
+ mem_right_track_22.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_26.mux_l2_in_0__A0 _032_/HI vgnd vpwr scs8hd_diode_2
XFILLER_41_140 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.mux_l3_in_0__S mux_right_track_6.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_0.mux_l3_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ mem_top_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_top_track_2.mux_l1_in_0_ chanx_right_in[9] chanx_right_in[2] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l1_in_0_ right_top_grid_pin_42_ chany_top_in[18] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_107 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_051_ _051_/HI _051_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_173 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_3
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D mux_top_track_24.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_6.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_6.mux_l1_in_0_/S mux_right_track_6.mux_l2_in_1_/S
+ mem_right_track_6.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_6.scs8hd_buf_4_0_ mux_right_track_6.mux_l3_in_0_/X _072_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_right_track_18.mux_l2_in_0__A1 mux_right_track_18.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.scs8hd_buf_4_0__A mux_right_track_16.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_254 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_20_165 vpwr vgnd scs8hd_fill_2
XFILLER_28_210 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l3_in_0_/S mem_bottom_track_25.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _103_/A chany_top_out[12] vgnd vpwr scs8hd_buf_2
X_034_ _034_/HI _034_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_7 vgnd vpwr scs8hd_decap_12
XFILLER_19_221 vpwr vgnd scs8hd_fill_2
XFILLER_19_232 vpwr vgnd scs8hd_fill_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_1__S mux_bottom_track_33.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_205 vgnd vpwr scs8hd_decap_8
XFILLER_4_139 vpwr vgnd scs8hd_fill_2
XFILLER_4_117 vgnd vpwr scs8hd_fill_1
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0__S mux_right_track_12.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_1_ chanx_right_in[12] chanx_right_in[5] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_205 vpwr vgnd scs8hd_fill_2
XFILLER_0_175 vgnd vpwr scs8hd_decap_4
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D mux_top_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A1 mux_bottom_track_25.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_231 vpwr vgnd scs8hd_fill_2
XFILLER_12_260 vpwr vgnd scs8hd_fill_2
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XFILLER_39_146 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_201 vpwr vgnd scs8hd_fill_2
XFILLER_5_245 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_36_149 vgnd vpwr scs8hd_fill_1
XFILLER_36_105 vgnd vpwr scs8hd_decap_3
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__D mux_right_track_10.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_237 vpwr vgnd scs8hd_fill_2
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_26.mux_l2_in_0__A1 mux_right_track_26.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XFILLER_41_152 vpwr vgnd scs8hd_fill_2
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_160 vgnd vpwr scs8hd_decap_3
XFILLER_32_174 vpwr vgnd scs8hd_fill_2
X_050_ _050_/HI _050_/LO vgnd vpwr scs8hd_conb_1
Xmem_right_track_6.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_4.mux_l3_in_0_/S mux_right_track_6.mux_l1_in_0_/S
+ mem_right_track_6.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_163 vpwr vgnd scs8hd_fill_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__S mux_bottom_track_25.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l3_in_0__S mux_right_track_10.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 _050_/HI vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/S mem_bottom_track_25.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
X_033_ _033_/HI _033_/LO vgnd vpwr scs8hd_conb_1
X_102_ chany_bottom_in[12] chany_top_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_7_148 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D mux_top_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_192 vpwr vgnd scs8hd_fill_2
XFILLER_25_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D mux_right_track_26.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_217 vpwr vgnd scs8hd_fill_2
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_228 vpwr vgnd scs8hd_fill_2
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__104__A chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_3_162 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_2__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__D mux_right_track_10.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_fill_1
XFILLER_8_254 vgnd vpwr scs8hd_decap_8
XFILLER_8_265 vgnd vpwr scs8hd_decap_8
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_12_272 vgnd vpwr scs8hd_decap_3
XFILLER_5_98 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_117 vpwr vgnd scs8hd_fill_2
XFILLER_29_191 vpwr vgnd scs8hd_fill_2
XFILLER_18_117 vpwr vgnd scs8hd_fill_2
XFILLER_18_128 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_131 vpwr vgnd scs8hd_fill_2
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_194 vgnd vpwr scs8hd_decap_8
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XANTENNA__112__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_271 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D mux_top_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_172 vpwr vgnd scs8hd_fill_2
XFILLER_32_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__S mux_right_track_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_186 vpwr vgnd scs8hd_fill_2
XFILLER_14_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_201 vgnd vpwr scs8hd_decap_4
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_19 vgnd vpwr scs8hd_decap_12
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_17.mux_l3_in_0_/S
+ mux_bottom_track_25.mux_l1_in_1_/S mem_bottom_track_25.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
X_101_ chany_bottom_in[13] chany_top_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_127 vgnd vpwr scs8hd_fill_1
X_032_ _032_/HI _032_/LO vgnd vpwr scs8hd_conb_1
XFILLER_19_245 vgnd vpwr scs8hd_decap_8
XFILLER_34_248 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_8
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_25_237 vgnd vpwr scs8hd_decap_4
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vpwr vgnd scs8hd_fill_2
XFILLER_16_226 vgnd vpwr scs8hd_decap_4
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_152 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.scs8hd_buf_4_0__A mux_right_track_2.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_159 vpwr vgnd scs8hd_fill_2
XFILLER_39_115 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_20.mux_l1_in_1__S mux_right_track_20.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_4
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_2__D mux_right_track_14.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_206 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_165 vgnd vpwr scs8hd_decap_4
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_fill_1
XFILLER_32_143 vgnd vpwr scs8hd_decap_4
Xmem_right_track_12.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_12.mux_l2_in_0_/S mux_right_track_12.mux_l3_in_0_/S
+ mem_right_track_12.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_24.scs8hd_buf_4_0__A mux_top_track_24.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_110 vgnd vpwr scs8hd_decap_12
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_11_98 vgnd vpwr scs8hd_decap_8
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
XFILLER_37_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_135 vgnd vpwr scs8hd_fill_1
XFILLER_9_191 vpwr vgnd scs8hd_fill_2
XFILLER_28_224 vpwr vgnd scs8hd_fill_2
X_100_ chany_bottom_in[14] chany_top_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_7_139 vpwr vgnd scs8hd_fill_2
XFILLER_11_146 vpwr vgnd scs8hd_fill_2
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
X_031_ _031_/HI _031_/LO vgnd vpwr scs8hd_conb_1
XFILLER_34_205 vgnd vpwr scs8hd_decap_6
Xmux_top_track_16.scs8hd_buf_4_0_ mux_top_track_16.mux_l3_in_0_/X _107_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_6_150 vgnd vpwr scs8hd_fill_1
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_249 vpwr vgnd scs8hd_fill_2
XFILLER_25_216 vpwr vgnd scs8hd_fill_2
XFILLER_33_271 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A mux_bottom_track_1.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_249 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XFILLER_22_208 vgnd vpwr scs8hd_decap_6
XFILLER_22_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.scs8hd_buf_4_0__A mux_right_track_24.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_1__S mux_right_track_12.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_230 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D mux_right_track_16.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S mux_top_track_32.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_3__A0 _028_/HI vgnd vpwr scs8hd_diode_2
XFILLER_12_230 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_3_ _034_/HI chany_bottom_in[6] mux_right_track_6.mux_l1_in_0_/S
+ mux_right_track_6.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_35_174 vpwr vgnd scs8hd_fill_2
XFILLER_35_141 vpwr vgnd scs8hd_fill_2
Xmux_top_track_32.mux_l2_in_1_ _040_/HI chany_bottom_in[10] mux_top_track_32.mux_l2_in_1_/S
+ mux_top_track_32.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_229 vpwr vgnd scs8hd_fill_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_163 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_86 vgnd vpwr scs8hd_decap_12
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_240 vgnd vpwr scs8hd_fill_1
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_199 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D mux_top_track_8.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_12.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_12.mux_l1_in_0_/S mux_right_track_12.mux_l2_in_0_/S
+ mem_right_track_12.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_144 vgnd vpwr scs8hd_decap_3
XFILLER_23_177 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S mux_right_track_6.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_24.scs8hd_buf_4_0_ mux_top_track_24.mux_l3_in_0_/X _103_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_37_258 vgnd vpwr scs8hd_decap_4
XFILLER_20_169 vpwr vgnd scs8hd_fill_2
XFILLER_28_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
X_030_ _030_/HI _030_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_169 vgnd vpwr scs8hd_decap_4
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__D mux_right_track_16.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_225 vpwr vgnd scs8hd_fill_2
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l2_in_1_ mux_right_track_6.mux_l1_in_3_/X mux_right_track_6.mux_l1_in_2_/X
+ mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1__A0 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_4
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_110 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_176 vgnd vpwr scs8hd_decap_4
XFILLER_30_231 vpwr vgnd scs8hd_fill_2
XFILLER_15_272 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_3.scs8hd_buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _094_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_13_209 vpwr vgnd scs8hd_fill_2
XFILLER_21_220 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.scs8hd_buf_4_0_ mux_right_track_10.mux_l3_in_0_/X _070_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_0_135 vpwr vgnd scs8hd_fill_2
XFILLER_0_179 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l1_in_3__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_264 vgnd vpwr scs8hd_decap_8
Xmux_right_track_6.mux_l1_in_2_ right_top_grid_pin_49_ right_top_grid_pin_47_ mux_right_track_6.mux_l1_in_0_/S
+ mux_right_track_6.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_33.mux_l1_in_1_/S
+ ccff_tail mem_bottom_track_33.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_106 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 mux_top_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_183 vgnd vpwr scs8hd_fill_1
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A0 chany_top_in[15] vgnd vpwr scs8hd_diode_2
Xmux_top_track_32.mux_l2_in_0_ chanx_right_in[14] mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_1_/S mux_top_track_32.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_32.scs8hd_buf_4_0_ mux_top_track_32.mux_l3_in_0_/X _099_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_4
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_120 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XFILLER_25_98 vgnd vpwr scs8hd_decap_8
XFILLER_1_263 vpwr vgnd scs8hd_fill_2
XFILLER_1_230 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vpwr vgnd scs8hd_fill_2
Xmem_right_track_12.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_10.mux_l3_in_0_/S mux_right_track_12.mux_l1_in_0_/S
+ mem_right_track_12.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_123 vgnd vpwr scs8hd_decap_6
XFILLER_23_156 vpwr vgnd scs8hd_fill_2
XFILLER_14_134 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
XFILLER_14_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_26.mux_l1_in_0__S mux_right_track_26.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_226 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_16.mux_l2_in_1_/S mux_top_track_16.mux_l3_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 _046_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D mux_top_track_32.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_1__A0 _051_/HI vgnd vpwr scs8hd_diode_2
XFILLER_19_204 vpwr vgnd scs8hd_fill_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A mux_bottom_track_9.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
Xmux_right_track_18.mux_l2_in_0_ mux_right_track_18.mux_l1_in_1_/X mux_right_track_18.mux_l1_in_0_/X
+ mux_right_track_18.mux_l2_in_0_/S mux_right_track_18.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
X_089_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_163 vgnd vpwr scs8hd_decap_4
XFILLER_6_196 vgnd vpwr scs8hd_decap_4
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__060__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
Xmux_right_track_20.mux_l2_in_0_ mux_right_track_20.mux_l1_in_1_/X mux_right_track_20.mux_l1_in_0_/X
+ mux_right_track_20.mux_l2_in_0_/S mux_right_track_20.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D mux_bottom_track_9.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l3_in_0__A0 mux_right_track_10.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_80 vpwr vgnd scs8hd_fill_2
XFILLER_21_254 vgnd vpwr scs8hd_decap_6
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_20.mux_l1_in_0__A0 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_125 vgnd vpwr scs8hd_decap_4
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
Xmux_right_track_18.mux_l1_in_1_ _055_/HI chany_bottom_in[14] mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_243 vpwr vgnd scs8hd_fill_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l1_in_1_ right_top_grid_pin_45_ right_top_grid_pin_43_ mux_right_track_6.mux_l1_in_0_/S
+ mux_right_track_6.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_33.mux_l1_in_1_/S mem_bottom_track_33.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
Xmux_top_track_8.mux_l2_in_1_ _042_/HI mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_20.mux_l1_in_1_ _029_/HI chany_bottom_in[16] mux_right_track_20.mux_l1_in_0_/S
+ mux_right_track_20.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D mux_right_track_0.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.scs8hd_buf_4_0_ mux_top_track_0.mux_l3_in_0_/X _115_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1__S mux_bottom_track_9.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_4_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
XFILLER_35_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_41_179 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_2_ chany_bottom_in[16] chany_bottom_in[6] mux_top_track_8.mux_l1_in_2_/S
+ mux_top_track_8.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_18.mux_l2_in_0__S mux_right_track_18.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_110 vgnd vpwr scs8hd_fill_1
XFILLER_17_121 vgnd vpwr scs8hd_fill_1
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_17_176 vgnd vpwr scs8hd_decap_4
XFILLER_40_190 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_2__A0 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XANTENNA__063__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_top_track_32.mux_l1_in_0_ chanx_right_in[7] chanx_right_in[0] mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_16.mux_l1_in_1_/S mux_top_track_16.mux_l2_in_1_/S
+ mem_top_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_149 vpwr vgnd scs8hd_fill_2
XFILLER_28_249 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_1__A1 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.scs8hd_buf_4_0__A mux_top_track_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_142 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l2_in_1__A0 mux_right_track_6.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
X_088_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D mux_right_track_0.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_271 vgnd vpwr scs8hd_decap_4
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_11 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.scs8hd_buf_4_0__A mux_top_track_32.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_200 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l3_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_230 vpwr vgnd scs8hd_fill_2
XFILLER_30_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D mux_top_track_8.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l3_in_0__A1 mux_right_track_10.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_92 vgnd vpwr scs8hd_fill_1
XFILLER_21_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_20.mux_l1_in_0__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_0_104 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
Xmux_right_track_18.mux_l1_in_0_ right_top_grid_pin_47_ chany_top_in[14] mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_6.mux_l3_in_0__A0 mux_right_track_6.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_211 vgnd vpwr scs8hd_fill_1
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_204 vgnd vpwr scs8hd_decap_8
XFILLER_8_215 vgnd vpwr scs8hd_decap_3
Xmux_right_track_6.mux_l1_in_0_ chany_top_in[6] chany_top_in[3] mux_right_track_6.mux_l1_in_0_/S
+ mux_right_track_6.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_119 vgnd vpwr scs8hd_decap_3
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__S mux_top_track_32.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_20.mux_l1_in_0_ right_top_grid_pin_48_ chany_top_in[16] mux_right_track_20.mux_l1_in_0_/S
+ mux_right_track_20.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__D mux_right_track_18.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_152 vgnd vpwr scs8hd_fill_1
XFILLER_38_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__066__A _066_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_218 vpwr vgnd scs8hd_fill_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l1_in_2__S mux_right_track_6.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_174 vpwr vgnd scs8hd_fill_2
XFILLER_29_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XFILLER_26_133 vgnd vpwr scs8hd_decap_3
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l1_in_1_ chanx_right_in[18] chanx_right_in[11] mux_top_track_8.mux_l1_in_2_/S
+ mux_top_track_8.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
XFILLER_17_155 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.mux_l1_in_2__A1 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_23_136 vgnd vpwr scs8hd_decap_6
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_22_191 vpwr vgnd scs8hd_fill_2
XFILLER_37_239 vgnd vpwr scs8hd_decap_3
Xmem_top_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_8.mux_l3_in_0_/S mux_top_track_16.mux_l1_in_1_/S
+ mem_top_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vpwr vgnd scs8hd_fill_2
XFILLER_9_195 vpwr vgnd scs8hd_fill_2
XFILLER_28_228 vgnd vpwr scs8hd_decap_8
XFILLER_28_206 vpwr vgnd scs8hd_fill_2
XFILLER_11_106 vgnd vpwr scs8hd_decap_3
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_231 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_087_ _087_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_10_161 vgnd vpwr scs8hd_decap_4
XFILLER_10_183 vpwr vgnd scs8hd_fill_2
XFILLER_10_194 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l2_in_1__A1 mux_right_track_6.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 _038_/HI vgnd vpwr scs8hd_diode_2
XFILLER_33_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_22.mux_l1_in_0__S mux_right_track_22.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_23 vgnd vpwr scs8hd_decap_12
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_253 vpwr vgnd scs8hd_fill_2
Xmem_right_track_20.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_20.mux_l1_in_0_/S mux_right_track_20.mux_l2_in_0_/S
+ mem_right_track_20.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_264 vpwr vgnd scs8hd_fill_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l3_in_0__A1 mux_right_track_6.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_227 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_260 vpwr vgnd scs8hd_fill_2
XFILLER_38_186 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D mux_right_track_4.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0__A0 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_35_178 vgnd vpwr scs8hd_decap_3
XFILLER_35_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_26_145 vpwr vgnd scs8hd_fill_2
XANTENNA__077__A chany_top_in[17] vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_148 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_1_222 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[4] top_left_grid_pin_1_ mux_top_track_8.mux_l1_in_2_/S
+ mux_top_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_22_181 vgnd vpwr scs8hd_decap_3
XFILLER_9_152 vgnd vpwr scs8hd_decap_8
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XFILLER_20_129 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_14.mux_l2_in_0__S mux_right_track_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l3_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_22.mux_l1_in_1__A0 _030_/HI vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_42_243 vgnd vpwr scs8hd_decap_4
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l3_in_0__S mux_top_track_16.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_086_ chany_top_in[8] chany_bottom_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__D mux_right_track_6.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l3_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_35 vgnd vpwr scs8hd_decap_12
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
Xmem_right_track_20.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_18.mux_l2_in_0_/S mux_right_track_20.mux_l1_in_0_/S
+ mem_right_track_20.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_158 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_top_track_0.mux_l1_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_235 vgnd vpwr scs8hd_fill_1
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_22.mux_l2_in_0__A0 mux_right_track_22.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
X_069_ _069_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_191 vpwr vgnd scs8hd_fill_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_6
XFILLER_21_224 vgnd vpwr scs8hd_decap_6
XFILLER_0_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
Xmem_top_track_24.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_24.mux_l2_in_1_/S mux_top_track_24.mux_l3_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_4.mux_l1_in_2_/S mux_right_track_4.mux_l2_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_14.scs8hd_buf_4_0__A mux_right_track_14.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.scs8hd_buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _074_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_38_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0__A1 mux_right_track_14.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D mux_right_track_24.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_187 vpwr vgnd scs8hd_fill_2
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_168 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_267 vpwr vgnd scs8hd_fill_2
XFILLER_1_245 vpwr vgnd scs8hd_fill_2
XFILLER_17_113 vpwr vgnd scs8hd_fill_2
XFILLER_32_149 vgnd vpwr scs8hd_decap_4
XFILLER_32_116 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l1_in_2__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XFILLER_23_149 vpwr vgnd scs8hd_fill_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D mux_right_track_6.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__088__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_105 vgnd vpwr scs8hd_fill_1
XFILLER_14_138 vpwr vgnd scs8hd_fill_2
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0__S mux_right_track_6.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_131 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_36_274 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_5.mux_l1_in_0_/S mux_bottom_track_5.mux_l2_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_22.mux_l1_in_1__A1 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_208 vpwr vgnd scs8hd_fill_2
XFILLER_10_130 vgnd vpwr scs8hd_decap_4
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
X_085_ chany_top_in[9] chany_bottom_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_8.mux_l1_in_2_/S mux_top_track_8.mux_l2_in_1_/S
+ mem_top_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_47 vgnd vpwr scs8hd_decap_12
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_222 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_22.mux_l2_in_0__A1 mux_right_track_22.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
X_068_ _068_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_84 vgnd vpwr scs8hd_decap_8
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 mux_bottom_track_17.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_203 vpwr vgnd scs8hd_fill_2
Xmem_top_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_24.mux_l1_in_0_/S mux_top_track_24.mux_l2_in_1_/S
+ mem_top_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_2_/S
+ mem_right_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_247 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.scs8hd_buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X _091_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_32.mux_l2_in_1__S mux_top_track_32.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_16.scs8hd_buf_4_0_ mux_right_track_16.mux_l2_in_0_/X _067_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_158 vpwr vgnd scs8hd_fill_2
XFILLER_35_136 vgnd vpwr scs8hd_decap_3
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D mux_bottom_track_33.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_18.mux_l1_in_0__A0 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_34_191 vgnd vpwr scs8hd_fill_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_125 vgnd vpwr scs8hd_decap_8
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_91 vpwr vgnd scs8hd_fill_2
XFILLER_16_191 vgnd vpwr scs8hd_decap_3
XFILLER_31_161 vpwr vgnd scs8hd_fill_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A0 bottom_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_14_117 vpwr vgnd scs8hd_fill_2
XFILLER_22_161 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A0 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_110 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_231 vpwr vgnd scs8hd_fill_2
XFILLER_36_220 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_5.mux_l1_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_264 vpwr vgnd scs8hd_fill_2
XFILLER_27_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
X_084_ chany_top_in[10] chany_bottom_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
XFILLER_33_267 vpwr vgnd scs8hd_fill_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_3
Xmux_right_track_2.mux_l1_in_3_ _028_/HI chany_bottom_in[4] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 _049_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__S mux_bottom_track_25.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 mux_bottom_track_25.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0__S mux_right_track_10.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_4.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_2_/S
+ mem_top_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_24_245 vgnd vpwr scs8hd_decap_8
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_127 vgnd vpwr scs8hd_decap_4
Xmux_right_track_24.scs8hd_buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _063_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_30_215 vgnd vpwr scs8hd_decap_3
XFILLER_15_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
X_067_ _067_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_0_30 vgnd vpwr scs8hd_fill_1
XFILLER_0_52 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_0_108 vgnd vpwr scs8hd_decap_4
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
Xmem_top_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_16.mux_l3_in_0_/S mux_top_track_24.mux_l1_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XFILLER_12_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A0 mux_bottom_track_9.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_26.mux_l1_in_0__A0 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_38_145 vgnd vpwr scs8hd_decap_4
Xmux_right_track_14.mux_l3_in_0_ mux_right_track_14.mux_l2_in_1_/X mux_right_track_14.mux_l2_in_0_/X
+ mux_right_track_14.mux_l3_in_0_/S mux_right_track_14.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_178 vpwr vgnd scs8hd_fill_2
XFILLER_29_167 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_8
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_4_211 vgnd vpwr scs8hd_fill_1
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_34_170 vpwr vgnd scs8hd_fill_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A0 _047_/HI vgnd vpwr scs8hd_diode_2
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_236 vgnd vpwr scs8hd_decap_4
Xmux_right_track_14.mux_l2_in_1_ _053_/HI chany_bottom_in[12] mux_right_track_14.mux_l2_in_0_/S
+ mux_right_track_14.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.scs8hd_buf_4_0__A mux_right_track_0.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_39_240 vgnd vpwr scs8hd_decap_4
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l3_in_0__S mux_bottom_track_9.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A1 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_140 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A0 mux_bottom_track_33.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 _031_/HI vgnd vpwr scs8hd_diode_2
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_1__S mux_bottom_track_17.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_210 vgnd vpwr scs8hd_decap_4
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_1__A0 _037_/HI vgnd vpwr scs8hd_diode_2
X_083_ _083_/A chany_bottom_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_10_143 vgnd vpwr scs8hd_decap_6
XFILLER_10_165 vgnd vpwr scs8hd_fill_1
XFILLER_10_198 vgnd vpwr scs8hd_fill_1
XFILLER_6_169 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_2_ right_top_grid_pin_49_ right_top_grid_pin_47_ mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_210 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_224 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 mux_bottom_track_9.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_15_213 vpwr vgnd scs8hd_fill_2
XFILLER_15_268 vpwr vgnd scs8hd_fill_2
X_066_ _066_/A chanx_right_out[9] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_fill_1
Xmem_right_track_10.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_10.mux_l2_in_0_/S mux_right_track_10.mux_l3_in_0_/S
+ mem_right_track_10.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l3_in_0__A0 mux_top_track_16.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A1 mux_bottom_track_9.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D mux_top_track_16.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
X_049_ _049_/HI _049_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_264 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_38_179 vgnd vpwr scs8hd_decap_4
XFILLER_38_124 vpwr vgnd scs8hd_fill_2
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D mux_bottom_track_17.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_234 vpwr vgnd scs8hd_fill_2
XFILLER_26_149 vpwr vgnd scs8hd_fill_2
XFILLER_26_138 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_259 vpwr vgnd scs8hd_fill_2
XFILLER_1_226 vpwr vgnd scs8hd_fill_2
XFILLER_25_160 vgnd vpwr scs8hd_decap_4
XFILLER_40_196 vgnd vpwr scs8hd_decap_4
XFILLER_40_152 vgnd vpwr scs8hd_fill_1
XFILLER_40_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
Xmem_top_track_32.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_32.mux_l2_in_1_/S mux_top_track_32.mux_l3_in_0_/S
+ mem_top_track_32.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_14.mux_l2_in_0_ right_top_grid_pin_45_ mux_right_track_14.mux_l1_in_0_/X
+ mux_right_track_14.mux_l2_in_0_/S mux_right_track_14.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_171 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_22.scs8hd_buf_4_0__A mux_right_track_22.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_24.mux_l2_in_1__A0 _039_/HI vgnd vpwr scs8hd_diode_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XFILLER_13_174 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A1 mux_bottom_track_33.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_247 vgnd vpwr scs8hd_fill_1
XFILLER_42_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A1 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
X_082_ chany_top_in[12] chany_bottom_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_10_177 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_1_ right_top_grid_pin_45_ right_top_grid_pin_43_ mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_236 vgnd vpwr scs8hd_decap_6
XFILLER_33_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l3_in_0__A0 mux_top_track_24.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_1_ _041_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_1_/S
+ mux_top_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 _042_/HI vgnd vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_6
XFILLER_30_206 vgnd vpwr scs8hd_decap_6
X_065_ _065_/A chanx_right_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_2_162 vgnd vpwr scs8hd_fill_1
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_10.mux_l1_in_0_/S mux_right_track_10.mux_l2_in_0_/S
+ mem_right_track_10.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l3_in_0__A1 mux_top_track_16.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_2_ chany_bottom_in[14] chany_bottom_in[5] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
X_048_ _048_/HI _048_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_276 vgnd vpwr scs8hd_fill_1
XFILLER_38_158 vpwr vgnd scs8hd_fill_2
XFILLER_14_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l3_in_0__A0 mux_top_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_35_106 vpwr vgnd scs8hd_fill_2
XFILLER_28_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_32.mux_l2_in_1__A0 _040_/HI vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_180 vgnd vpwr scs8hd_fill_1
XFILLER_19_191 vpwr vgnd scs8hd_fill_2
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_249 vgnd vpwr scs8hd_decap_4
XFILLER_1_205 vpwr vgnd scs8hd_fill_2
XFILLER_17_117 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.scs8hd_buf_4_0__A mux_right_track_8.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA__102__A chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_top_track_32.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_32.mux_l1_in_0_/S mux_top_track_32.mux_l2_in_1_/S
+ mem_top_track_32.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_197 vgnd vpwr scs8hd_decap_3
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l2_in_1__A1 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_2__D mux_right_track_10.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_186 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_32.mux_l3_in_0__A0 mux_top_track_32.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_135 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S mux_bottom_track_17.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_226 vgnd vpwr scs8hd_fill_1
XFILLER_42_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_ chany_top_in[19] chany_top_in[12] mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
X_081_ chany_top_in[13] chany_bottom_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_6_138 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[4] chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l3_in_0__A1 mux_top_track_24.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_5_160 vpwr vgnd scs8hd_fill_2
Xmux_right_track_26.mux_l2_in_0_ _032_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_204 vgnd vpwr scs8hd_decap_3
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 mux_top_track_8.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
X_064_ _064_/A chanx_right_out[11] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_17.mux_l2_in_1_ _044_/HI chanx_right_in[15] mux_bottom_track_17.mux_l2_in_1_/S
+ mux_bottom_track_17.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D mux_top_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__110__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_2_185 vgnd vpwr scs8hd_decap_4
XFILLER_0_22 vpwr vgnd scs8hd_fill_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_4
Xmem_right_track_10.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_8.mux_l3_in_0_/S mux_right_track_10.mux_l1_in_0_/S
+ mem_right_track_10.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_207 vgnd vpwr scs8hd_decap_4
XFILLER_20_251 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_4.mux_l1_in_1_ chanx_right_in[17] chanx_right_in[10] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__105__A chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
X_047_ _047_/HI _047_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_8.mux_l3_in_0__A1 mux_top_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__D mux_right_track_12.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.scs8hd_buf_4_0_ mux_right_track_8.mux_l3_in_0_/X _071_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_94 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l2_in_1__A1 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_34_184 vgnd vpwr scs8hd_decap_4
XFILLER_26_107 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l2_in_1_ _046_/HI chanx_right_in[18] mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_40_154 vpwr vgnd scs8hd_fill_2
XFILLER_40_143 vgnd vpwr scs8hd_decap_6
XFILLER_25_184 vgnd vpwr scs8hd_decap_4
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_31_95 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
Xmem_top_track_32.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_24.mux_l3_in_0_/S mux_top_track_32.mux_l1_in_0_/S
+ mem_top_track_32.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_165 vpwr vgnd scs8hd_fill_2
XFILLER_31_132 vgnd vpwr scs8hd_decap_4
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_32.mux_l3_in_0__A1 mux_top_track_32.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D mux_top_track_4.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_235 vpwr vgnd scs8hd_fill_2
XFILLER_36_224 vpwr vgnd scs8hd_fill_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_4
XFILLER_27_268 vgnd vpwr scs8hd_decap_8
XFILLER_27_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D mux_bottom_track_1.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_080_ chany_top_in[14] chany_bottom_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_10_157 vpwr vgnd scs8hd_fill_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_12_97 vgnd vpwr scs8hd_decap_8
XFILLER_33_227 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.scs8hd_buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X _087_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__D mux_right_track_12.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_238 vgnd vpwr scs8hd_decap_4
Xmem_right_track_18.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_18.mux_l1_in_1_/S mux_right_track_18.mux_l2_in_0_/S
+ mem_right_track_18.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S mux_bottom_track_17.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
X_063_ _063_/A chanx_right_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_2__A0 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_ chanx_right_in[3] top_left_grid_pin_1_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_26.mux_l1_in_0_ chany_bottom_in[15] right_top_grid_pin_43_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
X_115_ _115_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_046_ _046_/HI _046_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_223 vpwr vgnd scs8hd_fill_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_4
XFILLER_38_149 vgnd vpwr scs8hd_fill_1
XFILLER_37_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_ chanx_right_in[8] chanx_right_in[1] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.scs8hd_buf_4_0__A mux_top_track_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_28_171 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
X_029_ _029_/HI _029_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_174 vgnd vpwr scs8hd_fill_1
XFILLER_34_163 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 mux_right_track_2.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_25_130 vgnd vpwr scs8hd_decap_8
XFILLER_40_177 vpwr vgnd scs8hd_fill_2
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XFILLER_16_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
.ends

