VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2203.920 BY 2005.840 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.130 1961.720 1193.410 1964.120 ;
    END
  END address[0]
  PIN address[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1675.670 44.120 1675.950 46.520 ;
    END
  END address[10]
  PIN address[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1676.160 2154.480 1676.760 ;
    END
  END address[11]
  PIN address[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1740.080 2154.480 1740.680 ;
    END
  END address[12]
  PIN address[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.610 44.120 1739.890 46.520 ;
    END
  END address[13]
  PIN address[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1808.760 51.880 1809.360 ;
    END
  END address[14]
  PIN address[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1803.550 44.120 1803.830 46.520 ;
    END
  END address[15]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1561.240 51.880 1561.840 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1612.240 2154.480 1612.840 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1623.120 51.880 1623.720 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1284.670 1961.720 1284.950 1964.120 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1685.000 51.880 1685.600 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.210 1961.720 1376.490 1964.120 ;
    END
  END address[6]
  PIN address[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1746.880 51.880 1747.480 ;
    END
  END address[7]
  PIN address[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1467.750 1961.720 1468.030 1964.120 ;
    END
  END address[8]
  PIN address[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1612.190 44.120 1612.470 46.520 ;
    END
  END address[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1559.290 1961.720 1559.570 1964.120 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1650.830 1961.720 1651.110 1964.120 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1870.640 51.880 1871.240 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 95.110 1961.720 95.390 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 460.810 1961.720 461.090 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[10]
  PIN gfpga_pad_GPIO_PAD[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 552.350 1961.720 552.630 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[11]
  PIN gfpga_pad_GPIO_PAD[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 643.890 1961.720 644.170 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[12]
  PIN gfpga_pad_GPIO_PAD[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 735.430 1961.720 735.710 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[13]
  PIN gfpga_pad_GPIO_PAD[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1994.910 44.120 1995.190 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[14]
  PIN gfpga_pad_GPIO_PAD[15]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1804.000 2154.480 1804.600 ;
    END
  END gfpga_pad_GPIO_PAD[15]
  PIN gfpga_pad_GPIO_PAD[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2016.990 1961.720 2017.270 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[16]
  PIN gfpga_pad_GPIO_PAD[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1867.920 2154.480 1868.520 ;
    END
  END gfpga_pad_GPIO_PAD[17]
  PIN gfpga_pad_GPIO_PAD[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2108.530 1961.720 2108.810 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[18]
  PIN gfpga_pad_GPIO_PAD[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2058.390 44.120 2058.670 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[19]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 186.190 1961.720 186.470 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 826.970 1961.720 827.250 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[20]
  PIN gfpga_pad_GPIO_PAD[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 918.510 1961.720 918.790 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[21]
  PIN gfpga_pad_GPIO_PAD[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1010.050 1961.720 1010.330 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[22]
  PIN gfpga_pad_GPIO_PAD[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1101.590 1961.720 1101.870 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[23]
  PIN gfpga_pad_GPIO_PAD[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 76.120 2154.480 76.720 ;
    END
  END gfpga_pad_GPIO_PAD[24]
  PIN gfpga_pad_GPIO_PAD[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 140.040 2154.480 140.640 ;
    END
  END gfpga_pad_GPIO_PAD[25]
  PIN gfpga_pad_GPIO_PAD[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 203.960 2154.480 204.560 ;
    END
  END gfpga_pad_GPIO_PAD[26]
  PIN gfpga_pad_GPIO_PAD[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 267.880 2154.480 268.480 ;
    END
  END gfpga_pad_GPIO_PAD[27]
  PIN gfpga_pad_GPIO_PAD[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 331.800 2154.480 332.400 ;
    END
  END gfpga_pad_GPIO_PAD[28]
  PIN gfpga_pad_GPIO_PAD[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 395.720 2154.480 396.320 ;
    END
  END gfpga_pad_GPIO_PAD[29]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 277.730 1961.720 278.010 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 459.640 2154.480 460.240 ;
    END
  END gfpga_pad_GPIO_PAD[30]
  PIN gfpga_pad_GPIO_PAD[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 523.560 2154.480 524.160 ;
    END
  END gfpga_pad_GPIO_PAD[31]
  PIN gfpga_pad_GPIO_PAD[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 588.160 2154.480 588.760 ;
    END
  END gfpga_pad_GPIO_PAD[32]
  PIN gfpga_pad_GPIO_PAD[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 652.080 2154.480 652.680 ;
    END
  END gfpga_pad_GPIO_PAD[33]
  PIN gfpga_pad_GPIO_PAD[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 716.000 2154.480 716.600 ;
    END
  END gfpga_pad_GPIO_PAD[34]
  PIN gfpga_pad_GPIO_PAD[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 779.920 2154.480 780.520 ;
    END
  END gfpga_pad_GPIO_PAD[35]
  PIN gfpga_pad_GPIO_PAD[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 843.840 2154.480 844.440 ;
    END
  END gfpga_pad_GPIO_PAD[36]
  PIN gfpga_pad_GPIO_PAD[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 907.760 2154.480 908.360 ;
    END
  END gfpga_pad_GPIO_PAD[37]
  PIN gfpga_pad_GPIO_PAD[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 971.680 2154.480 972.280 ;
    END
  END gfpga_pad_GPIO_PAD[38]
  PIN gfpga_pad_GPIO_PAD[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1036.280 2154.480 1036.880 ;
    END
  END gfpga_pad_GPIO_PAD[39]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 369.270 1961.720 369.550 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1100.200 2154.480 1100.800 ;
    END
  END gfpga_pad_GPIO_PAD[40]
  PIN gfpga_pad_GPIO_PAD[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1164.120 2154.480 1164.720 ;
    END
  END gfpga_pad_GPIO_PAD[41]
  PIN gfpga_pad_GPIO_PAD[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1228.040 2154.480 1228.640 ;
    END
  END gfpga_pad_GPIO_PAD[42]
  PIN gfpga_pad_GPIO_PAD[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1291.960 2154.480 1292.560 ;
    END
  END gfpga_pad_GPIO_PAD[43]
  PIN gfpga_pad_GPIO_PAD[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1355.880 2154.480 1356.480 ;
    END
  END gfpga_pad_GPIO_PAD[44]
  PIN gfpga_pad_GPIO_PAD[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1419.800 2154.480 1420.400 ;
    END
  END gfpga_pad_GPIO_PAD[45]
  PIN gfpga_pad_GPIO_PAD[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1483.720 2154.480 1484.320 ;
    END
  END gfpga_pad_GPIO_PAD[46]
  PIN gfpga_pad_GPIO_PAD[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1548.320 2154.480 1548.920 ;
    END
  END gfpga_pad_GPIO_PAD[47]
  PIN gfpga_pad_GPIO_PAD[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.310 44.120 81.590 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[48]
  PIN gfpga_pad_GPIO_PAD[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 144.790 44.120 145.070 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[49]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1867.030 44.120 1867.310 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 208.730 44.120 209.010 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[50]
  PIN gfpga_pad_GPIO_PAD[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 272.670 44.120 272.950 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[51]
  PIN gfpga_pad_GPIO_PAD[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 336.150 44.120 336.430 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[52]
  PIN gfpga_pad_GPIO_PAD[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 400.090 44.120 400.370 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[53]
  PIN gfpga_pad_GPIO_PAD[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 464.030 44.120 464.310 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[54]
  PIN gfpga_pad_GPIO_PAD[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 527.510 44.120 527.790 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[55]
  PIN gfpga_pad_GPIO_PAD[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 591.450 44.120 591.730 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[56]
  PIN gfpga_pad_GPIO_PAD[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 655.390 44.120 655.670 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[57]
  PIN gfpga_pad_GPIO_PAD[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 718.870 44.120 719.150 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[58]
  PIN gfpga_pad_GPIO_PAD[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 782.810 44.120 783.090 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[59]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1742.370 1961.720 1742.650 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 846.750 44.120 847.030 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[60]
  PIN gfpga_pad_GPIO_PAD[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 910.230 44.120 910.510 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[61]
  PIN gfpga_pad_GPIO_PAD[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 974.170 44.120 974.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[62]
  PIN gfpga_pad_GPIO_PAD[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1038.110 44.120 1038.390 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[63]
  PIN gfpga_pad_GPIO_PAD[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1101.590 44.120 1101.870 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[64]
  PIN gfpga_pad_GPIO_PAD[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1165.530 44.120 1165.810 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[65]
  PIN gfpga_pad_GPIO_PAD[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1229.470 44.120 1229.750 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[66]
  PIN gfpga_pad_GPIO_PAD[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1292.950 44.120 1293.230 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[67]
  PIN gfpga_pad_GPIO_PAD[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1356.890 44.120 1357.170 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[68]
  PIN gfpga_pad_GPIO_PAD[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1420.830 44.120 1421.110 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[69]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1930.970 44.120 1931.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1484.310 44.120 1484.590 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[70]
  PIN gfpga_pad_GPIO_PAD[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1548.250 44.120 1548.530 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[71]
  PIN gfpga_pad_GPIO_PAD[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 74.760 51.880 75.360 ;
    END
  END gfpga_pad_GPIO_PAD[72]
  PIN gfpga_pad_GPIO_PAD[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 136.640 51.880 137.240 ;
    END
  END gfpga_pad_GPIO_PAD[73]
  PIN gfpga_pad_GPIO_PAD[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 198.520 51.880 199.120 ;
    END
  END gfpga_pad_GPIO_PAD[74]
  PIN gfpga_pad_GPIO_PAD[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 260.400 51.880 261.000 ;
    END
  END gfpga_pad_GPIO_PAD[75]
  PIN gfpga_pad_GPIO_PAD[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 322.280 51.880 322.880 ;
    END
  END gfpga_pad_GPIO_PAD[76]
  PIN gfpga_pad_GPIO_PAD[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 384.160 51.880 384.760 ;
    END
  END gfpga_pad_GPIO_PAD[77]
  PIN gfpga_pad_GPIO_PAD[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 446.040 51.880 446.640 ;
    END
  END gfpga_pad_GPIO_PAD[78]
  PIN gfpga_pad_GPIO_PAD[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 507.920 51.880 508.520 ;
    END
  END gfpga_pad_GPIO_PAD[79]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1833.910 1961.720 1834.190 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN gfpga_pad_GPIO_PAD[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 569.800 51.880 570.400 ;
    END
  END gfpga_pad_GPIO_PAD[80]
  PIN gfpga_pad_GPIO_PAD[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 631.680 51.880 632.280 ;
    END
  END gfpga_pad_GPIO_PAD[81]
  PIN gfpga_pad_GPIO_PAD[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 693.560 51.880 694.160 ;
    END
  END gfpga_pad_GPIO_PAD[82]
  PIN gfpga_pad_GPIO_PAD[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 756.120 51.880 756.720 ;
    END
  END gfpga_pad_GPIO_PAD[83]
  PIN gfpga_pad_GPIO_PAD[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 818.000 51.880 818.600 ;
    END
  END gfpga_pad_GPIO_PAD[84]
  PIN gfpga_pad_GPIO_PAD[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 879.880 51.880 880.480 ;
    END
  END gfpga_pad_GPIO_PAD[85]
  PIN gfpga_pad_GPIO_PAD[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 941.760 51.880 942.360 ;
    END
  END gfpga_pad_GPIO_PAD[86]
  PIN gfpga_pad_GPIO_PAD[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1003.640 51.880 1004.240 ;
    END
  END gfpga_pad_GPIO_PAD[87]
  PIN gfpga_pad_GPIO_PAD[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1065.520 51.880 1066.120 ;
    END
  END gfpga_pad_GPIO_PAD[88]
  PIN gfpga_pad_GPIO_PAD[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1127.400 51.880 1128.000 ;
    END
  END gfpga_pad_GPIO_PAD[89]
  PIN gfpga_pad_GPIO_PAD[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1932.520 51.880 1933.120 ;
    END
  END gfpga_pad_GPIO_PAD[8]
  PIN gfpga_pad_GPIO_PAD[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1189.280 51.880 1189.880 ;
    END
  END gfpga_pad_GPIO_PAD[90]
  PIN gfpga_pad_GPIO_PAD[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1251.160 51.880 1251.760 ;
    END
  END gfpga_pad_GPIO_PAD[91]
  PIN gfpga_pad_GPIO_PAD[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1313.040 51.880 1313.640 ;
    END
  END gfpga_pad_GPIO_PAD[92]
  PIN gfpga_pad_GPIO_PAD[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1375.600 51.880 1376.200 ;
    END
  END gfpga_pad_GPIO_PAD[93]
  PIN gfpga_pad_GPIO_PAD[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1437.480 51.880 1438.080 ;
    END
  END gfpga_pad_GPIO_PAD[94]
  PIN gfpga_pad_GPIO_PAD[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1499.360 51.880 1499.960 ;
    END
  END gfpga_pad_GPIO_PAD[95]
  PIN gfpga_pad_GPIO_PAD[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1925.450 1961.720 1925.730 1964.120 ;
    END
  END gfpga_pad_GPIO_PAD[9]
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2122.330 44.120 2122.610 46.520 ;
    END
  END reset
  PIN set
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2152.080 1931.840 2154.480 1932.440 ;
    END
  END set
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 2178.920 45.000 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 2203.920 20.000 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 105.000 92.485 2103.235 1914.035 ;
      LAYER met1 ;
        RECT 63.350 61.160 2139.190 1945.700 ;
      LAYER met2 ;
        RECT 63.370 1961.440 94.830 1961.720 ;
        RECT 95.670 1961.440 185.910 1961.720 ;
        RECT 186.750 1961.440 277.450 1961.720 ;
        RECT 278.290 1961.440 368.990 1961.720 ;
        RECT 369.830 1961.440 460.530 1961.720 ;
        RECT 461.370 1961.440 552.070 1961.720 ;
        RECT 552.910 1961.440 643.610 1961.720 ;
        RECT 644.450 1961.440 735.150 1961.720 ;
        RECT 735.990 1961.440 826.690 1961.720 ;
        RECT 827.530 1961.440 918.230 1961.720 ;
        RECT 919.070 1961.440 1009.770 1961.720 ;
        RECT 1010.610 1961.440 1101.310 1961.720 ;
        RECT 1102.150 1961.440 1192.850 1961.720 ;
        RECT 1193.690 1961.440 1284.390 1961.720 ;
        RECT 1285.230 1961.440 1375.930 1961.720 ;
        RECT 1376.770 1961.440 1467.470 1961.720 ;
        RECT 1468.310 1961.440 1559.010 1961.720 ;
        RECT 1559.850 1961.440 1650.550 1961.720 ;
        RECT 1651.390 1961.440 1742.090 1961.720 ;
        RECT 1742.930 1961.440 1833.630 1961.720 ;
        RECT 1834.470 1961.440 1925.170 1961.720 ;
        RECT 1926.010 1961.440 2016.710 1961.720 ;
        RECT 2017.550 1961.440 2108.250 1961.720 ;
        RECT 2109.090 1961.440 2139.170 1961.720 ;
        RECT 63.370 46.800 2139.170 1961.440 ;
        RECT 63.370 46.520 81.030 46.800 ;
        RECT 81.870 46.520 144.510 46.800 ;
        RECT 145.350 46.520 208.450 46.800 ;
        RECT 209.290 46.520 272.390 46.800 ;
        RECT 273.230 46.520 335.870 46.800 ;
        RECT 336.710 46.520 399.810 46.800 ;
        RECT 400.650 46.520 463.750 46.800 ;
        RECT 464.590 46.520 527.230 46.800 ;
        RECT 528.070 46.520 591.170 46.800 ;
        RECT 592.010 46.520 655.110 46.800 ;
        RECT 655.950 46.520 718.590 46.800 ;
        RECT 719.430 46.520 782.530 46.800 ;
        RECT 783.370 46.520 846.470 46.800 ;
        RECT 847.310 46.520 909.950 46.800 ;
        RECT 910.790 46.520 973.890 46.800 ;
        RECT 974.730 46.520 1037.830 46.800 ;
        RECT 1038.670 46.520 1101.310 46.800 ;
        RECT 1102.150 46.520 1165.250 46.800 ;
        RECT 1166.090 46.520 1229.190 46.800 ;
        RECT 1230.030 46.520 1292.670 46.800 ;
        RECT 1293.510 46.520 1356.610 46.800 ;
        RECT 1357.450 46.520 1420.550 46.800 ;
        RECT 1421.390 46.520 1484.030 46.800 ;
        RECT 1484.870 46.520 1547.970 46.800 ;
        RECT 1548.810 46.520 1611.910 46.800 ;
        RECT 1612.750 46.520 1675.390 46.800 ;
        RECT 1676.230 46.520 1739.330 46.800 ;
        RECT 1740.170 46.520 1803.270 46.800 ;
        RECT 1804.110 46.520 1866.750 46.800 ;
        RECT 1867.590 46.520 1930.690 46.800 ;
        RECT 1931.530 46.520 1994.630 46.800 ;
        RECT 1995.470 46.520 2058.110 46.800 ;
        RECT 2058.950 46.520 2122.050 46.800 ;
        RECT 2122.890 46.520 2139.170 46.800 ;
      LAYER met3 ;
        RECT 51.880 1933.520 2152.080 1945.905 ;
        RECT 52.280 1932.840 2152.080 1933.520 ;
        RECT 52.280 1932.120 2151.680 1932.840 ;
        RECT 51.880 1931.440 2151.680 1932.120 ;
        RECT 51.880 1871.640 2152.080 1931.440 ;
        RECT 52.280 1870.240 2152.080 1871.640 ;
        RECT 51.880 1868.920 2152.080 1870.240 ;
        RECT 51.880 1867.520 2151.680 1868.920 ;
        RECT 51.880 1809.760 2152.080 1867.520 ;
        RECT 52.280 1808.360 2152.080 1809.760 ;
        RECT 51.880 1805.000 2152.080 1808.360 ;
        RECT 51.880 1803.600 2151.680 1805.000 ;
        RECT 51.880 1747.880 2152.080 1803.600 ;
        RECT 52.280 1746.480 2152.080 1747.880 ;
        RECT 51.880 1741.080 2152.080 1746.480 ;
        RECT 51.880 1739.680 2151.680 1741.080 ;
        RECT 51.880 1686.000 2152.080 1739.680 ;
        RECT 52.280 1684.600 2152.080 1686.000 ;
        RECT 51.880 1677.160 2152.080 1684.600 ;
        RECT 51.880 1675.760 2151.680 1677.160 ;
        RECT 51.880 1624.120 2152.080 1675.760 ;
        RECT 52.280 1622.720 2152.080 1624.120 ;
        RECT 51.880 1613.240 2152.080 1622.720 ;
        RECT 51.880 1611.840 2151.680 1613.240 ;
        RECT 51.880 1562.240 2152.080 1611.840 ;
        RECT 52.280 1560.840 2152.080 1562.240 ;
        RECT 51.880 1549.320 2152.080 1560.840 ;
        RECT 51.880 1547.920 2151.680 1549.320 ;
        RECT 51.880 1500.360 2152.080 1547.920 ;
        RECT 52.280 1498.960 2152.080 1500.360 ;
        RECT 51.880 1484.720 2152.080 1498.960 ;
        RECT 51.880 1483.320 2151.680 1484.720 ;
        RECT 51.880 1438.480 2152.080 1483.320 ;
        RECT 52.280 1437.080 2152.080 1438.480 ;
        RECT 51.880 1420.800 2152.080 1437.080 ;
        RECT 51.880 1419.400 2151.680 1420.800 ;
        RECT 51.880 1376.600 2152.080 1419.400 ;
        RECT 52.280 1375.200 2152.080 1376.600 ;
        RECT 51.880 1356.880 2152.080 1375.200 ;
        RECT 51.880 1355.480 2151.680 1356.880 ;
        RECT 51.880 1314.040 2152.080 1355.480 ;
        RECT 52.280 1312.640 2152.080 1314.040 ;
        RECT 51.880 1292.960 2152.080 1312.640 ;
        RECT 51.880 1291.560 2151.680 1292.960 ;
        RECT 51.880 1252.160 2152.080 1291.560 ;
        RECT 52.280 1250.760 2152.080 1252.160 ;
        RECT 51.880 1229.040 2152.080 1250.760 ;
        RECT 51.880 1227.640 2151.680 1229.040 ;
        RECT 51.880 1190.280 2152.080 1227.640 ;
        RECT 52.280 1188.880 2152.080 1190.280 ;
        RECT 51.880 1165.120 2152.080 1188.880 ;
        RECT 51.880 1163.720 2151.680 1165.120 ;
        RECT 51.880 1128.400 2152.080 1163.720 ;
        RECT 52.280 1127.000 2152.080 1128.400 ;
        RECT 51.880 1101.200 2152.080 1127.000 ;
        RECT 51.880 1099.800 2151.680 1101.200 ;
        RECT 51.880 1066.520 2152.080 1099.800 ;
        RECT 52.280 1065.120 2152.080 1066.520 ;
        RECT 51.880 1037.280 2152.080 1065.120 ;
        RECT 51.880 1035.880 2151.680 1037.280 ;
        RECT 51.880 1004.640 2152.080 1035.880 ;
        RECT 52.280 1003.240 2152.080 1004.640 ;
        RECT 51.880 972.680 2152.080 1003.240 ;
        RECT 51.880 971.280 2151.680 972.680 ;
        RECT 51.880 942.760 2152.080 971.280 ;
        RECT 52.280 941.360 2152.080 942.760 ;
        RECT 51.880 908.760 2152.080 941.360 ;
        RECT 51.880 907.360 2151.680 908.760 ;
        RECT 51.880 880.880 2152.080 907.360 ;
        RECT 52.280 879.480 2152.080 880.880 ;
        RECT 51.880 844.840 2152.080 879.480 ;
        RECT 51.880 843.440 2151.680 844.840 ;
        RECT 51.880 819.000 2152.080 843.440 ;
        RECT 52.280 817.600 2152.080 819.000 ;
        RECT 51.880 780.920 2152.080 817.600 ;
        RECT 51.880 779.520 2151.680 780.920 ;
        RECT 51.880 757.120 2152.080 779.520 ;
        RECT 52.280 755.720 2152.080 757.120 ;
        RECT 51.880 717.000 2152.080 755.720 ;
        RECT 51.880 715.600 2151.680 717.000 ;
        RECT 51.880 694.560 2152.080 715.600 ;
        RECT 52.280 693.160 2152.080 694.560 ;
        RECT 51.880 653.080 2152.080 693.160 ;
        RECT 51.880 651.680 2151.680 653.080 ;
        RECT 51.880 632.680 2152.080 651.680 ;
        RECT 52.280 631.280 2152.080 632.680 ;
        RECT 51.880 589.160 2152.080 631.280 ;
        RECT 51.880 587.760 2151.680 589.160 ;
        RECT 51.880 570.800 2152.080 587.760 ;
        RECT 52.280 569.400 2152.080 570.800 ;
        RECT 51.880 524.560 2152.080 569.400 ;
        RECT 51.880 523.160 2151.680 524.560 ;
        RECT 51.880 508.920 2152.080 523.160 ;
        RECT 52.280 507.520 2152.080 508.920 ;
        RECT 51.880 460.640 2152.080 507.520 ;
        RECT 51.880 459.240 2151.680 460.640 ;
        RECT 51.880 447.040 2152.080 459.240 ;
        RECT 52.280 445.640 2152.080 447.040 ;
        RECT 51.880 396.720 2152.080 445.640 ;
        RECT 51.880 395.320 2151.680 396.720 ;
        RECT 51.880 385.160 2152.080 395.320 ;
        RECT 52.280 383.760 2152.080 385.160 ;
        RECT 51.880 332.800 2152.080 383.760 ;
        RECT 51.880 331.400 2151.680 332.800 ;
        RECT 51.880 323.280 2152.080 331.400 ;
        RECT 52.280 321.880 2152.080 323.280 ;
        RECT 51.880 268.880 2152.080 321.880 ;
        RECT 51.880 267.480 2151.680 268.880 ;
        RECT 51.880 261.400 2152.080 267.480 ;
        RECT 52.280 260.000 2152.080 261.400 ;
        RECT 51.880 204.960 2152.080 260.000 ;
        RECT 51.880 203.560 2151.680 204.960 ;
        RECT 51.880 199.520 2152.080 203.560 ;
        RECT 52.280 198.120 2152.080 199.520 ;
        RECT 51.880 141.040 2152.080 198.120 ;
        RECT 51.880 139.640 2151.680 141.040 ;
        RECT 51.880 137.640 2152.080 139.640 ;
        RECT 52.280 136.240 2152.080 137.640 ;
        RECT 51.880 77.120 2152.080 136.240 ;
        RECT 51.880 75.760 2151.680 77.120 ;
        RECT 52.280 75.720 2151.680 75.760 ;
        RECT 52.280 74.360 2152.080 75.720 ;
        RECT 51.880 60.615 2152.080 74.360 ;
      LAYER met4 ;
        RECT 0.000 0.000 2203.920 2005.840 ;
      LAYER met5 ;
        RECT 0.000 70.850 2203.920 2005.840 ;
  END
END fpga_top
END LIBRARY

