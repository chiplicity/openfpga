* NGSPICE file created from cbx_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt cbx_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_4_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_0_ top_grid_pin_10_ top_grid_pin_12_ top_grid_pin_14_
+ top_grid_pin_2_ top_grid_pin_4_ top_grid_pin_6_ top_grid_pin_8_ vpwr vgnd
XFILLER_10_317 vpwr vgnd scs8hd_fill_2
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_166 vpwr vgnd scs8hd_fill_2
XFILLER_9_148 vpwr vgnd scs8hd_fill_2
XFILLER_9_159 vgnd vpwr scs8hd_decap_3
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_170 vpwr vgnd scs8hd_fill_2
XFILLER_10_169 vpwr vgnd scs8hd_fill_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_6
XFILLER_2_335 vgnd vpwr scs8hd_fill_1
XFILLER_18_247 vpwr vgnd scs8hd_fill_2
XANTENNA__124__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vpwr vgnd scs8hd_fill_2
XFILLER_5_195 vpwr vgnd scs8hd_fill_2
XFILLER_17_291 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_4.LATCH_4_.latch data_in mem_bottom_ipin_4.LATCH_4_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_200_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__209__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_131_ _112_/A _133_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XANTENNA__110__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_44 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_242 vgnd vpwr scs8hd_decap_6
XFILLER_18_20 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_264 vgnd vpwr scs8hd_fill_1
X_114_ _140_/A _111_/X _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_224 vgnd vpwr scs8hd_fill_1
XFILLER_11_297 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_342 vgnd vpwr scs8hd_decap_12
XFILLER_6_290 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_6
XFILLER_16_389 vgnd vpwr scs8hd_decap_8
XANTENNA__116__B _111_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_282 vpwr vgnd scs8hd_fill_2
XFILLER_3_293 vpwr vgnd scs8hd_fill_2
XANTENNA__132__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_45 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_65 vgnd vpwr scs8hd_decap_8
XFILLER_0_274 vpwr vgnd scs8hd_fill_2
XFILLER_0_263 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _105_/A vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XFILLER_8_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.LATCH_0_.latch data_in mem_bottom_ipin_5.LATCH_0_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_189 vpwr vgnd scs8hd_fill_2
XFILLER_5_300 vpwr vgnd scs8hd_fill_2
XFILLER_9_127 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_108 vgnd vpwr scs8hd_decap_8
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_7.LATCH_3_.latch data_in mem_bottom_ipin_7.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_391 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XFILLER_15_229 vgnd vpwr scs8hd_decap_4
XFILLER_15_218 vpwr vgnd scs8hd_fill_2
X_130_ _129_/X _133_/B vgnd vpwr scs8hd_buf_1
XFILLER_2_122 vpwr vgnd scs8hd_fill_2
XANTENNA__110__D _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA__119__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_14_273 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
X_113_ _113_/A _140_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_276 vpwr vgnd scs8hd_fill_2
XFILLER_19_354 vgnd vpwr scs8hd_decap_12
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_16_346 vgnd vpwr scs8hd_decap_12
XFILLER_3_250 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__132__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_15_33 vpwr vgnd scs8hd_fill_2
XFILLER_15_22 vpwr vgnd scs8hd_fill_2
XFILLER_15_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_132 vgnd vpwr scs8hd_decap_12
XFILLER_16_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_165 vgnd vpwr scs8hd_decap_12
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XANTENNA__127__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_375 vgnd vpwr scs8hd_decap_4
XANTENNA__143__A _105_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _150_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_9_117 vpwr vgnd scs8hd_fill_2
XFILLER_5_378 vgnd vpwr scs8hd_fill_1
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_149 vgnd vpwr scs8hd_decap_4
XFILLER_12_23 vgnd vpwr scs8hd_decap_8
XFILLER_12_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_337 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _159_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__140__B _141_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_145 vgnd vpwr scs8hd_decap_4
XFILLER_2_112 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_252 vpwr vgnd scs8hd_fill_2
XANTENNA__119__C _119_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_285 vgnd vpwr scs8hd_decap_4
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__135__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__151__A _175_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_211 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _166_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_99 vgnd vpwr scs8hd_decap_8
X_112_ _112_/A _111_/X _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A _145_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_80 vpwr vgnd scs8hd_fill_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_6
XFILLER_4_218 vgnd vpwr scs8hd_decap_4
XFILLER_16_369 vpwr vgnd scs8hd_fill_2
XFILLER_16_358 vgnd vpwr scs8hd_decap_3
XFILLER_6_25 vpwr vgnd scs8hd_fill_2
XFILLER_6_58 vpwr vgnd scs8hd_fill_2
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_0_.latch data_in _160_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_380 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_13_317 vpwr vgnd scs8hd_fill_2
XFILLER_0_287 vgnd vpwr scs8hd_decap_4
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XFILLER_16_144 vgnd vpwr scs8hd_decap_8
XFILLER_0_298 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_188 vgnd vpwr scs8hd_decap_8
XFILLER_16_177 vgnd vpwr scs8hd_decap_8
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_354 vpwr vgnd scs8hd_fill_2
XFILLER_12_350 vpwr vgnd scs8hd_fill_2
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
XANTENNA__143__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_147 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_107 vpwr vgnd scs8hd_fill_2
XFILLER_5_313 vpwr vgnd scs8hd_fill_2
XFILLER_5_324 vgnd vpwr scs8hd_decap_4
XFILLER_5_335 vpwr vgnd scs8hd_fill_2
XFILLER_5_357 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_128 vpwr vgnd scs8hd_fill_2
XFILLER_2_349 vgnd vpwr scs8hd_decap_12
XFILLER_18_239 vgnd vpwr scs8hd_decap_8
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_1.LATCH_0_.latch data_in mem_bottom_ipin_1.LATCH_0_.latch/Q _178_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_143 vpwr vgnd scs8hd_fill_2
XANTENNA__149__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_404 vgnd vpwr scs8hd_decap_3
XFILLER_11_404 vgnd vpwr scs8hd_decap_3
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_3_.latch data_in mem_bottom_ipin_3.LATCH_3_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_69 vpwr vgnd scs8hd_fill_2
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__B _150_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _161_/A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
X_111_ _110_/X _111_/X vgnd vpwr scs8hd_buf_1
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_216 vpwr vgnd scs8hd_fill_2
XFILLER_11_234 vpwr vgnd scs8hd_fill_2
XFILLER_11_256 vpwr vgnd scs8hd_fill_2
XFILLER_19_367 vgnd vpwr scs8hd_decap_12
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_271 vpwr vgnd scs8hd_fill_2
XFILLER_1_70 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__072__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_7 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_392 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_79 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_244 vgnd vpwr scs8hd_fill_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_388 vgnd vpwr scs8hd_decap_8
XFILLER_12_384 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_38 vpwr vgnd scs8hd_fill_2
XFILLER_8_174 vgnd vpwr scs8hd_decap_3
XANTENNA__154__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_170 vgnd vpwr scs8hd_decap_8
XFILLER_12_181 vgnd vpwr scs8hd_fill_1
XANTENNA__170__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_317 vgnd vpwr scs8hd_decap_12
XANTENNA__080__A _080_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_177 vgnd vpwr scs8hd_decap_4
XFILLER_17_251 vpwr vgnd scs8hd_fill_2
XANTENNA__149__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_81 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_6.LATCH_2_.latch data_in mem_bottom_ipin_6.LATCH_2_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_158 vpwr vgnd scs8hd_fill_2
XFILLER_14_265 vgnd vpwr scs8hd_decap_6
XFILLER_9_48 vgnd vpwr scs8hd_fill_1
XFILLER_13_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_191 vgnd vpwr scs8hd_decap_4
XFILLER_9_280 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
X_110_ _163_/A address[4] address[3] _121_/A _110_/X vgnd vpwr scs8hd_or4_4
XFILLER_11_213 vpwr vgnd scs8hd_fill_2
XFILLER_19_302 vgnd vpwr scs8hd_decap_3
XFILLER_19_379 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_294 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__072__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_286 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XFILLER_3_297 vpwr vgnd scs8hd_fill_2
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_15_360 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA__083__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_278 vgnd vpwr scs8hd_fill_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_396 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__168__A _168_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_92 vgnd vpwr scs8hd_fill_1
XFILLER_13_138 vpwr vgnd scs8hd_fill_2
XANTENNA__078__A _077_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_304 vgnd vpwr scs8hd_fill_1
XFILLER_3_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _159_/A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__170__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_329 vgnd vpwr scs8hd_decap_6
XANTENNA__080__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_4
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XFILLER_1_351 vgnd vpwr scs8hd_decap_12
XANTENNA__165__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA__075__B _137_/B vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_126 vpwr vgnd scs8hd_fill_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_4
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__176__A _168_/A vgnd vpwr scs8hd_diode_2
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
X_169_ _104_/A _168_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_251 vpwr vgnd scs8hd_fill_2
XFILLER_10_291 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_328 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_17 vpwr vgnd scs8hd_fill_2
XFILLER_3_210 vpwr vgnd scs8hd_fill_2
XFILLER_3_265 vpwr vgnd scs8hd_fill_2
XANTENNA__157__C _157_/C vgnd vpwr scs8hd_diode_2
XANTENNA__173__B _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_37 vpwr vgnd scs8hd_fill_2
XFILLER_15_26 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__083__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vgnd vpwr scs8hd_fill_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_4
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _180_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_38 vgnd vpwr scs8hd_fill_1
XANTENNA__080__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__089__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_363 vgnd vpwr scs8hd_decap_3
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XANTENNA__075__C address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_7 vgnd vpwr scs8hd_fill_1
XFILLER_0_19 vgnd vpwr scs8hd_decap_12
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_289 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__176__B _172_/X vgnd vpwr scs8hd_diode_2
XANTENNA__192__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__086__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _082_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
X_168_ _168_/A _168_/B _168_/Y vgnd vpwr scs8hd_nor2_4
X_099_ _098_/X _113_/A vgnd vpwr scs8hd_buf_1
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XFILLER_1_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_5_.latch data_in mem_bottom_ipin_4.LATCH_5_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__097__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_29 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_60 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_4
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__C _157_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XFILLER_0_225 vpwr vgnd scs8hd_fill_2
XFILLER_16_104 vpwr vgnd scs8hd_fill_2
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_310 vgnd vpwr scs8hd_decap_4
XFILLER_12_365 vpwr vgnd scs8hd_fill_2
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_358 vgnd vpwr scs8hd_decap_4
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_391 vgnd vpwr scs8hd_decap_12
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_5_339 vgnd vpwr scs8hd_decap_12
XFILLER_4_361 vgnd vpwr scs8hd_decap_12
XANTENNA__179__B _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA__195__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_320 vpwr vgnd scs8hd_fill_2
XFILLER_5_114 vgnd vpwr scs8hd_decap_4
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_106 vgnd vpwr scs8hd_decap_6
XFILLER_14_224 vgnd vpwr scs8hd_decap_12
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.LATCH_1_.latch data_in mem_bottom_ipin_5.LATCH_1_.latch/Q _127_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_249 vgnd vpwr scs8hd_decap_12
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_238 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_098_ address[1] _090_/B address[0] _098_/X vgnd vpwr scs8hd_or3_4
X_167_ _175_/A _168_/B _167_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_ipin_7.LATCH_4_.latch data_in mem_bottom_ipin_7.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__097__B _105_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_363 vgnd vpwr scs8hd_decap_3
XANTENNA__198__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_190 vgnd vpwr scs8hd_decap_6
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_348 vgnd vpwr scs8hd_decap_4
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_388 vgnd vpwr scs8hd_decap_8
XFILLER_11_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vpwr vgnd scs8hd_fill_2
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XFILLER_7_381 vgnd vpwr scs8hd_decap_3
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XFILLER_16_71 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_185 vpwr vgnd scs8hd_fill_2
XFILLER_4_373 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ _162_/A mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_4_41 vgnd vpwr scs8hd_decap_6
XFILLER_4_85 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_236 vgnd vpwr scs8hd_decap_3
XFILLER_13_94 vpwr vgnd scs8hd_fill_2
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _149_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XFILLER_9_262 vgnd vpwr scs8hd_decap_4
XFILLER_9_284 vpwr vgnd scs8hd_fill_2
XFILLER_18_28 vgnd vpwr scs8hd_decap_3
XFILLER_11_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_306 vgnd vpwr scs8hd_decap_12
X_097_ _112_/A _105_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_276 vgnd vpwr scs8hd_decap_3
X_166_ _140_/A _168_/B _166_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_31 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_18_372 vgnd vpwr scs8hd_fill_1
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_73 vgnd vpwr scs8hd_decap_8
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_10_84 vgnd vpwr scs8hd_decap_8
X_149_ _112_/A _150_/B _149_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_18 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_249 vgnd vpwr scs8hd_fill_1
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_316 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _165_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_30 vpwr vgnd scs8hd_fill_2
XFILLER_13_109 vgnd vpwr scs8hd_decap_3
XFILLER_17_404 vgnd vpwr scs8hd_decap_3
XFILLER_8_135 vgnd vpwr scs8hd_fill_1
XFILLER_4_385 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_1_.latch data_in _159_/A _155_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_127 vgnd vpwr scs8hd_fill_1
XFILLER_17_267 vgnd vpwr scs8hd_decap_12
XFILLER_17_256 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_4
XFILLER_17_201 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_182 vpwr vgnd scs8hd_fill_2
XFILLER_4_75 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__100__A _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_318 vgnd vpwr scs8hd_decap_12
X_165_ _092_/A _168_/B _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_255 vgnd vpwr scs8hd_decap_4
XFILLER_6_266 vgnd vpwr scs8hd_decap_3
X_096_ _096_/A _105_/B vgnd vpwr scs8hd_buf_1
XFILLER_20_19 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_1.LATCH_1_.latch data_in mem_bottom_ipin_1.LATCH_1_.latch/Q _177_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_3_214 vgnd vpwr scs8hd_decap_3
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vpwr vgnd scs8hd_fill_2
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XFILLER_19_159 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _160_/A mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_15_376 vpwr vgnd scs8hd_fill_2
XFILLER_15_343 vpwr vgnd scs8hd_fill_2
XFILLER_15_310 vgnd vpwr scs8hd_fill_1
X_148_ _147_/X _150_/B vgnd vpwr scs8hd_buf_1
X_079_ _141_/A _180_/A _079_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_ipin_3.LATCH_4_.latch data_in mem_bottom_ipin_3.LATCH_4_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_328 vgnd vpwr scs8hd_decap_8
XFILLER_12_346 vpwr vgnd scs8hd_fill_2
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_309 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_84 vgnd vpwr scs8hd_decap_8
XFILLER_12_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_158 vgnd vpwr scs8hd_fill_1
XANTENNA__103__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_301 vpwr vgnd scs8hd_fill_2
XFILLER_5_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XFILLER_17_279 vgnd vpwr scs8hd_decap_12
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XFILLER_4_161 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _161_/Y mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_205 vpwr vgnd scs8hd_fill_2
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XFILLER_1_164 vpwr vgnd scs8hd_fill_2
XANTENNA__100__B _113_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_260 vpwr vgnd scs8hd_fill_2
XFILLER_9_297 vgnd vpwr scs8hd_decap_4
XFILLER_1_8 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__201__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_0_.latch data_in mem_bottom_ipin_4.LATCH_0_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_164_ _163_/X _168_/B vgnd vpwr scs8hd_buf_1
X_095_ _163_/A _137_/B _119_/C _077_/A _096_/A vgnd vpwr scs8hd_or4_4
XFILLER_6_201 vpwr vgnd scs8hd_fill_2
XFILLER_6_234 vgnd vpwr scs8hd_decap_6
XFILLER_10_230 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__111__A _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_22 vpwr vgnd scs8hd_fill_2
XFILLER_1_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_53 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_6.LATCH_3_.latch data_in mem_bottom_ipin_6.LATCH_3_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_399 vpwr vgnd scs8hd_fill_2
XFILLER_15_388 vpwr vgnd scs8hd_fill_2
XFILLER_15_322 vpwr vgnd scs8hd_fill_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_147_ _163_/A address[4] address[3] _157_/B _147_/X vgnd vpwr scs8hd_or4_4
X_078_ _077_/X _180_/A vgnd vpwr scs8hd_buf_1
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
XFILLER_0_229 vpwr vgnd scs8hd_fill_2
XFILLER_16_108 vgnd vpwr scs8hd_decap_4
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_369 vpwr vgnd scs8hd_fill_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_43 vpwr vgnd scs8hd_fill_2
XFILLER_11_380 vpwr vgnd scs8hd_fill_2
XFILLER_7_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_104 vgnd vpwr scs8hd_decap_12
XFILLER_12_100 vpwr vgnd scs8hd_fill_2
XFILLER_12_133 vgnd vpwr scs8hd_fill_1
XANTENNA__103__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_170 vpwr vgnd scs8hd_fill_2
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__204__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vgnd vpwr scs8hd_fill_1
XFILLER_1_379 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_75 vgnd vpwr scs8hd_decap_4
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
X_180_ _180_/A _113_/A _180_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_42 vpwr vgnd scs8hd_fill_2
XFILLER_1_143 vgnd vpwr scs8hd_decap_4
XFILLER_1_187 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_9_210 vpwr vgnd scs8hd_fill_2
XFILLER_9_232 vpwr vgnd scs8hd_fill_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_094_ address[3] _119_/C vgnd vpwr scs8hd_inv_8
X_163_ _163_/A address[4] address[3] _077_/A _163_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_224 vgnd vpwr scs8hd_decap_3
XFILLER_10_253 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_364 vgnd vpwr scs8hd_decap_8
XFILLER_1_45 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_7.LATCH_3_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_15_301 vpwr vgnd scs8hd_fill_2
XFILLER_15_356 vgnd vpwr scs8hd_decap_4
X_146_ _145_/X _157_/B vgnd vpwr scs8hd_buf_1
XANTENNA__122__A _121_/X vgnd vpwr scs8hd_diode_2
X_077_ _077_/A _129_/A _077_/X vgnd vpwr scs8hd_or2_4
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_308 vgnd vpwr scs8hd_decap_8
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_175 vgnd vpwr scs8hd_decap_6
XFILLER_15_164 vgnd vpwr scs8hd_decap_4
XPHY_6 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _159_/Y mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XFILLER_7_11 vpwr vgnd scs8hd_fill_2
XFILLER_7_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__117__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_392 vgnd vpwr scs8hd_decap_12
XFILLER_7_99 vgnd vpwr scs8hd_decap_3
X_129_ _129_/A _121_/A _129_/X vgnd vpwr scs8hd_or2_4
XFILLER_8_116 vpwr vgnd scs8hd_fill_2
XFILLER_8_138 vpwr vgnd scs8hd_fill_2
XFILLER_12_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_178 vgnd vpwr scs8hd_fill_1
XFILLER_12_189 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__114__B _111_/X vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_4
XFILLER_4_89 vgnd vpwr scs8hd_fill_1
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _154_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_21 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_4
XFILLER_13_284 vpwr vgnd scs8hd_fill_2
XFILLER_13_273 vgnd vpwr scs8hd_decap_3
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _145_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_266 vgnd vpwr scs8hd_fill_1
XANTENNA__125__A _141_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_162_ _162_/A _162_/Y vgnd vpwr scs8hd_inv_8
X_093_ _075_/A _163_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_265 vpwr vgnd scs8hd_fill_2
XFILLER_10_287 vpwr vgnd scs8hd_fill_2
XFILLER_1_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_291 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_22 vgnd vpwr scs8hd_decap_3
XFILLER_10_99 vgnd vpwr scs8hd_decap_3
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
X_145_ address[5] _145_/B _145_/X vgnd vpwr scs8hd_or2_4
XFILLER_2_283 vgnd vpwr scs8hd_decap_6
XFILLER_2_272 vgnd vpwr scs8hd_fill_1
X_076_ _075_/X _129_/A vgnd vpwr scs8hd_buf_1
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_209 vgnd vpwr scs8hd_decap_4
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_316 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vgnd vpwr scs8hd_decap_6
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
X_128_ _144_/A _124_/B _128_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _079_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__133__A _141_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B _111_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_216 vpwr vgnd scs8hd_fill_2
XFILLER_17_205 vgnd vpwr scs8hd_decap_8
XFILLER_9_404 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_6.LATCH_3_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_11 vgnd vpwr scs8hd_fill_1
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _141_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
X_161_ _161_/A _161_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
X_092_ _092_/A _112_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_299 vgnd vpwr scs8hd_decap_3
XFILLER_18_300 vgnd vpwr scs8hd_decap_8
XFILLER_18_377 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _162_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_45 vpwr vgnd scs8hd_fill_2
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
X_144_ _144_/A _141_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_075_ _075_/A _137_/B address[3] _075_/X vgnd vpwr scs8hd_or3_4
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_90 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_5.LATCH_2_.latch data_in mem_bottom_ipin_5.LATCH_2_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_328 vgnd vpwr scs8hd_decap_8
XFILLER_15_111 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
X_127_ _105_/A _124_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_321 vgnd vpwr scs8hd_decap_3
XFILLER_7_354 vpwr vgnd scs8hd_fill_2
XFILLER_7_376 vgnd vpwr scs8hd_decap_3
XFILLER_7_387 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _133_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_7.LATCH_5_.latch data_in mem_bottom_ipin_7.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_158 vgnd vpwr scs8hd_fill_1
XFILLER_20_180 vgnd vpwr scs8hd_decap_6
XFILLER_4_302 vgnd vpwr scs8hd_decap_8
XFILLER_4_313 vpwr vgnd scs8hd_fill_2
XFILLER_4_335 vgnd vpwr scs8hd_fill_1
XFILLER_8_129 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_327 vgnd vpwr scs8hd_decap_12
XFILLER_1_316 vpwr vgnd scs8hd_fill_2
XFILLER_4_58 vgnd vpwr scs8hd_decap_6
XFILLER_4_132 vpwr vgnd scs8hd_fill_2
XFILLER_4_165 vgnd vpwr scs8hd_fill_1
XFILLER_16_261 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _112_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vpwr vgnd scs8hd_fill_2
XFILLER_13_231 vgnd vpwr scs8hd_decap_3
XFILLER_13_297 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_160_ _160_/A _160_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_205 vpwr vgnd scs8hd_fill_2
X_091_ _090_/X _092_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_245 vpwr vgnd scs8hd_fill_2
XFILLER_18_312 vgnd vpwr scs8hd_decap_12
XFILLER_1_26 vpwr vgnd scs8hd_fill_2
XFILLER_18_389 vgnd vpwr scs8hd_decap_8
XANTENNA__136__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_271 vpwr vgnd scs8hd_fill_2
XANTENNA__152__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_219 vpwr vgnd scs8hd_fill_2
XFILLER_10_57 vgnd vpwr scs8hd_fill_1
XFILLER_19_11 vpwr vgnd scs8hd_fill_2
XFILLER_15_326 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_074_ address[4] _137_/B vgnd vpwr scs8hd_inv_8
X_143_ _105_/A _141_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__147__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_373 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
X_126_ _142_/A _124_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_47 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_5.LATCH_3_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ _162_/Y mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_104 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _141_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_174 vgnd vpwr scs8hd_decap_4
X_109_ address[5] _145_/B _121_/A vgnd vpwr scs8hd_nand2_4
XFILLER_3_391 vgnd vpwr scs8hd_decap_12
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_270 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_306 vgnd vpwr scs8hd_fill_1
XFILLER_1_339 vgnd vpwr scs8hd_decap_12
XANTENNA__070__A _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_199 vpwr vgnd scs8hd_fill_2
XFILLER_16_273 vpwr vgnd scs8hd_fill_2
XFILLER_16_240 vgnd vpwr scs8hd_fill_1
XANTENNA__139__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_46 vpwr vgnd scs8hd_fill_2
XFILLER_1_158 vgnd vpwr scs8hd_decap_4
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_203 vpwr vgnd scs8hd_fill_2
XFILLER_9_214 vgnd vpwr scs8hd_decap_4
XFILLER_9_236 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_8_280 vpwr vgnd scs8hd_fill_2
XFILLER_8_291 vgnd vpwr scs8hd_decap_6
X_090_ address[1] _090_/B _157_/C _090_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_324 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__152__B _150_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_142_ _142_/A _141_/B _142_/Y vgnd vpwr scs8hd_nor2_4
X_073_ enable _075_/A vgnd vpwr scs8hd_inv_8
XFILLER_2_253 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XFILLER_18_110 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_81 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_385 vgnd vpwr scs8hd_decap_12
XANTENNA__073__A enable vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
X_125_ _141_/A _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_15 vpwr vgnd scs8hd_fill_2
XFILLER_7_26 vpwr vgnd scs8hd_fill_2
XFILLER_7_301 vpwr vgnd scs8hd_fill_2
XFILLER_11_363 vgnd vpwr scs8hd_fill_1
XANTENNA__158__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_35 vgnd vpwr scs8hd_decap_12
XANTENNA__068__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_79 vpwr vgnd scs8hd_fill_2
XFILLER_4_337 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_1.LATCH_2_.latch data_in mem_bottom_ipin_1.LATCH_2_.latch/Q _176_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_108_ address[6] _145_/B vgnd vpwr scs8hd_inv_8
XFILLER_7_120 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_282 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_3.LATCH_5_.latch data_in mem_bottom_ipin_3.LATCH_5_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_fill_1
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_4_178 vpwr vgnd scs8hd_fill_2
XANTENNA__155__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _077_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_25 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A _080_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_192 vpwr vgnd scs8hd_fill_2
XFILLER_0_181 vpwr vgnd scs8hd_fill_2
XFILLER_0_170 vpwr vgnd scs8hd_fill_2
XANTENNA__166__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_5_92 vgnd vpwr scs8hd_fill_1
XANTENNA__076__A _075_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_4.LATCH_3_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_229 vgnd vpwr scs8hd_decap_3
XFILLER_10_269 vgnd vpwr scs8hd_decap_6
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _160_/Y mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_295 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_339 vpwr vgnd scs8hd_fill_2
XFILLER_15_306 vgnd vpwr scs8hd_decap_4
X_141_ _141_/A _141_/B _141_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_232 vpwr vgnd scs8hd_fill_2
X_072_ address[5] address[6] _077_/A vgnd vpwr scs8hd_or2_4
XFILLER_18_122 vgnd vpwr scs8hd_decap_12
XFILLER_18_9 vgnd vpwr scs8hd_decap_8
XFILLER_18_199 vgnd vpwr scs8hd_decap_12
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_372 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__147__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__163__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_60 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_342 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_397 vgnd vpwr scs8hd_decap_6
XFILLER_15_136 vgnd vpwr scs8hd_decap_4
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
X_124_ _140_/A _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_335 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__158__B _157_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_1_.latch data_in mem_bottom_ipin_4.LATCH_1_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__174__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_47 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_349 vgnd vpwr scs8hd_decap_12
X_107_ _144_/A _105_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_161 vpwr vgnd scs8hd_fill_2
XFILLER_11_194 vpwr vgnd scs8hd_fill_2
XFILLER_3_360 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_4_.latch data_in mem_bottom_ipin_6.LATCH_4_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XFILLER_19_294 vgnd vpwr scs8hd_decap_8
XANTENNA__169__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_70 vgnd vpwr scs8hd_decap_3
XANTENNA__079__A _141_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XFILLER_4_168 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _161_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__155__C _157_/C vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_105 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_13_278 vgnd vpwr scs8hd_decap_4
XFILLER_13_256 vpwr vgnd scs8hd_fill_2
XFILLER_13_212 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_204 vpwr vgnd scs8hd_fill_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_4
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_18 vpwr vgnd scs8hd_fill_2
XFILLER_18_337 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_392 vgnd vpwr scs8hd_decap_12
XFILLER_17_381 vgnd vpwr scs8hd_decap_4
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
X_140_ _140_/A _141_/B _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ _175_/A _141_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_266 vgnd vpwr scs8hd_decap_6
XFILLER_18_134 vgnd vpwr scs8hd_decap_12
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_384 vpwr vgnd scs8hd_fill_2
XANTENNA__147__D _157_/B vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_354 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_7.LATCH_0_.latch data_in mem_bottom_ipin_7.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_358 vpwr vgnd scs8hd_fill_2
X_123_ _112_/A _124_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_376 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vgnd vpwr scs8hd_decap_8
XANTENNA__158__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_192 vpwr vgnd scs8hd_fill_2
XANTENNA__174__B _172_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_59 vgnd vpwr scs8hd_decap_12
XFILLER_12_129 vgnd vpwr scs8hd_decap_4
XFILLER_4_317 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
X_106_ _106_/A _144_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_184 vgnd vpwr scs8hd_fill_1
XANTENNA__169__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_3.LATCH_3_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__079__B _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_405 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _163_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_114 vgnd vpwr scs8hd_decap_3
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XFILLER_0_342 vgnd vpwr scs8hd_decap_12
XFILLER_0_331 vpwr vgnd scs8hd_fill_2
XFILLER_0_320 vgnd vpwr scs8hd_decap_8
XFILLER_16_287 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_0_ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_139 vpwr vgnd scs8hd_fill_2
XFILLER_8_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_290 vgnd vpwr scs8hd_decap_6
XFILLER_5_72 vgnd vpwr scs8hd_decap_3
XFILLER_6_209 vgnd vpwr scs8hd_decap_3
XFILLER_10_249 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_7.LATCH_4_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_349 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_242 vpwr vgnd scs8hd_fill_2
XFILLER_5_275 vgnd vpwr scs8hd_decap_4
XANTENNA__177__B _172_/X vgnd vpwr scs8hd_diode_2
XANTENNA__193__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _153_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ _069_/X _175_/A vgnd vpwr scs8hd_buf_1
XFILLER_18_146 vgnd vpwr scs8hd_decap_6
XFILLER_14_396 vgnd vpwr scs8hd_fill_1
XFILLER_14_341 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__163__D _077_/A vgnd vpwr scs8hd_diode_2
X_199_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_20_366 vgnd vpwr scs8hd_decap_6
XFILLER_20_311 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_315 vgnd vpwr scs8hd_decap_4
XFILLER_11_355 vpwr vgnd scs8hd_fill_2
X_122_ _121_/X _124_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_82 vgnd vpwr scs8hd_decap_4
XFILLER_11_93 vpwr vgnd scs8hd_fill_2
XFILLER_11_388 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_119 vgnd vpwr scs8hd_decap_4
XFILLER_4_329 vgnd vpwr scs8hd_decap_6
X_105_ _105_/A _105_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_7_145 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vpwr vgnd scs8hd_fill_2
XFILLER_7_178 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__095__B _137_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_354 vgnd vpwr scs8hd_decap_12
XFILLER_16_299 vgnd vpwr scs8hd_decap_12
XFILLER_16_244 vgnd vpwr scs8hd_decap_8
XANTENNA__196__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _180_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_1_129 vgnd vpwr scs8hd_fill_1
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_218 vgnd vpwr scs8hd_fill_1
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XFILLER_6_7 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_18 vpwr vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_2_279 vpwr vgnd scs8hd_fill_2
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_198_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_52 vgnd vpwr scs8hd_decap_4
XFILLER_20_323 vgnd vpwr scs8hd_decap_12
XANTENNA__098__B _090_/B vgnd vpwr scs8hd_diode_2
X_121_ _121_/A _121_/B _121_/X vgnd vpwr scs8hd_or2_4
XFILLER_11_301 vpwr vgnd scs8hd_fill_2
XFILLER_11_323 vpwr vgnd scs8hd_fill_2
XFILLER_11_334 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_371 vpwr vgnd scs8hd_fill_2
XFILLER_6_382 vpwr vgnd scs8hd_fill_2
XANTENNA__199__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _162_/Y vgnd vpwr
+ scs8hd_diode_2
X_104_ _104_/A _105_/A vgnd vpwr scs8hd_buf_1
Xmem_bottom_ipin_3.LATCH_0_.latch data_in mem_bottom_ipin_3.LATCH_0_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_113 vgnd vpwr scs8hd_decap_4
XFILLER_11_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_6.LATCH_4_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__095__C _119_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XFILLER_0_366 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_5.LATCH_3_.latch data_in mem_bottom_ipin_5.LATCH_3_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_29 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XFILLER_0_185 vgnd vpwr scs8hd_fill_1
XFILLER_0_130 vpwr vgnd scs8hd_fill_2
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_362 vpwr vgnd scs8hd_fill_2
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_332 vgnd vpwr scs8hd_decap_4
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_335 vgnd vpwr scs8hd_decap_6
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_380 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_107 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_120_ _119_/X _121_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_339 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_394 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
X_103_ _142_/A _105_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_3_320 vpwr vgnd scs8hd_fill_2
XFILLER_11_198 vpwr vgnd scs8hd_fill_2
XFILLER_19_254 vpwr vgnd scs8hd_fill_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_180 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__D _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_106 vgnd vpwr scs8hd_decap_8
XFILLER_4_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_50 vgnd vpwr scs8hd_decap_8
XFILLER_16_224 vgnd vpwr scs8hd_decap_12
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_94 vgnd vpwr scs8hd_fill_1
XFILLER_16_279 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_1.LATCH_3_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vgnd vpwr scs8hd_decap_4
XFILLER_5_20 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_10_208 vgnd vpwr scs8hd_decap_6
XFILLER_18_308 vgnd vpwr scs8hd_fill_1
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_14_73 vgnd vpwr scs8hd_decap_8
XFILLER_14_62 vgnd vpwr scs8hd_decap_8
XFILLER_5_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_234 vpwr vgnd scs8hd_fill_2
XFILLER_17_330 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _141_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_14_388 vgnd vpwr scs8hd_decap_8
XFILLER_14_355 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_196_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_5.LATCH_4_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_87 vgnd vpwr scs8hd_fill_1
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_392 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_41 vgnd vpwr scs8hd_fill_1
XFILLER_2_3 vgnd vpwr scs8hd_decap_3
XFILLER_11_74 vpwr vgnd scs8hd_fill_2
XFILLER_19_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
X_179_ _180_/A _092_/A _179_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_340 vgnd vpwr scs8hd_decap_3
XFILLER_10_380 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_19 vgnd vpwr scs8hd_decap_12
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_102_ _168_/A _142_/A vgnd vpwr scs8hd_buf_1
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_75 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_335 vgnd vpwr scs8hd_decap_6
XFILLER_0_302 vgnd vpwr scs8hd_fill_1
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_16_236 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_280 vpwr vgnd scs8hd_fill_2
XFILLER_5_405 vpwr vgnd scs8hd_fill_2
XFILLER_0_187 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_3_.latch data_in mem_bottom_ipin_1.LATCH_3_.latch/Q _175_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_243 vgnd vpwr scs8hd_decap_3
XFILLER_8_276 vpwr vgnd scs8hd_fill_2
XFILLER_12_272 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_43 vgnd vpwr scs8hd_decap_4
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_279 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__101__B _105_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_2_249 vpwr vgnd scs8hd_fill_2
XFILLER_2_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_14_345 vgnd vpwr scs8hd_fill_1
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_195_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_77 vpwr vgnd scs8hd_fill_2
XFILLER_1_293 vpwr vgnd scs8hd_fill_2
XFILLER_1_282 vpwr vgnd scs8hd_fill_2
XFILLER_1_260 vpwr vgnd scs8hd_fill_2
XFILLER_17_161 vgnd vpwr scs8hd_decap_12
XFILLER_20_304 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_359 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__107__A _144_/A vgnd vpwr scs8hd_diode_2
X_178_ _106_/A _172_/X _178_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_392 vgnd vpwr scs8hd_decap_4
XFILLER_20_156 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_101_ _141_/A _105_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_112 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
XFILLER_11_178 vgnd vpwr scs8hd_decap_3
XFILLER_7_149 vgnd vpwr scs8hd_decap_4
XFILLER_19_245 vgnd vpwr scs8hd_decap_6
XFILLER_8_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _119_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_2_.latch data_in mem_bottom_ipin_4.LATCH_2_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_4.LATCH_4_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__205__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_177 vpwr vgnd scs8hd_fill_2
XFILLER_0_166 vpwr vgnd scs8hd_fill_2
XFILLER_8_211 vgnd vpwr scs8hd_fill_1
XFILLER_12_262 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__115__A _141_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_255 vgnd vpwr scs8hd_decap_8
XFILLER_8_266 vgnd vpwr scs8hd_decap_3
XFILLER_5_88 vgnd vpwr scs8hd_decap_4
XFILLER_5_99 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_6.LATCH_5_.latch data_in mem_bottom_ipin_6.LATCH_5_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_97 vpwr vgnd scs8hd_fill_2
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XFILLER_17_354 vgnd vpwr scs8hd_fill_1
XFILLER_17_321 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_228 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _161_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_14_313 vpwr vgnd scs8hd_fill_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_194_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__112__B _111_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_fill_1
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_6
XFILLER_17_173 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_327 vpwr vgnd scs8hd_fill_2
XFILLER_11_21 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
XFILLER_14_110 vgnd vpwr scs8hd_decap_8
XANTENNA__107__B _105_/B vgnd vpwr scs8hd_diode_2
X_177_ _104_/A _172_/X _177_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__123__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_375 vgnd vpwr scs8hd_decap_4
XFILLER_6_386 vgnd vpwr scs8hd_decap_8
XFILLER_20_168 vgnd vpwr scs8hd_decap_12
XFILLER_9_180 vgnd vpwr scs8hd_decap_3
XFILLER_7_117 vgnd vpwr scs8hd_fill_1
X_100_ _105_/B _113_/A _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_157 vpwr vgnd scs8hd_fill_2
XANTENNA__208__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_301 vgnd vpwr scs8hd_decap_4
XFILLER_3_367 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_88 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_17_86 vgnd vpwr scs8hd_decap_8
XFILLER_3_142 vgnd vpwr scs8hd_decap_4
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_7.LATCH_1_.latch data_in mem_bottom_ipin_7.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_208 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_fill_1
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_285 vgnd vpwr scs8hd_decap_3
XFILLER_12_296 vgnd vpwr scs8hd_fill_1
XANTENNA__115__B _111_/X vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_43 vgnd vpwr scs8hd_decap_12
XFILLER_14_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_388 vpwr vgnd scs8hd_fill_2
XFILLER_17_377 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_270 vgnd vpwr scs8hd_decap_4
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
X_193_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XFILLER_2_46 vgnd vpwr scs8hd_decap_4
XFILLER_2_35 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_306 vgnd vpwr scs8hd_decap_6
XFILLER_11_339 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
XFILLER_14_188 vpwr vgnd scs8hd_fill_2
XFILLER_14_177 vpwr vgnd scs8hd_fill_2
X_176_ _168_/A _172_/X _176_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_354 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_3.LATCH_4_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_3 vgnd vpwr scs8hd_decap_6
XFILLER_3_313 vpwr vgnd scs8hd_fill_2
XFILLER_3_324 vgnd vpwr scs8hd_decap_12
XFILLER_3_379 vgnd vpwr scs8hd_decap_12
XFILLER_19_258 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _152_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_3
XANTENNA__118__B _111_/X vgnd vpwr scs8hd_diode_2
X_159_ _159_/A _159_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_184 vgnd vpwr scs8hd_decap_4
XFILLER_10_191 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_305 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_132 vgnd vpwr scs8hd_decap_4
XFILLER_15_250 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _129_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_bottom_ipin_7.LATCH_5_.latch/Q
+ mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_224 vpwr vgnd scs8hd_fill_2
XFILLER_8_235 vgnd vpwr scs8hd_decap_8
XANTENNA__131__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_24 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_88 vgnd vpwr scs8hd_decap_4
XFILLER_14_55 vgnd vpwr scs8hd_decap_4
XFILLER_5_238 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_367 vgnd vpwr scs8hd_decap_4
XFILLER_17_334 vgnd vpwr scs8hd_decap_12
XANTENNA__126__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_14_359 vgnd vpwr scs8hd_decap_4
XFILLER_14_337 vpwr vgnd scs8hd_fill_2
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _179_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_21 vgnd vpwr scs8hd_decap_3
X_192_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_341 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_78 vpwr vgnd scs8hd_fill_2
XFILLER_11_89 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_6
X_175_ _175_/A _172_/X _175_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_311 vgnd vpwr scs8hd_decap_4
XFILLER_10_351 vgnd vpwr scs8hd_fill_1
XFILLER_20_137 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_336 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_089_ address[2] _090_/B vgnd vpwr scs8hd_inv_8
X_158_ _129_/A _157_/B address[0] _158_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_163 vgnd vpwr scs8hd_decap_3
XANTENNA__134__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _140_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_12_ vgnd vpwr scs8hd_inv_1
XFILLER_17_22 vpwr vgnd scs8hd_fill_2
XFILLER_17_11 vpwr vgnd scs8hd_fill_2
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XFILLER_15_284 vpwr vgnd scs8hd_fill_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__129__B _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_47 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_3.LATCH_1_.latch data_in mem_bottom_ipin_3.LATCH_1_.latch/Q _105_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_280 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_5_217 vpwr vgnd scs8hd_fill_2
XFILLER_5_228 vgnd vpwr scs8hd_decap_4
XFILLER_17_346 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _141_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.LATCH_4_.latch data_in mem_bottom_ipin_5.LATCH_4_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_209 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_14_327 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_15 vpwr vgnd scs8hd_fill_2
XFILLER_1_297 vpwr vgnd scs8hd_fill_2
XFILLER_1_286 vpwr vgnd scs8hd_fill_2
XFILLER_1_264 vpwr vgnd scs8hd_fill_2
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
XFILLER_13_393 vgnd vpwr scs8hd_decap_12
XFILLER_13_382 vpwr vgnd scs8hd_fill_2
XANTENNA__137__B _137_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _105_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_14_135 vgnd vpwr scs8hd_fill_1
X_174_ _113_/A _172_/X _174_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_345 vgnd vpwr scs8hd_decap_6
XFILLER_10_363 vgnd vpwr scs8hd_decap_4
XFILLER_10_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _147_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_149 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_bottom_ipin_6.LATCH_5_.latch/Q
+ mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_116 vgnd vpwr scs8hd_decap_6
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XFILLER_3_348 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_157_ _129_/A _157_/B _157_/C _157_/Y vgnd vpwr scs8hd_nor3_4
X_088_ _180_/A _106_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_263 vpwr vgnd scs8hd_fill_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
X_209_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_90 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A _175_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_0_.latch data_in mem_bottom_ipin_6.LATCH_0_.latch/Q _136_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_266 vgnd vpwr scs8hd_decap_6
XANTENNA__156__A _121_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_358 vpwr vgnd scs8hd_fill_2
XFILLER_17_303 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_14_317 vgnd vpwr scs8hd_fill_1
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_210 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_155 vgnd vpwr scs8hd_decap_3
XFILLER_13_350 vpwr vgnd scs8hd_fill_2
XANTENNA__137__C _119_/C vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_310 vgnd vpwr scs8hd_decap_3
XFILLER_9_376 vpwr vgnd scs8hd_fill_2
XFILLER_11_25 vpwr vgnd scs8hd_fill_2
XFILLER_14_169 vgnd vpwr scs8hd_decap_8
XFILLER_14_158 vpwr vgnd scs8hd_fill_2
X_173_ _092_/A _172_/X _173_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_324 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_92 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _160_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__074__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
X_156_ _121_/B _157_/B address[0] _156_/Y vgnd vpwr scs8hd_nor3_4
X_087_ _086_/X _106_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _080_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_209 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_1.LATCH_4_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_113 vgnd vpwr scs8hd_decap_3
XFILLER_3_146 vgnd vpwr scs8hd_fill_1
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_297 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
X_139_ _112_/A _141_/B _139_/Y vgnd vpwr scs8hd_nor2_4
X_208_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_190 vpwr vgnd scs8hd_fill_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_8_205 vgnd vpwr scs8hd_decap_6
XFILLER_12_223 vpwr vgnd scs8hd_fill_2
XFILLER_5_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _157_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_260 vgnd vpwr scs8hd_decap_3
XANTENNA__082__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_208 vpwr vgnd scs8hd_fill_2
XFILLER_1_403 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _186_/HI mem_bottom_ipin_5.LATCH_5_.latch/Q
+ mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_241 vgnd vpwr scs8hd_decap_4
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XFILLER_4_285 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_81 vpwr vgnd scs8hd_fill_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3 vgnd vpwr scs8hd_decap_4
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XANTENNA__137__D _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_90 vpwr vgnd scs8hd_fill_2
XFILLER_13_362 vpwr vgnd scs8hd_fill_2
XFILLER_9_388 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_1.LATCH_4_.latch data_in mem_bottom_ipin_1.LATCH_4_.latch/Q _174_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_37 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_172_ _172_/A _172_/X vgnd vpwr scs8hd_buf_1
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_118 vgnd vpwr scs8hd_decap_6
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__090__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_086_ address[1] address[2] address[0] _086_/X vgnd vpwr scs8hd_or3_4
X_155_ _121_/B _157_/B _157_/C _155_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_10_173 vgnd vpwr scs8hd_decap_4
XFILLER_2_361 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_2.LATCH_0_.latch data_in _162_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_309 vgnd vpwr scs8hd_fill_1
XANTENNA__069__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_58 vgnd vpwr scs8hd_decap_3
XANTENNA__085__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_158 vpwr vgnd scs8hd_fill_2
X_207_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_138_ _137_/X _141_/B vgnd vpwr scs8hd_buf_1
X_069_ _080_/A address[2] _157_/C _069_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_228 vpwr vgnd scs8hd_fill_2
XFILLER_12_202 vpwr vgnd scs8hd_fill_2
XFILLER_5_39 vpwr vgnd scs8hd_fill_2
XANTENNA__156__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _168_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_253 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _168_/B vgnd vpwr scs8hd_diode_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _129_/A vgnd vpwr scs8hd_diode_2
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_256 vpwr vgnd scs8hd_fill_2
XFILLER_17_135 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_4.LATCH_3_.latch data_in mem_bottom_ipin_4.LATCH_3_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_301 vgnd vpwr scs8hd_fill_1
XFILLER_9_345 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _106_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__088__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_127 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _077_/A _121_/B _172_/A vgnd vpwr scs8hd_or2_4
XFILLER_10_344 vgnd vpwr scs8hd_decap_4
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_131 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vgnd vpwr scs8hd_decap_3
XANTENNA__180__B _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_370 vpwr vgnd scs8hd_fill_2
XFILLER_5_381 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_108 vpwr vgnd scs8hd_fill_2
XANTENNA__090__B _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_15_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_085_ _180_/A _104_/A _085_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
X_154_ _144_/A _150_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_373 vgnd vpwr scs8hd_decap_12
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_252 vgnd vpwr scs8hd_decap_8
XANTENNA__175__B _172_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_26 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__069__C _157_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _185_/HI mem_bottom_ipin_4.LATCH_5_.latch/Q
+ mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__B _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_206_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_137_ _163_/A _137_/B _119_/C _121_/A _137_/X vgnd vpwr scs8hd_or4_4
X_068_ address[0] _157_/C vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_107 vgnd vpwr scs8hd_decap_6
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_280 vgnd vpwr scs8hd_decap_12
XFILLER_12_258 vpwr vgnd scs8hd_fill_2
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_7_284 vpwr vgnd scs8hd_fill_2
XFILLER_11_280 vpwr vgnd scs8hd_fill_2
XFILLER_19_391 vgnd vpwr scs8hd_decap_12
XFILLER_17_317 vpwr vgnd scs8hd_fill_2
XFILLER_17_306 vgnd vpwr scs8hd_decap_8
XFILLER_4_210 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_ipin_7.LATCH_2_.latch data_in mem_bottom_ipin_7.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_14_309 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XFILLER_2_19 vpwr vgnd scs8hd_fill_2
XFILLER_1_268 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_147 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_331 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__178__B _172_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _106_/A vgnd vpwr scs8hd_diode_2
X_170_ _106_/A _168_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_121 vgnd vpwr scs8hd_fill_1
XFILLER_5_360 vpwr vgnd scs8hd_fill_2
XFILLER_5_393 vgnd vpwr scs8hd_decap_12
XFILLER_3_95 vgnd vpwr scs8hd_fill_1
XANTENNA__090__C _157_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _098_/X vgnd vpwr scs8hd_diode_2
X_153_ _105_/A _150_/B _153_/Y vgnd vpwr scs8hd_nor2_4
X_084_ _083_/X _104_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_168 vgnd vpwr scs8hd_decap_3
XFILLER_12_71 vgnd vpwr scs8hd_decap_4
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_385 vgnd vpwr scs8hd_decap_12
XFILLER_17_38 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_105 vpwr vgnd scs8hd_fill_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_267 vpwr vgnd scs8hd_fill_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_3
XFILLER_15_201 vpwr vgnd scs8hd_fill_2
X_205_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_136_ _144_/A _133_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_171 vpwr vgnd scs8hd_fill_2
X_067_ address[1] _080_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_74 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_292 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_119_ _163_/A address[4] _119_/C _119_/X vgnd vpwr scs8hd_or3_4
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _151_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__197__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_222 vgnd vpwr scs8hd_fill_1
XFILLER_4_266 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _159_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_16 vgnd vpwr scs8hd_decap_3
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_1_225 vpwr vgnd scs8hd_fill_2
XFILLER_13_376 vgnd vpwr scs8hd_decap_4
XFILLER_13_354 vpwr vgnd scs8hd_fill_2
XFILLER_13_321 vpwr vgnd scs8hd_fill_2
XFILLER_9_358 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _184_/HI mem_bottom_ipin_3.LATCH_5_.latch/Q
+ mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_313 vpwr vgnd scs8hd_fill_2
XFILLER_10_324 vgnd vpwr scs8hd_decap_12
XFILLER_6_328 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_13_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_111 vgnd vpwr scs8hd_decap_4
XFILLER_9_144 vpwr vgnd scs8hd_fill_2
XFILLER_9_155 vpwr vgnd scs8hd_fill_2
XFILLER_9_199 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_309 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
X_083_ address[1] address[2] _157_/C _083_/X vgnd vpwr scs8hd_or3_4
X_152_ _142_/A _150_/B _152_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_132 vpwr vgnd scs8hd_fill_2
XFILLER_10_165 vpwr vgnd scs8hd_fill_2
XFILLER_10_187 vpwr vgnd scs8hd_fill_2
XFILLER_12_50 vgnd vpwr scs8hd_decap_8
XFILLER_18_276 vgnd vpwr scs8hd_decap_12
XFILLER_5_191 vpwr vgnd scs8hd_fill_2
X_204_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_135_ _105_/A _133_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_194 vpwr vgnd scs8hd_fill_2
XFILLER_9_51 vgnd vpwr scs8hd_decap_4
XFILLER_9_84 vgnd vpwr scs8hd_decap_4
XFILLER_12_227 vgnd vpwr scs8hd_decap_3
XFILLER_18_93 vgnd vpwr scs8hd_decap_4
XFILLER_7_220 vgnd vpwr scs8hd_decap_4
XFILLER_11_260 vgnd vpwr scs8hd_decap_4
XFILLER_7_297 vpwr vgnd scs8hd_fill_2
X_118_ _144_/A _111_/X _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_94 vgnd vpwr scs8hd_decap_12
XFILLER_4_256 vgnd vpwr scs8hd_fill_1
XFILLER_4_289 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_85 vgnd vpwr scs8hd_decap_6
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_15_94 vpwr vgnd scs8hd_fill_2
XFILLER_15_83 vpwr vgnd scs8hd_fill_2
XFILLER_9_304 vgnd vpwr scs8hd_fill_1
XFILLER_9_326 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_270 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_307 vpwr vgnd scs8hd_fill_2
XFILLER_10_369 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_2_.latch data_in mem_bottom_ipin_3.LATCH_2_.latch/Q _103_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_9_123 vgnd vpwr scs8hd_fill_1
XFILLER_3_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_42 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_5.LATCH_5_.latch data_in mem_bottom_ipin_5.LATCH_5_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_082_ _180_/A _168_/A _082_/Y vgnd vpwr scs8hd_nor2_4
X_151_ _175_/A _150_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_104 vpwr vgnd scs8hd_fill_2
XFILLER_10_111 vgnd vpwr scs8hd_decap_8
XFILLER_10_177 vgnd vpwr scs8hd_fill_1
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XFILLER_18_288 vgnd vpwr scs8hd_decap_12
XFILLER_18_211 vgnd vpwr scs8hd_decap_3
XFILLER_17_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_225 vpwr vgnd scs8hd_fill_2
XFILLER_15_214 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_203_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
X_134_ _142_/A _133_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_151 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vgnd vpwr scs8hd_decap_6
XFILLER_12_239 vgnd vpwr scs8hd_decap_6
XFILLER_20_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _183_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_7_265 vpwr vgnd scs8hd_fill_2
X_117_ _105_/A _111_/X _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_320 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_75 vgnd vpwr scs8hd_decap_4
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_17_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_73 vgnd vpwr scs8hd_decap_3
XFILLER_13_301 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _168_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_1_.latch data_in mem_bottom_ipin_6.LATCH_1_.latch/Q _135_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_371 vpwr vgnd scs8hd_fill_2
XFILLER_10_337 vpwr vgnd scs8hd_fill_2
XFILLER_10_348 vgnd vpwr scs8hd_fill_1
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_5_374 vgnd vpwr scs8hd_decap_4
XFILLER_3_21 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_150_ _140_/A _150_/B _150_/Y vgnd vpwr scs8hd_nor2_4
X_081_ _080_/X _168_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_300 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_116 vgnd vpwr scs8hd_fill_1
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_12_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__200__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_202_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_7_403 vgnd vpwr scs8hd_decap_4
X_133_ _141_/A _133_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_130 vgnd vpwr scs8hd_decap_6
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_11 vgnd vpwr scs8hd_fill_1
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_292 vgnd vpwr scs8hd_decap_6
XFILLER_20_273 vgnd vpwr scs8hd_decap_6
XFILLER_12_218 vgnd vpwr scs8hd_decap_3
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_284 vpwr vgnd scs8hd_fill_2
X_116_ _142_/A _111_/X _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _160_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_63 vgnd vpwr scs8hd_decap_12
XFILLER_4_225 vgnd vpwr scs8hd_decap_3
XFILLER_4_247 vgnd vpwr scs8hd_decap_6
XFILLER_16_332 vgnd vpwr scs8hd_decap_4
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
XFILLER_16_365 vpwr vgnd scs8hd_fill_2
XFILLER_6_21 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_1_206 vpwr vgnd scs8hd_fill_2
XFILLER_9_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_41 vgnd vpwr scs8hd_decap_12
XFILLER_13_335 vpwr vgnd scs8hd_fill_2
XFILLER_9_306 vpwr vgnd scs8hd_fill_2
XFILLER_0_294 vpwr vgnd scs8hd_fill_2
XFILLER_0_283 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__203__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_143 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vgnd vpwr scs8hd_decap_4
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_320 vpwr vgnd scs8hd_fill_2
XFILLER_5_331 vpwr vgnd scs8hd_fill_2
XFILLER_5_353 vgnd vpwr scs8hd_decap_4
XFILLER_5_364 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _182_/HI mem_bottom_ipin_1.LATCH_5_.latch/Q
+ mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_080_ _080_/A address[2] address[0] _080_/X vgnd vpwr scs8hd_or3_4
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XFILLER_6_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__108__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_109 vpwr vgnd scs8hd_fill_2
X_201_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
Xmem_bottom_ipin_1.LATCH_5_.latch data_in mem_bottom_ipin_1.LATCH_5_.latch/Q _173_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_132_ _140_/A _133_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_175 vgnd vpwr scs8hd_decap_4
XANTENNA__110__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_56 vgnd vpwr scs8hd_decap_4
XFILLER_0_78 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_9_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_230 vgnd vpwr scs8hd_decap_12
XFILLER_11_230 vpwr vgnd scs8hd_fill_2
XANTENNA__105__B _105_/B vgnd vpwr scs8hd_diode_2
X_115_ _141_/A _111_/X _115_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_201 vpwr vgnd scs8hd_fill_2
XFILLER_7_256 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_330 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_1_.latch data_in _161_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__206__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_75 vgnd vpwr scs8hd_decap_12
XFILLER_16_377 vgnd vpwr scs8hd_decap_8
XANTENNA__116__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_229 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vgnd vpwr scs8hd_decap_8
XFILLER_13_358 vpwr vgnd scs8hd_fill_2
XFILLER_13_325 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_240 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

