magic
tech sky130A
magscale 1 2
timestamp 1606930212
<< locali >>
rect 15393 7191 15427 7293
rect 15117 3383 15151 3689
rect 19257 3451 19291 3689
rect 14381 2907 14415 3145
rect 16037 2975 16071 3145
<< viali >>
rect 20729 20009 20763 20043
rect 20545 19873 20579 19907
rect 20177 19465 20211 19499
rect 16497 19261 16531 19295
rect 18337 19261 18371 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 16681 19125 16715 19159
rect 18521 19125 18555 19159
rect 20729 19125 20763 19159
rect 9965 18853 9999 18887
rect 15945 18853 15979 18887
rect 17877 18853 17911 18887
rect 19901 18853 19935 18887
rect 9689 18785 9723 18819
rect 12081 18785 12115 18819
rect 15669 18785 15703 18819
rect 17601 18785 17635 18819
rect 19625 18785 19659 18819
rect 12357 18717 12391 18751
rect 20177 18377 20211 18411
rect 20729 18377 20763 18411
rect 7757 18173 7791 18207
rect 19999 18173 20033 18207
rect 20545 18173 20579 18207
rect 8033 18105 8067 18139
rect 15485 17833 15519 17867
rect 20453 17833 20487 17867
rect 11437 17697 11471 17731
rect 15301 17697 15335 17731
rect 20269 17697 20303 17731
rect 11713 17629 11747 17663
rect 20177 17289 20211 17323
rect 20729 17289 20763 17323
rect 14473 17153 14507 17187
rect 14197 17085 14231 17119
rect 19993 17085 20027 17119
rect 20545 17085 20579 17119
rect 17325 16677 17359 16711
rect 19901 16677 19935 16711
rect 17049 16609 17083 16643
rect 19625 16609 19659 16643
rect 20177 16201 20211 16235
rect 20729 16201 20763 16235
rect 19993 15997 20027 16031
rect 20545 15997 20579 16031
rect 20453 15657 20487 15691
rect 14197 15589 14231 15623
rect 11805 15521 11839 15555
rect 13921 15521 13955 15555
rect 20269 15521 20303 15555
rect 12081 15453 12115 15487
rect 20729 15113 20763 15147
rect 9597 14909 9631 14943
rect 20545 14909 20579 14943
rect 9873 14841 9907 14875
rect 19901 14569 19935 14603
rect 20453 14569 20487 14603
rect 8401 14433 8435 14467
rect 19717 14433 19751 14467
rect 20269 14433 20303 14467
rect 8677 14365 8711 14399
rect 17509 14025 17543 14059
rect 19441 14025 19475 14059
rect 11069 13889 11103 13923
rect 20177 13889 20211 13923
rect 10793 13821 10827 13855
rect 16129 13821 16163 13855
rect 16396 13821 16430 13855
rect 19257 13821 19291 13855
rect 19993 13821 20027 13855
rect 19257 13481 19291 13515
rect 19901 13413 19935 13447
rect 19073 13345 19107 13379
rect 19625 13345 19659 13379
rect 15117 12937 15151 12971
rect 16957 12937 16991 12971
rect 19257 12937 19291 12971
rect 15669 12801 15703 12835
rect 17601 12801 17635 12835
rect 19901 12801 19935 12835
rect 19073 12733 19107 12767
rect 19625 12733 19659 12767
rect 20361 12733 20395 12767
rect 17417 12665 17451 12699
rect 20637 12665 20671 12699
rect 15485 12597 15519 12631
rect 15577 12597 15611 12631
rect 17325 12597 17359 12631
rect 15393 12393 15427 12427
rect 17325 12393 17359 12427
rect 20453 12393 20487 12427
rect 13522 12325 13556 12359
rect 17846 12325 17880 12359
rect 19717 12325 19751 12359
rect 13277 12257 13311 12291
rect 15945 12257 15979 12291
rect 16212 12257 16246 12291
rect 19441 12257 19475 12291
rect 20269 12257 20303 12291
rect 17601 12189 17635 12223
rect 14657 12053 14691 12087
rect 18981 12053 19015 12087
rect 15117 11849 15151 11883
rect 16773 11849 16807 11883
rect 13369 11713 13403 11747
rect 15393 11713 15427 11747
rect 17509 11713 17543 11747
rect 20729 11713 20763 11747
rect 20821 11713 20855 11747
rect 13093 11645 13127 11679
rect 13737 11645 13771 11679
rect 15660 11645 15694 11679
rect 18061 11645 18095 11679
rect 18620 11645 18654 11679
rect 18880 11645 18914 11679
rect 14004 11577 14038 11611
rect 12725 11509 12759 11543
rect 13185 11509 13219 11543
rect 18245 11509 18279 11543
rect 19993 11509 20027 11543
rect 20269 11509 20303 11543
rect 20637 11509 20671 11543
rect 14105 11305 14139 11339
rect 15301 11305 15335 11339
rect 15761 11305 15795 11339
rect 18705 11305 18739 11339
rect 20545 11305 20579 11339
rect 15669 11237 15703 11271
rect 16129 11237 16163 11271
rect 19432 11237 19466 11271
rect 12716 11169 12750 11203
rect 16497 11169 16531 11203
rect 17132 11169 17166 11203
rect 12449 11101 12483 11135
rect 15853 11101 15887 11135
rect 16865 11101 16899 11135
rect 19165 11101 19199 11135
rect 13829 11033 13863 11067
rect 16313 10965 16347 10999
rect 18245 10965 18279 10999
rect 15393 10761 15427 10795
rect 19073 10693 19107 10727
rect 16037 10625 16071 10659
rect 17049 10625 17083 10659
rect 18613 10625 18647 10659
rect 19717 10625 19751 10659
rect 20545 10625 20579 10659
rect 20637 10625 20671 10659
rect 12449 10557 12483 10591
rect 18429 10557 18463 10591
rect 19441 10557 19475 10591
rect 19533 10557 19567 10591
rect 12725 10489 12759 10523
rect 15853 10489 15887 10523
rect 18521 10489 18555 10523
rect 15761 10421 15795 10455
rect 16497 10421 16531 10455
rect 16865 10421 16899 10455
rect 16957 10421 16991 10455
rect 18061 10421 18095 10455
rect 20085 10421 20119 10455
rect 20453 10421 20487 10455
rect 13277 10217 13311 10251
rect 16957 10217 16991 10251
rect 17868 10149 17902 10183
rect 13645 10081 13679 10115
rect 15301 10081 15335 10115
rect 15568 10081 15602 10115
rect 19625 10081 19659 10115
rect 19717 10081 19751 10115
rect 20269 10081 20303 10115
rect 13737 10013 13771 10047
rect 13829 10013 13863 10047
rect 17601 10013 17635 10047
rect 19809 10013 19843 10047
rect 18981 9945 19015 9979
rect 16681 9877 16715 9911
rect 19257 9877 19291 9911
rect 20453 9877 20487 9911
rect 11069 9605 11103 9639
rect 11621 9537 11655 9571
rect 13001 9537 13035 9571
rect 17509 9537 17543 9571
rect 10977 9469 11011 9503
rect 13461 9469 13495 9503
rect 13728 9469 13762 9503
rect 15393 9469 15427 9503
rect 15660 9469 15694 9503
rect 18429 9469 18463 9503
rect 18696 9469 18730 9503
rect 20545 9469 20579 9503
rect 11437 9401 11471 9435
rect 10793 9333 10827 9367
rect 11529 9333 11563 9367
rect 14841 9333 14875 9367
rect 16773 9333 16807 9367
rect 19809 9333 19843 9367
rect 20729 9333 20763 9367
rect 9689 9129 9723 9163
rect 13829 9129 13863 9163
rect 15301 9129 15335 9163
rect 15761 9129 15795 9163
rect 16405 9129 16439 9163
rect 15669 9061 15703 9095
rect 19318 9061 19352 9095
rect 9137 8993 9171 9027
rect 10057 8993 10091 9027
rect 11060 8993 11094 9027
rect 12449 8993 12483 9027
rect 12716 8993 12750 9027
rect 13921 8993 13955 9027
rect 16773 8993 16807 9027
rect 19073 8993 19107 9027
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 10793 8925 10827 8959
rect 14105 8925 14139 8959
rect 15853 8925 15887 8959
rect 16865 8925 16899 8959
rect 17049 8925 17083 8959
rect 18613 8925 18647 8959
rect 12173 8789 12207 8823
rect 20453 8789 20487 8823
rect 11621 8585 11655 8619
rect 18613 8585 18647 8619
rect 21097 8585 21131 8619
rect 15577 8517 15611 8551
rect 11897 8449 11931 8483
rect 17509 8449 17543 8483
rect 19073 8449 19107 8483
rect 19257 8449 19291 8483
rect 8585 8381 8619 8415
rect 10241 8381 10275 8415
rect 13001 8381 13035 8415
rect 14841 8381 14875 8415
rect 15761 8381 15795 8415
rect 15853 8381 15887 8415
rect 18981 8381 19015 8415
rect 19717 8381 19751 8415
rect 19984 8381 20018 8415
rect 8852 8313 8886 8347
rect 10486 8313 10520 8347
rect 15117 8313 15151 8347
rect 16120 8313 16154 8347
rect 9965 8245 9999 8279
rect 14289 8245 14323 8279
rect 17233 8245 17267 8279
rect 9321 8041 9355 8075
rect 10609 8041 10643 8075
rect 13185 8041 13219 8075
rect 16221 8041 16255 8075
rect 19257 8041 19291 8075
rect 19809 8041 19843 8075
rect 10977 7973 11011 8007
rect 16589 7973 16623 8007
rect 16681 7973 16715 8007
rect 17509 7973 17543 8007
rect 19165 7973 19199 8007
rect 20913 7973 20947 8007
rect 7941 7905 7975 7939
rect 8208 7905 8242 7939
rect 12072 7905 12106 7939
rect 13461 7905 13495 7939
rect 13728 7905 13762 7939
rect 17233 7905 17267 7939
rect 20177 7905 20211 7939
rect 11069 7837 11103 7871
rect 11161 7837 11195 7871
rect 11805 7837 11839 7871
rect 16773 7837 16807 7871
rect 19349 7837 19383 7871
rect 20269 7837 20303 7871
rect 20453 7837 20487 7871
rect 14841 7701 14875 7735
rect 18797 7701 18831 7735
rect 11069 7497 11103 7531
rect 11345 7497 11379 7531
rect 12817 7497 12851 7531
rect 19625 7429 19659 7463
rect 11989 7361 12023 7395
rect 13369 7361 13403 7395
rect 13829 7361 13863 7395
rect 20269 7361 20303 7395
rect 11253 7293 11287 7327
rect 14096 7293 14130 7327
rect 15393 7293 15427 7327
rect 15485 7293 15519 7327
rect 17325 7293 17359 7327
rect 11713 7225 11747 7259
rect 13185 7225 13219 7259
rect 15730 7225 15764 7259
rect 19993 7225 20027 7259
rect 11805 7157 11839 7191
rect 13277 7157 13311 7191
rect 15209 7157 15243 7191
rect 15393 7157 15427 7191
rect 16865 7157 16899 7191
rect 17141 7157 17175 7191
rect 20085 7157 20119 7191
rect 12081 6953 12115 6987
rect 12357 6953 12391 6987
rect 14565 6953 14599 6987
rect 15301 6953 15335 6987
rect 13185 6885 13219 6919
rect 13277 6885 13311 6919
rect 10057 6817 10091 6851
rect 10968 6817 11002 6851
rect 15669 6817 15703 6851
rect 15761 6817 15795 6851
rect 16569 6817 16603 6851
rect 18236 6817 18270 6851
rect 19993 6817 20027 6851
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 10701 6749 10735 6783
rect 13369 6749 13403 6783
rect 14657 6749 14691 6783
rect 14841 6749 14875 6783
rect 15853 6749 15887 6783
rect 16313 6749 16347 6783
rect 17969 6749 18003 6783
rect 20085 6749 20119 6783
rect 20177 6749 20211 6783
rect 9689 6681 9723 6715
rect 12817 6681 12851 6715
rect 17693 6681 17727 6715
rect 19625 6681 19659 6715
rect 14197 6613 14231 6647
rect 19349 6613 19383 6647
rect 10885 6409 10919 6443
rect 11161 6409 11195 6443
rect 13461 6409 13495 6443
rect 15301 6409 15335 6443
rect 20361 6409 20395 6443
rect 11713 6273 11747 6307
rect 14105 6273 14139 6307
rect 14841 6273 14875 6307
rect 15853 6273 15887 6307
rect 16865 6273 16899 6307
rect 20913 6273 20947 6307
rect 7849 6205 7883 6239
rect 9505 6205 9539 6239
rect 9772 6205 9806 6239
rect 11621 6205 11655 6239
rect 16681 6205 16715 6239
rect 16773 6205 16807 6239
rect 18705 6205 18739 6239
rect 18972 6205 19006 6239
rect 20729 6205 20763 6239
rect 8116 6137 8150 6171
rect 15669 6137 15703 6171
rect 7389 6069 7423 6103
rect 9229 6069 9263 6103
rect 11529 6069 11563 6103
rect 13829 6069 13863 6103
rect 13921 6069 13955 6103
rect 15761 6069 15795 6103
rect 16313 6069 16347 6103
rect 18245 6069 18279 6103
rect 20085 6069 20119 6103
rect 20821 6069 20855 6103
rect 6653 5865 6687 5899
rect 9689 5865 9723 5899
rect 10425 5865 10459 5899
rect 14473 5865 14507 5899
rect 15301 5865 15335 5899
rect 16313 5865 16347 5899
rect 16773 5865 16807 5899
rect 19257 5865 19291 5899
rect 6745 5797 6779 5831
rect 11704 5797 11738 5831
rect 19349 5797 19383 5831
rect 7564 5729 7598 5763
rect 10333 5729 10367 5763
rect 10793 5729 10827 5763
rect 11437 5729 11471 5763
rect 13093 5729 13127 5763
rect 13360 5729 13394 5763
rect 15669 5729 15703 5763
rect 16681 5729 16715 5763
rect 20269 5729 20303 5763
rect 6929 5661 6963 5695
rect 7297 5661 7331 5695
rect 10885 5661 10919 5695
rect 10977 5661 11011 5695
rect 14749 5661 14783 5695
rect 15761 5661 15795 5695
rect 15945 5661 15979 5695
rect 16865 5661 16899 5695
rect 19533 5661 19567 5695
rect 18889 5593 18923 5627
rect 6285 5525 6319 5559
rect 8677 5525 8711 5559
rect 10149 5525 10183 5559
rect 12817 5525 12851 5559
rect 20453 5525 20487 5559
rect 8217 5321 8251 5355
rect 13001 5321 13035 5355
rect 14013 5321 14047 5355
rect 18061 5321 18095 5355
rect 19625 5321 19659 5355
rect 8493 5253 8527 5287
rect 9045 5185 9079 5219
rect 13645 5185 13679 5219
rect 14565 5185 14599 5219
rect 18613 5185 18647 5219
rect 20269 5185 20303 5219
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 10241 5117 10275 5151
rect 11897 5117 11931 5151
rect 13369 5117 13403 5151
rect 19073 5117 19107 5151
rect 20085 5117 20119 5151
rect 20637 5117 20671 5151
rect 8953 5049 8987 5083
rect 10508 5049 10542 5083
rect 14381 5049 14415 5083
rect 18429 5049 18463 5083
rect 18521 5049 18555 5083
rect 8861 4981 8895 5015
rect 11621 4981 11655 5015
rect 13461 4981 13495 5015
rect 14473 4981 14507 5015
rect 19257 4981 19291 5015
rect 19993 4981 20027 5015
rect 20821 4981 20855 5015
rect 7665 4777 7699 4811
rect 10609 4777 10643 4811
rect 14197 4777 14231 4811
rect 14289 4777 14323 4811
rect 6552 4709 6586 4743
rect 19432 4709 19466 4743
rect 6285 4641 6319 4675
rect 8953 4641 8987 4675
rect 9045 4641 9079 4675
rect 10977 4641 11011 4675
rect 17049 4641 17083 4675
rect 17316 4641 17350 4675
rect 19165 4641 19199 4675
rect 9137 4573 9171 4607
rect 11069 4573 11103 4607
rect 11253 4573 11287 4607
rect 14381 4573 14415 4607
rect 8585 4505 8619 4539
rect 13829 4437 13863 4471
rect 18429 4437 18463 4471
rect 20545 4437 20579 4471
rect 9229 4233 9263 4267
rect 16957 4233 16991 4267
rect 19441 4233 19475 4267
rect 19717 4233 19751 4267
rect 7849 4097 7883 4131
rect 10057 4097 10091 4131
rect 11069 4097 11103 4131
rect 13093 4097 13127 4131
rect 14657 4097 14691 4131
rect 15209 4097 15243 4131
rect 17509 4097 17543 4131
rect 18061 4097 18095 4131
rect 20269 4097 20303 4131
rect 9965 4029 9999 4063
rect 13001 4029 13035 4063
rect 15476 4029 15510 4063
rect 20729 4029 20763 4063
rect 8116 3961 8150 3995
rect 9873 3961 9907 3995
rect 18328 3961 18362 3995
rect 9505 3893 9539 3927
rect 10517 3893 10551 3927
rect 10885 3893 10919 3927
rect 10977 3893 11011 3927
rect 11805 3893 11839 3927
rect 12541 3893 12575 3927
rect 12909 3893 12943 3927
rect 14105 3893 14139 3927
rect 14473 3893 14507 3927
rect 14565 3893 14599 3927
rect 16589 3893 16623 3927
rect 17325 3893 17359 3927
rect 17417 3893 17451 3927
rect 20085 3893 20119 3927
rect 20177 3893 20211 3927
rect 20913 3893 20947 3927
rect 8493 3689 8527 3723
rect 9137 3689 9171 3723
rect 12725 3689 12759 3723
rect 14657 3689 14691 3723
rect 15117 3689 15151 3723
rect 17049 3689 17083 3723
rect 17509 3689 17543 3723
rect 17877 3689 17911 3723
rect 17969 3689 18003 3723
rect 19257 3689 19291 3723
rect 19441 3689 19475 3723
rect 9956 3621 9990 3655
rect 7113 3553 7147 3587
rect 7380 3553 7414 3587
rect 11612 3553 11646 3587
rect 13544 3553 13578 3587
rect 9689 3485 9723 3519
rect 11345 3485 11379 3519
rect 13277 3485 13311 3519
rect 15301 3553 15335 3587
rect 15568 3553 15602 3587
rect 18889 3553 18923 3587
rect 18153 3485 18187 3519
rect 19809 3553 19843 3587
rect 19901 3485 19935 3519
rect 20085 3485 20119 3519
rect 19257 3417 19291 3451
rect 11069 3349 11103 3383
rect 15117 3349 15151 3383
rect 16681 3349 16715 3383
rect 19073 3349 19107 3383
rect 8217 3145 8251 3179
rect 8493 3145 8527 3179
rect 10977 3145 11011 3179
rect 11345 3145 11379 3179
rect 14289 3145 14323 3179
rect 14381 3145 14415 3179
rect 14749 3145 14783 3179
rect 15117 3145 15151 3179
rect 16037 3145 16071 3179
rect 19441 3145 19475 3179
rect 6837 3009 6871 3043
rect 9045 3009 9079 3043
rect 11989 3009 12023 3043
rect 7104 2941 7138 2975
rect 8861 2941 8895 2975
rect 9597 2941 9631 2975
rect 9864 2941 9898 2975
rect 11713 2941 11747 2975
rect 12909 2941 12943 2975
rect 13176 2941 13210 2975
rect 15761 3009 15795 3043
rect 18245 3077 18279 3111
rect 20729 3077 20763 3111
rect 16681 3009 16715 3043
rect 19993 3009 20027 3043
rect 14565 2941 14599 2975
rect 16037 2941 16071 2975
rect 17417 2941 17451 2975
rect 18061 2941 18095 2975
rect 18705 2941 18739 2975
rect 20545 2941 20579 2975
rect 8953 2873 8987 2907
rect 11805 2873 11839 2907
rect 14381 2873 14415 2907
rect 18981 2873 19015 2907
rect 12449 2805 12483 2839
rect 15485 2805 15519 2839
rect 15577 2805 15611 2839
rect 16129 2805 16163 2839
rect 16497 2805 16531 2839
rect 16589 2805 16623 2839
rect 17601 2805 17635 2839
rect 19809 2805 19843 2839
rect 19901 2805 19935 2839
rect 7389 2601 7423 2635
rect 8401 2601 8435 2635
rect 10149 2601 10183 2635
rect 13369 2601 13403 2635
rect 15853 2601 15887 2635
rect 16221 2601 16255 2635
rect 17877 2601 17911 2635
rect 20729 2601 20763 2635
rect 10517 2533 10551 2567
rect 10609 2533 10643 2567
rect 7757 2465 7791 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 16313 2465 16347 2499
rect 16957 2465 16991 2499
rect 17693 2465 17727 2499
rect 18429 2465 18463 2499
rect 19441 2465 19475 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 7849 2397 7883 2431
rect 8033 2397 8067 2431
rect 10793 2397 10827 2431
rect 13461 2397 13495 2431
rect 13645 2397 13679 2431
rect 16405 2397 16439 2431
rect 13001 2329 13035 2363
rect 19625 2329 19659 2363
rect 11621 2261 11655 2295
rect 12173 2261 12207 2295
rect 17141 2261 17175 2295
rect 18613 2261 18647 2295
rect 20177 2261 20211 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 19886 19864 19892 19916
rect 19944 19904 19950 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 19944 19876 20545 19904
rect 19944 19864 19950 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 20162 19496 20168 19508
rect 20123 19468 20168 19496
rect 20162 19456 20168 19468
rect 20220 19456 20226 19508
rect 15930 19252 15936 19304
rect 15988 19292 15994 19304
rect 16485 19295 16543 19301
rect 16485 19292 16497 19295
rect 15988 19264 16497 19292
rect 15988 19252 15994 19264
rect 16485 19261 16497 19264
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18325 19295 18383 19301
rect 18325 19292 18337 19295
rect 17920 19264 18337 19292
rect 17920 19252 17926 19264
rect 18325 19261 18337 19264
rect 18371 19261 18383 19295
rect 18325 19255 18383 19261
rect 18874 19252 18880 19304
rect 18932 19292 18938 19304
rect 19058 19292 19064 19304
rect 18932 19264 19064 19292
rect 18932 19252 18938 19264
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 19978 19292 19984 19304
rect 19939 19264 19984 19292
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 5718 19184 5724 19236
rect 5776 19224 5782 19236
rect 20548 19224 20576 19255
rect 5776 19196 20576 19224
rect 5776 19184 5782 19196
rect 16669 19159 16727 19165
rect 16669 19125 16681 19159
rect 16715 19156 16727 19159
rect 17770 19156 17776 19168
rect 16715 19128 17776 19156
rect 16715 19125 16727 19128
rect 16669 19119 16727 19125
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18506 19156 18512 19168
rect 18467 19128 18512 19156
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 20717 19159 20775 19165
rect 20717 19125 20729 19159
rect 20763 19156 20775 19159
rect 20806 19156 20812 19168
rect 20763 19128 20812 19156
rect 20763 19125 20775 19128
rect 20717 19119 20775 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 9953 18887 10011 18893
rect 9953 18853 9965 18887
rect 9999 18884 10011 18887
rect 15746 18884 15752 18896
rect 9999 18856 15752 18884
rect 9999 18853 10011 18856
rect 9953 18847 10011 18853
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 15930 18884 15936 18896
rect 15891 18856 15936 18884
rect 15930 18844 15936 18856
rect 15988 18844 15994 18896
rect 17862 18884 17868 18896
rect 17823 18856 17868 18884
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 19886 18884 19892 18896
rect 19847 18856 19892 18884
rect 19886 18844 19892 18856
rect 19944 18844 19950 18896
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 12069 18819 12127 18825
rect 12069 18816 12081 18819
rect 11756 18788 12081 18816
rect 11756 18776 11762 18788
rect 12069 18785 12081 18788
rect 12115 18785 12127 18819
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 12069 18779 12127 18785
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 17586 18816 17592 18828
rect 17547 18788 17592 18816
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 19610 18816 19616 18828
rect 19571 18788 19616 18816
rect 19610 18776 19616 18788
rect 19668 18776 19674 18828
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 12360 18680 12388 18711
rect 19978 18680 19984 18692
rect 12360 18652 19984 18680
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 20162 18408 20168 18420
rect 20123 18380 20168 18408
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 15746 18232 15752 18284
rect 15804 18272 15810 18284
rect 15804 18244 20576 18272
rect 15804 18232 15810 18244
rect 7650 18164 7656 18216
rect 7708 18204 7714 18216
rect 20548 18213 20576 18244
rect 7745 18207 7803 18213
rect 7745 18204 7757 18207
rect 7708 18176 7757 18204
rect 7708 18164 7714 18176
rect 7745 18173 7757 18176
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 19987 18207 20045 18213
rect 19987 18173 19999 18207
rect 20033 18173 20045 18207
rect 19987 18167 20045 18173
rect 20533 18207 20591 18213
rect 20533 18173 20545 18207
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 8021 18139 8079 18145
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 19996 18136 20024 18167
rect 8067 18108 20024 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 15473 17867 15531 17873
rect 15473 17833 15485 17867
rect 15519 17864 15531 17867
rect 17862 17864 17868 17876
rect 15519 17836 17868 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 20438 17864 20444 17876
rect 20399 17836 20444 17864
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 11425 17731 11483 17737
rect 11425 17697 11437 17731
rect 11471 17728 11483 17731
rect 11882 17728 11888 17740
rect 11471 17700 11888 17728
rect 11471 17697 11483 17700
rect 11425 17691 11483 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 14458 17688 14464 17740
rect 14516 17728 14522 17740
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 14516 17700 15301 17728
rect 14516 17688 14522 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17697 20315 17731
rect 20257 17691 20315 17697
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 20272 17660 20300 17691
rect 11747 17632 20300 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 14458 17184 14464 17196
rect 14419 17156 14464 17184
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 14182 17116 14188 17128
rect 14143 17088 14188 17116
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 19944 17088 19993 17116
rect 19944 17076 19950 17088
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 17310 17008 17316 17060
rect 17368 17048 17374 17060
rect 20548 17048 20576 17079
rect 17368 17020 20576 17048
rect 17368 17008 17374 17020
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 17310 16708 17316 16720
rect 17271 16680 17316 16708
rect 17310 16668 17316 16680
rect 17368 16668 17374 16720
rect 19886 16708 19892 16720
rect 19847 16680 19892 16708
rect 19886 16668 19892 16680
rect 19944 16668 19950 16720
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 17037 16643 17095 16649
rect 17037 16640 17049 16643
rect 16448 16612 17049 16640
rect 16448 16600 16454 16612
rect 17037 16609 17049 16612
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 19613 16643 19671 16649
rect 19613 16640 19625 16643
rect 19576 16612 19625 16640
rect 19576 16600 19582 16612
rect 19613 16609 19625 16612
rect 19659 16609 19671 16643
rect 19613 16603 19671 16609
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 19978 16028 19984 16040
rect 19939 16000 19984 16028
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20530 16028 20536 16040
rect 20491 16000 20536 16028
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 14185 15623 14243 15629
rect 14185 15589 14197 15623
rect 14231 15620 14243 15623
rect 20530 15620 20536 15632
rect 14231 15592 20536 15620
rect 14231 15589 14243 15592
rect 14185 15583 14243 15589
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 11790 15552 11796 15564
rect 11751 15524 11796 15552
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 13906 15552 13912 15564
rect 13867 15524 13912 15552
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 20254 15552 20260 15564
rect 20215 15524 20260 15552
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 12084 15416 12112 15447
rect 19978 15416 19984 15428
rect 12084 15388 19984 15416
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 20714 15144 20720 15156
rect 20675 15116 20720 15144
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 9582 14940 9588 14952
rect 9543 14912 9588 14940
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 16482 14900 16488 14952
rect 16540 14940 16546 14952
rect 20533 14943 20591 14949
rect 20533 14940 20545 14943
rect 16540 14912 20545 14940
rect 16540 14900 16546 14912
rect 20533 14909 20545 14912
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 9861 14875 9919 14881
rect 9861 14841 9873 14875
rect 9907 14872 9919 14875
rect 20254 14872 20260 14884
rect 9907 14844 20260 14872
rect 9907 14841 9919 14844
rect 9861 14835 9919 14841
rect 20254 14832 20260 14844
rect 20312 14832 20318 14884
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 19886 14600 19892 14612
rect 19847 14572 19892 14600
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 20438 14600 20444 14612
rect 20399 14572 20444 14600
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 8386 14464 8392 14476
rect 8347 14436 8392 14464
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 19702 14464 19708 14476
rect 19663 14436 19708 14464
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 20257 14467 20315 14473
rect 20257 14433 20269 14467
rect 20303 14433 20315 14467
rect 20257 14427 20315 14433
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 16482 14396 16488 14408
rect 8711 14368 16488 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 20272 14328 20300 14427
rect 11112 14300 20300 14328
rect 11112 14288 11118 14300
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 16356 14028 17509 14056
rect 16356 14016 16362 14028
rect 17497 14025 17509 14028
rect 17543 14025 17555 14059
rect 17497 14019 17555 14025
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19429 14059 19487 14065
rect 19429 14056 19441 14059
rect 19300 14028 19441 14056
rect 19300 14016 19306 14028
rect 19429 14025 19441 14028
rect 19475 14025 19487 14059
rect 19429 14019 19487 14025
rect 11054 13920 11060 13932
rect 11015 13892 11060 13920
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 19886 13880 19892 13932
rect 19944 13920 19950 13932
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 19944 13892 20177 13920
rect 19944 13880 19950 13892
rect 20165 13889 20177 13892
rect 20211 13889 20223 13923
rect 20165 13883 20223 13889
rect 10502 13812 10508 13864
rect 10560 13852 10566 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10560 13824 10793 13852
rect 10560 13812 10566 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 16114 13852 16120 13864
rect 16075 13824 16120 13852
rect 10781 13815 10839 13821
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 16384 13855 16442 13861
rect 16384 13821 16396 13855
rect 16430 13852 16442 13855
rect 17126 13852 17132 13864
rect 16430 13824 17132 13852
rect 16430 13821 16442 13824
rect 16384 13815 16442 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19426 13852 19432 13864
rect 19291 13824 19432 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19981 13855 20039 13861
rect 19981 13821 19993 13855
rect 20027 13852 20039 13855
rect 20070 13852 20076 13864
rect 20027 13824 20076 13852
rect 20027 13821 20039 13824
rect 19981 13815 20039 13821
rect 20070 13812 20076 13824
rect 20128 13812 20134 13864
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 19242 13512 19248 13524
rect 19203 13484 19248 13512
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19702 13404 19708 13456
rect 19760 13444 19766 13456
rect 19889 13447 19947 13453
rect 19889 13444 19901 13447
rect 19760 13416 19901 13444
rect 19760 13404 19766 13416
rect 19889 13413 19901 13416
rect 19935 13413 19947 13447
rect 19889 13407 19947 13413
rect 19061 13379 19119 13385
rect 19061 13345 19073 13379
rect 19107 13376 19119 13379
rect 19334 13376 19340 13388
rect 19107 13348 19340 13376
rect 19107 13345 19119 13348
rect 19061 13339 19119 13345
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13345 19671 13379
rect 19613 13339 19671 13345
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 19628 13308 19656 13339
rect 12584 13280 19656 13308
rect 12584 13268 12590 13280
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 15105 12971 15163 12977
rect 15105 12937 15117 12971
rect 15151 12968 15163 12971
rect 15654 12968 15660 12980
rect 15151 12940 15660 12968
rect 15151 12937 15163 12940
rect 15105 12931 15163 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 16945 12971 17003 12977
rect 16945 12937 16957 12971
rect 16991 12968 17003 12971
rect 17586 12968 17592 12980
rect 16991 12940 17592 12968
rect 16991 12937 17003 12940
rect 16945 12931 17003 12937
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 19242 12968 19248 12980
rect 19203 12940 19248 12968
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 15654 12832 15660 12844
rect 15615 12804 15660 12832
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 17586 12832 17592 12844
rect 17547 12804 17592 12832
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 19484 12804 19901 12832
rect 19484 12792 19490 12804
rect 19889 12801 19901 12804
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14148 12736 17540 12764
rect 14148 12724 14154 12736
rect 16482 12656 16488 12708
rect 16540 12696 16546 12708
rect 17405 12699 17463 12705
rect 17405 12696 17417 12699
rect 16540 12668 17417 12696
rect 16540 12656 16546 12668
rect 17405 12665 17417 12668
rect 17451 12665 17463 12699
rect 17512 12696 17540 12736
rect 17678 12724 17684 12776
rect 17736 12764 17742 12776
rect 19061 12767 19119 12773
rect 19061 12764 19073 12767
rect 17736 12736 19073 12764
rect 17736 12724 17742 12736
rect 19061 12733 19073 12736
rect 19107 12733 19119 12767
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19061 12727 19119 12733
rect 19168 12736 19625 12764
rect 19168 12696 19196 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 19794 12724 19800 12776
rect 19852 12764 19858 12776
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 19852 12736 20361 12764
rect 19852 12724 19858 12736
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 17512 12668 19196 12696
rect 17405 12659 17463 12665
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 19886 12696 19892 12708
rect 19484 12668 19892 12696
rect 19484 12656 19490 12668
rect 19886 12656 19892 12668
rect 19944 12656 19950 12708
rect 20254 12656 20260 12708
rect 20312 12696 20318 12708
rect 20625 12699 20683 12705
rect 20625 12696 20637 12699
rect 20312 12668 20637 12696
rect 20312 12656 20318 12668
rect 20625 12665 20637 12668
rect 20671 12665 20683 12699
rect 20625 12659 20683 12665
rect 15470 12628 15476 12640
rect 15431 12600 15476 12628
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 17310 12628 17316 12640
rect 15620 12600 15665 12628
rect 17271 12600 17316 12628
rect 15620 12588 15626 12600
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 15381 12427 15439 12433
rect 15381 12393 15393 12427
rect 15427 12424 15439 12427
rect 15470 12424 15476 12436
rect 15427 12396 15476 12424
rect 15427 12393 15439 12396
rect 15381 12387 15439 12393
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 17313 12427 17371 12433
rect 17313 12393 17325 12427
rect 17359 12393 17371 12427
rect 20438 12424 20444 12436
rect 20399 12396 20444 12424
rect 17313 12387 17371 12393
rect 13446 12316 13452 12368
rect 13504 12365 13510 12368
rect 13504 12359 13568 12365
rect 13504 12325 13522 12359
rect 13556 12325 13568 12359
rect 16114 12356 16120 12368
rect 13504 12319 13568 12325
rect 15948 12328 16120 12356
rect 13504 12316 13510 12319
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 15378 12288 15384 12300
rect 13311 12260 15384 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 15378 12248 15384 12260
rect 15436 12288 15442 12300
rect 15948 12297 15976 12328
rect 16114 12316 16120 12328
rect 16172 12356 16178 12368
rect 17328 12356 17356 12387
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 17586 12356 17592 12368
rect 16172 12328 16896 12356
rect 17328 12328 17592 12356
rect 16172 12316 16178 12328
rect 15933 12291 15991 12297
rect 15933 12288 15945 12291
rect 15436 12260 15945 12288
rect 15436 12248 15442 12260
rect 15933 12257 15945 12260
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 16200 12291 16258 12297
rect 16200 12257 16212 12291
rect 16246 12288 16258 12291
rect 16758 12288 16764 12300
rect 16246 12260 16764 12288
rect 16246 12257 16258 12260
rect 16200 12251 16258 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16868 12288 16896 12328
rect 17586 12316 17592 12328
rect 17644 12356 17650 12368
rect 17834 12359 17892 12365
rect 17834 12356 17846 12359
rect 17644 12328 17846 12356
rect 17644 12316 17650 12328
rect 17834 12325 17846 12328
rect 17880 12325 17892 12359
rect 17834 12319 17892 12325
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19705 12359 19763 12365
rect 19705 12356 19717 12359
rect 19392 12328 19717 12356
rect 19392 12316 19398 12328
rect 19705 12325 19717 12328
rect 19751 12325 19763 12359
rect 19705 12319 19763 12325
rect 16868 12260 17632 12288
rect 17604 12232 17632 12260
rect 19150 12248 19156 12300
rect 19208 12288 19214 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19208 12260 19441 12288
rect 19208 12248 19214 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 20254 12288 20260 12300
rect 20215 12260 20260 12288
rect 19429 12251 19487 12257
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 17586 12220 17592 12232
rect 17547 12192 17592 12220
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 15838 12084 15844 12096
rect 14691 12056 15844 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 18969 12087 19027 12093
rect 18969 12084 18981 12087
rect 18932 12056 18981 12084
rect 18932 12044 18938 12056
rect 18969 12053 18981 12056
rect 19015 12053 19027 12087
rect 18969 12047 19027 12053
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 15105 11883 15163 11889
rect 15105 11849 15117 11883
rect 15151 11880 15163 11883
rect 15654 11880 15660 11892
rect 15151 11852 15660 11880
rect 15151 11849 15163 11852
rect 15105 11843 15163 11849
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16758 11880 16764 11892
rect 16719 11852 16764 11880
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13446 11744 13452 11756
rect 13403 11716 13452 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 15378 11744 15384 11756
rect 15339 11716 15384 11744
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 17310 11704 17316 11756
rect 17368 11744 17374 11756
rect 17497 11747 17555 11753
rect 17497 11744 17509 11747
rect 17368 11716 17509 11744
rect 17368 11704 17374 11716
rect 17497 11713 17509 11716
rect 17543 11713 17555 11747
rect 18506 11744 18512 11756
rect 17497 11707 17555 11713
rect 18064 11716 18512 11744
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 13630 11676 13636 11688
rect 13127 11648 13636 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 15396 11676 15424 11704
rect 15654 11685 15660 11688
rect 15648 11676 15660 11685
rect 13771 11648 15424 11676
rect 15615 11648 15660 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 15648 11639 15660 11648
rect 15654 11636 15660 11639
rect 15712 11636 15718 11688
rect 18064 11685 18092 11716
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 20622 11704 20628 11756
rect 20680 11744 20686 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20680 11716 20729 11744
rect 20680 11704 20686 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18874 11685 18880 11688
rect 18608 11679 18666 11685
rect 18608 11676 18620 11679
rect 18472 11648 18620 11676
rect 18472 11636 18478 11648
rect 18608 11645 18620 11648
rect 18654 11645 18666 11679
rect 18868 11676 18880 11685
rect 18787 11648 18880 11676
rect 18608 11639 18666 11645
rect 18868 11639 18880 11648
rect 18932 11676 18938 11688
rect 20824 11676 20852 11707
rect 18932 11648 20852 11676
rect 18874 11636 18880 11639
rect 18932 11636 18938 11648
rect 13992 11611 14050 11617
rect 12728 11580 13952 11608
rect 12728 11549 12756 11580
rect 12713 11543 12771 11549
rect 12713 11509 12725 11543
rect 12759 11509 12771 11543
rect 12713 11503 12771 11509
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 13924 11540 13952 11580
rect 13992 11577 14004 11611
rect 14038 11608 14050 11611
rect 15838 11608 15844 11620
rect 14038 11580 15844 11608
rect 14038 11577 14050 11580
rect 13992 11571 14050 11577
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 19610 11608 19616 11620
rect 16132 11580 19616 11608
rect 16132 11540 16160 11580
rect 19610 11568 19616 11580
rect 19668 11568 19674 11620
rect 21910 11608 21916 11620
rect 19812 11580 21916 11608
rect 13228 11512 13273 11540
rect 13924 11512 16160 11540
rect 18233 11543 18291 11549
rect 13228 11500 13234 11512
rect 18233 11509 18245 11543
rect 18279 11540 18291 11543
rect 19812 11540 19840 11580
rect 21910 11568 21916 11580
rect 21968 11568 21974 11620
rect 19978 11540 19984 11552
rect 18279 11512 19840 11540
rect 19939 11512 19984 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20254 11540 20260 11552
rect 20215 11512 20260 11540
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 20625 11543 20683 11549
rect 20625 11540 20637 11543
rect 20496 11512 20637 11540
rect 20496 11500 20502 11512
rect 20625 11509 20637 11512
rect 20671 11509 20683 11543
rect 20625 11503 20683 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 658 11296 664 11348
rect 716 11336 722 11348
rect 716 11308 13584 11336
rect 716 11296 722 11308
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 13556 11268 13584 11308
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13688 11308 14105 11336
rect 13688 11296 13694 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15562 11336 15568 11348
rect 15335 11308 15568 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 15930 11336 15936 11348
rect 15795 11308 15936 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 19334 11336 19340 11348
rect 18739 11308 19340 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 20533 11339 20591 11345
rect 20533 11305 20545 11339
rect 20579 11305 20591 11339
rect 20533 11299 20591 11305
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 4120 11240 13492 11268
rect 13556 11240 15669 11268
rect 4120 11228 4126 11240
rect 12704 11203 12762 11209
rect 12704 11169 12716 11203
rect 12750 11200 12762 11203
rect 13078 11200 13084 11212
rect 12750 11172 13084 11200
rect 12750 11169 12762 11172
rect 12704 11163 12762 11169
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 13464 11132 13492 11240
rect 15657 11237 15669 11240
rect 15703 11268 15715 11271
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 15703 11240 16129 11268
rect 15703 11237 15715 11240
rect 15657 11231 15715 11237
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 18874 11268 18880 11280
rect 16117 11231 16175 11237
rect 16776 11240 18880 11268
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 16485 11203 16543 11209
rect 16485 11200 16497 11203
rect 15620 11172 16497 11200
rect 15620 11160 15626 11172
rect 16485 11169 16497 11172
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 15838 11132 15844 11144
rect 12492 11104 12537 11132
rect 13464 11104 15700 11132
rect 15799 11104 15844 11132
rect 12492 11092 12498 11104
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13817 11067 13875 11073
rect 13817 11064 13829 11067
rect 13504 11036 13829 11064
rect 13504 11024 13510 11036
rect 13817 11033 13829 11036
rect 13863 11033 13875 11067
rect 15672 11064 15700 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 16776 11064 16804 11240
rect 18874 11228 18880 11240
rect 18932 11228 18938 11280
rect 19420 11271 19478 11277
rect 19420 11237 19432 11271
rect 19466 11268 19478 11271
rect 19978 11268 19984 11280
rect 19466 11240 19984 11268
rect 19466 11237 19478 11240
rect 19420 11231 19478 11237
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 17120 11203 17178 11209
rect 17120 11169 17132 11203
rect 17166 11200 17178 11203
rect 20548 11200 20576 11299
rect 20622 11200 20628 11212
rect 17166 11172 20628 11200
rect 17166 11169 17178 11172
rect 17120 11163 17178 11169
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 16853 11135 16911 11141
rect 16853 11101 16865 11135
rect 16899 11101 16911 11135
rect 18414 11132 18420 11144
rect 16853 11095 16911 11101
rect 17880 11104 18420 11132
rect 15672 11036 16804 11064
rect 13817 11027 13875 11033
rect 16301 10999 16359 11005
rect 16301 10965 16313 10999
rect 16347 10996 16359 10999
rect 16868 10996 16896 11095
rect 17586 10996 17592 11008
rect 16347 10968 17592 10996
rect 16347 10965 16359 10968
rect 16301 10959 16359 10965
rect 17586 10956 17592 10968
rect 17644 10996 17650 11008
rect 17880 10996 17908 11104
rect 18414 11092 18420 11104
rect 18472 11132 18478 11144
rect 19153 11135 19211 11141
rect 19153 11132 19165 11135
rect 18472 11104 19165 11132
rect 18472 11092 18478 11104
rect 19153 11101 19165 11104
rect 19199 11101 19211 11135
rect 19153 11095 19211 11101
rect 17644 10968 17908 10996
rect 17644 10956 17650 10968
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18233 10999 18291 11005
rect 18233 10996 18245 10999
rect 18012 10968 18245 10996
rect 18012 10956 18018 10968
rect 18233 10965 18245 10968
rect 18279 10965 18291 10999
rect 18233 10959 18291 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 19518 10792 19524 10804
rect 15427 10764 19524 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 19061 10727 19119 10733
rect 19061 10724 19073 10727
rect 12452 10696 19073 10724
rect 12452 10597 12480 10696
rect 19061 10693 19073 10696
rect 19107 10693 19119 10727
rect 19061 10687 19119 10693
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16482 10656 16488 10668
rect 16071 10628 16488 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16816 10628 17049 10656
rect 16816 10616 16822 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18012 10628 18613 10656
rect 18012 10616 18018 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 19978 10656 19984 10668
rect 19751 10628 19984 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20530 10656 20536 10668
rect 20491 10628 20536 10656
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 20622 10616 20628 10668
rect 20680 10656 20686 10668
rect 20680 10628 20725 10656
rect 20680 10616 20686 10628
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 16574 10588 16580 10600
rect 12437 10551 12495 10557
rect 16500 10560 16580 10588
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12713 10523 12771 10529
rect 12713 10520 12725 10523
rect 12032 10492 12725 10520
rect 12032 10480 12038 10492
rect 12713 10489 12725 10492
rect 12759 10489 12771 10523
rect 12713 10483 12771 10489
rect 15286 10480 15292 10532
rect 15344 10520 15350 10532
rect 15841 10523 15899 10529
rect 15841 10520 15853 10523
rect 15344 10492 15853 10520
rect 15344 10480 15350 10492
rect 15841 10489 15853 10492
rect 15887 10489 15899 10523
rect 15841 10483 15899 10489
rect 15746 10452 15752 10464
rect 15707 10424 15752 10452
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 16500 10461 16528 10560
rect 16574 10548 16580 10560
rect 16632 10548 16638 10600
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 18104 10560 18429 10588
rect 18104 10548 18110 10560
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19392 10560 19441 10588
rect 19392 10548 19398 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20254 10588 20260 10600
rect 19567 10560 20260 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 18509 10523 18567 10529
rect 18509 10489 18521 10523
rect 18555 10520 18567 10523
rect 18555 10492 20116 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 16485 10455 16543 10461
rect 16485 10421 16497 10455
rect 16531 10421 16543 10455
rect 16485 10415 16543 10421
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16632 10424 16865 10452
rect 16632 10412 16638 10424
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 16853 10415 16911 10421
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 18049 10455 18107 10461
rect 17000 10424 17045 10452
rect 17000 10412 17006 10424
rect 18049 10421 18061 10455
rect 18095 10452 18107 10455
rect 18598 10452 18604 10464
rect 18095 10424 18604 10452
rect 18095 10421 18107 10424
rect 18049 10415 18107 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 20088 10461 20116 10492
rect 20073 10455 20131 10461
rect 20073 10421 20085 10455
rect 20119 10421 20131 10455
rect 20438 10452 20444 10464
rect 20399 10424 20444 10452
rect 20073 10415 20131 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13906 10248 13912 10260
rect 13311 10220 13912 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 16945 10251 17003 10257
rect 16945 10248 16957 10251
rect 15804 10220 16957 10248
rect 15804 10208 15810 10220
rect 16945 10217 16957 10220
rect 16991 10217 17003 10251
rect 16945 10211 17003 10217
rect 17856 10183 17914 10189
rect 17856 10149 17868 10183
rect 17902 10180 17914 10183
rect 17954 10180 17960 10192
rect 17902 10152 17960 10180
rect 17902 10149 17914 10152
rect 17856 10143 17914 10149
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 20438 10180 20444 10192
rect 19628 10152 20444 10180
rect 19628 10124 19656 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13044 10084 13645 10112
rect 13044 10072 13050 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10112 15347 10115
rect 15378 10112 15384 10124
rect 15335 10084 15384 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15556 10115 15614 10121
rect 15556 10081 15568 10115
rect 15602 10112 15614 10115
rect 15838 10112 15844 10124
rect 15602 10084 15844 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 19610 10112 19616 10124
rect 19571 10084 19616 10112
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 20257 10115 20315 10121
rect 19760 10084 19805 10112
rect 19760 10072 19766 10084
rect 20257 10081 20269 10115
rect 20303 10112 20315 10115
rect 20346 10112 20352 10124
rect 20303 10084 20352 10112
rect 20303 10081 20315 10084
rect 20257 10075 20315 10081
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 12860 10016 13737 10044
rect 12860 10004 12866 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10013 13875 10047
rect 17586 10044 17592 10056
rect 17547 10016 17592 10044
rect 13817 10007 13875 10013
rect 13832 9976 13860 10007
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 18984 10016 19809 10044
rect 18984 9988 19012 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 18966 9976 18972 9988
rect 13740 9948 13860 9976
rect 18879 9948 18972 9976
rect 13740 9920 13768 9948
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 13722 9868 13728 9920
rect 13780 9868 13786 9920
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 16540 9880 16681 9908
rect 16540 9868 16546 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 19058 9868 19064 9920
rect 19116 9908 19122 9920
rect 19245 9911 19303 9917
rect 19245 9908 19257 9911
rect 19116 9880 19257 9908
rect 19116 9868 19122 9880
rect 19245 9877 19257 9880
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 20441 9911 20499 9917
rect 20441 9908 20453 9911
rect 19392 9880 20453 9908
rect 19392 9868 19398 9880
rect 20441 9877 20453 9880
rect 20487 9877 20499 9911
rect 20441 9871 20499 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 15378 9704 15384 9716
rect 11940 9676 12204 9704
rect 15291 9676 15384 9704
rect 11940 9664 11946 9676
rect 11057 9639 11115 9645
rect 11057 9605 11069 9639
rect 11103 9636 11115 9639
rect 11790 9636 11796 9648
rect 11103 9608 11796 9636
rect 11103 9605 11115 9608
rect 11057 9599 11115 9605
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 11606 9568 11612 9580
rect 11567 9540 11612 9568
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10928 9472 10977 9500
rect 10928 9460 10934 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 12176 9500 12204 9676
rect 15378 9664 15384 9676
rect 15436 9704 15442 9716
rect 17586 9704 17592 9716
rect 15436 9676 17592 9704
rect 15436 9664 15442 9676
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13722 9509 13728 9512
rect 10965 9463 11023 9469
rect 11063 9472 12204 9500
rect 13449 9503 13507 9509
rect 10410 9392 10416 9444
rect 10468 9432 10474 9444
rect 11063 9432 11091 9472
rect 13449 9469 13461 9503
rect 13495 9469 13507 9503
rect 13716 9500 13728 9509
rect 13683 9472 13728 9500
rect 13449 9463 13507 9469
rect 13716 9463 13728 9472
rect 10468 9404 11091 9432
rect 11425 9435 11483 9441
rect 10468 9392 10474 9404
rect 11425 9401 11437 9435
rect 11471 9432 11483 9435
rect 11882 9432 11888 9444
rect 11471 9404 11888 9432
rect 11471 9401 11483 9404
rect 11425 9395 11483 9401
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 13464 9432 13492 9463
rect 13722 9460 13728 9463
rect 13780 9460 13786 9512
rect 15396 9509 15424 9664
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 17954 9568 17960 9580
rect 17543 9540 17960 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 13832 9472 15393 9500
rect 13832 9432 13860 9472
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 15648 9503 15706 9509
rect 15648 9469 15660 9503
rect 15694 9500 15706 9503
rect 16482 9500 16488 9512
rect 15694 9472 16488 9500
rect 15694 9469 15706 9472
rect 15648 9463 15706 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 17586 9460 17592 9512
rect 17644 9500 17650 9512
rect 18414 9500 18420 9512
rect 17644 9472 18420 9500
rect 17644 9460 17650 9472
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 18684 9503 18742 9509
rect 18684 9469 18696 9503
rect 18730 9500 18742 9503
rect 18966 9500 18972 9512
rect 18730 9472 18972 9500
rect 18730 9469 18742 9472
rect 18684 9463 18742 9469
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 20533 9503 20591 9509
rect 20533 9500 20545 9503
rect 19300 9472 20545 9500
rect 19300 9460 19306 9472
rect 20533 9469 20545 9472
rect 20579 9469 20591 9503
rect 20533 9463 20591 9469
rect 13464 9404 13860 9432
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 15068 9404 20760 9432
rect 15068 9392 15074 9404
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 10376 9336 10793 9364
rect 10376 9324 10382 9336
rect 10781 9333 10793 9336
rect 10827 9333 10839 9367
rect 10781 9327 10839 9333
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11112 9336 11529 9364
rect 11112 9324 11118 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11517 9327 11575 9333
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 15838 9364 15844 9376
rect 14875 9336 15844 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 16758 9364 16764 9376
rect 16719 9336 16764 9364
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 19794 9364 19800 9376
rect 19755 9336 19800 9364
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 20732 9373 20760 9404
rect 20717 9367 20775 9373
rect 20717 9333 20729 9367
rect 20763 9333 20775 9367
rect 20717 9327 20775 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9640 9132 9689 9160
rect 9640 9120 9646 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 9784 9132 11836 9160
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 9784 9092 9812 9132
rect 11808 9092 11836 9132
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 13817 9163 13875 9169
rect 13817 9160 13829 9163
rect 13780 9132 13829 9160
rect 13780 9120 13786 9132
rect 13817 9129 13829 9132
rect 13863 9129 13875 9163
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 13817 9123 13875 9129
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15749 9163 15807 9169
rect 15749 9129 15761 9163
rect 15795 9160 15807 9163
rect 15930 9160 15936 9172
rect 15795 9132 15936 9160
rect 15795 9129 15807 9132
rect 15749 9123 15807 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16390 9160 16396 9172
rect 16351 9132 16396 9160
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 15657 9095 15715 9101
rect 15657 9092 15669 9095
rect 5132 9064 9812 9092
rect 10796 9064 11744 9092
rect 11808 9064 15669 9092
rect 5132 9052 5138 9064
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9171 8996 10057 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9548 8928 10149 8956
rect 9548 8916 9554 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10244 8888 10272 8919
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 10796 8965 10824 9064
rect 11048 9027 11106 9033
rect 11048 8993 11060 9027
rect 11094 9024 11106 9027
rect 11606 9024 11612 9036
rect 11094 8996 11612 9024
rect 11094 8993 11106 8996
rect 11048 8987 11106 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11716 9024 11744 9064
rect 15657 9061 15669 9064
rect 15703 9061 15715 9095
rect 18598 9092 18604 9104
rect 15657 9055 15715 9061
rect 16684 9064 18604 9092
rect 12434 9024 12440 9036
rect 11716 8996 12440 9024
rect 12434 8984 12440 8996
rect 12492 9024 12498 9036
rect 12710 9033 12716 9036
rect 12704 9024 12716 9033
rect 12492 8996 12537 9024
rect 12671 8996 12716 9024
rect 12492 8984 12498 8996
rect 12704 8987 12716 8996
rect 12710 8984 12716 8987
rect 12768 8984 12774 9036
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 9024 13967 9027
rect 16684 9024 16712 9064
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 19242 9052 19248 9104
rect 19300 9101 19306 9104
rect 19300 9095 19364 9101
rect 19300 9061 19318 9095
rect 19352 9092 19364 9095
rect 19794 9092 19800 9104
rect 19352 9064 19800 9092
rect 19352 9061 19364 9064
rect 19300 9055 19364 9061
rect 19300 9052 19306 9055
rect 19794 9052 19800 9064
rect 19852 9052 19858 9104
rect 13955 8996 16712 9024
rect 16761 9027 16819 9033
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 17494 9024 17500 9036
rect 16807 8996 17500 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 18414 8984 18420 9036
rect 18472 9024 18478 9036
rect 19061 9027 19119 9033
rect 19061 9024 19073 9027
rect 18472 8996 19073 9024
rect 18472 8984 18478 8996
rect 19061 8993 19073 8996
rect 19107 8993 19119 9027
rect 19061 8987 19119 8993
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10376 8928 10793 8956
rect 10376 8916 10382 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 14056 8928 14105 8956
rect 14056 8916 14062 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 15838 8956 15844 8968
rect 15799 8928 15844 8956
rect 14093 8919 14151 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16850 8956 16856 8968
rect 16811 8928 16856 8956
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8956 17095 8959
rect 17126 8956 17132 8968
rect 17083 8928 17132 8956
rect 17083 8925 17095 8928
rect 17037 8919 17095 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 18601 8959 18659 8965
rect 18601 8925 18613 8959
rect 18647 8956 18659 8959
rect 18966 8956 18972 8968
rect 18647 8928 18972 8956
rect 18647 8925 18659 8928
rect 18601 8919 18659 8925
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 9364 8860 10272 8888
rect 9364 8848 9370 8860
rect 12161 8823 12219 8829
rect 12161 8789 12173 8823
rect 12207 8820 12219 8823
rect 12710 8820 12716 8832
rect 12207 8792 12716 8820
rect 12207 8789 12219 8792
rect 12161 8783 12219 8789
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 19426 8820 19432 8832
rect 13412 8792 19432 8820
rect 13412 8780 13418 8792
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 20438 8820 20444 8832
rect 20399 8792 20444 8820
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 11606 8616 11612 8628
rect 11567 8588 11612 8616
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 18601 8619 18659 8625
rect 18601 8616 18613 8619
rect 14854 8588 18613 8616
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 8570 8412 8576 8424
rect 8483 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8412 8634 8424
rect 10229 8415 10287 8421
rect 10229 8412 10241 8415
rect 8628 8384 10241 8412
rect 8628 8372 8634 8384
rect 10229 8381 10241 8384
rect 10275 8412 10287 8415
rect 10318 8412 10324 8424
rect 10275 8384 10324 8412
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 12989 8415 13047 8421
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13354 8412 13360 8424
rect 13035 8384 13360 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 14854 8421 14882 8588
rect 18601 8585 18613 8588
rect 18647 8585 18659 8619
rect 18601 8579 18659 8585
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 21085 8619 21143 8625
rect 21085 8616 21097 8619
rect 18932 8588 21097 8616
rect 18932 8576 18938 8588
rect 21085 8585 21097 8588
rect 21131 8585 21143 8619
rect 21085 8579 21143 8585
rect 15562 8548 15568 8560
rect 15523 8520 15568 8548
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 17494 8480 17500 8492
rect 17455 8452 17500 8480
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 19058 8480 19064 8492
rect 19019 8452 19064 8480
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19242 8480 19248 8492
rect 19203 8452 19248 8480
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8381 15807 8415
rect 15749 8375 15807 8381
rect 15841 8415 15899 8421
rect 15841 8381 15853 8415
rect 15887 8412 15899 8415
rect 15930 8412 15936 8424
rect 15887 8384 15936 8412
rect 15887 8381 15899 8384
rect 15841 8375 15899 8381
rect 8840 8347 8898 8353
rect 8840 8313 8852 8347
rect 8886 8344 8898 8347
rect 9306 8344 9312 8356
rect 8886 8316 9312 8344
rect 8886 8313 8898 8316
rect 8840 8307 8898 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 10474 8347 10532 8353
rect 10474 8344 10486 8347
rect 9968 8316 10486 8344
rect 9968 8285 9996 8316
rect 10474 8313 10486 8316
rect 10520 8344 10532 8347
rect 10962 8344 10968 8356
rect 10520 8316 10968 8344
rect 10520 8313 10532 8316
rect 10474 8307 10532 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 14550 8304 14556 8356
rect 14608 8344 14614 8356
rect 15105 8347 15163 8353
rect 15105 8344 15117 8347
rect 14608 8316 15117 8344
rect 14608 8304 14614 8316
rect 15105 8313 15117 8316
rect 15151 8313 15163 8347
rect 15105 8307 15163 8313
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8245 10011 8279
rect 9953 8239 10011 8245
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14277 8279 14335 8285
rect 14277 8276 14289 8279
rect 13964 8248 14289 8276
rect 13964 8236 13970 8248
rect 14277 8245 14289 8248
rect 14323 8276 14335 8279
rect 15764 8276 15792 8375
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 18966 8412 18972 8424
rect 18927 8384 18972 8412
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8381 19763 8415
rect 19705 8375 19763 8381
rect 19972 8415 20030 8421
rect 19972 8381 19984 8415
rect 20018 8412 20030 8415
rect 20438 8412 20444 8424
rect 20018 8384 20444 8412
rect 20018 8381 20030 8384
rect 19972 8375 20030 8381
rect 16108 8347 16166 8353
rect 16108 8313 16120 8347
rect 16154 8344 16166 8347
rect 16758 8344 16764 8356
rect 16154 8316 16764 8344
rect 16154 8313 16166 8316
rect 16108 8307 16166 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 19720 8344 19748 8375
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 18840 8316 19748 8344
rect 18840 8304 18846 8316
rect 14323 8248 15792 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 17126 8236 17132 8288
rect 17184 8276 17190 8288
rect 17221 8279 17279 8285
rect 17221 8276 17233 8279
rect 17184 8248 17233 8276
rect 17184 8236 17190 8248
rect 17221 8245 17233 8248
rect 17267 8245 17279 8279
rect 17221 8239 17279 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9306 8072 9312 8084
rect 8352 8044 8708 8072
rect 9267 8044 9312 8072
rect 8352 8032 8358 8044
rect 8570 8004 8576 8016
rect 7944 7976 8576 8004
rect 7944 7945 7972 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 8680 8004 8708 8044
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 11054 8072 11060 8084
rect 10643 8044 11060 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 13078 8032 13084 8084
rect 13136 8072 13142 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 13136 8044 13185 8072
rect 13136 8032 13142 8044
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 13173 8035 13231 8041
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 16850 8072 16856 8084
rect 16255 8044 16856 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 19245 8075 19303 8081
rect 19245 8041 19257 8075
rect 19291 8072 19303 8075
rect 19797 8075 19855 8081
rect 19797 8072 19809 8075
rect 19291 8044 19809 8072
rect 19291 8041 19303 8044
rect 19245 8035 19303 8041
rect 19797 8041 19809 8044
rect 19843 8041 19855 8075
rect 19797 8035 19855 8041
rect 10965 8007 11023 8013
rect 10965 8004 10977 8007
rect 8680 7976 10977 8004
rect 10965 7973 10977 7976
rect 11011 7973 11023 8007
rect 16577 8007 16635 8013
rect 16577 8004 16589 8007
rect 10965 7967 11023 7973
rect 11256 7976 16589 8004
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8196 7939 8254 7945
rect 8196 7905 8208 7939
rect 8242 7936 8254 7939
rect 9214 7936 9220 7948
rect 8242 7908 9220 7936
rect 8242 7905 8254 7908
rect 8196 7899 8254 7905
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 11054 7868 11060 7880
rect 11015 7840 11060 7868
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 11164 7800 11192 7831
rect 11020 7772 11192 7800
rect 11020 7760 11026 7772
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 11256 7732 11284 7976
rect 16577 7973 16589 7976
rect 16623 7973 16635 8007
rect 16577 7967 16635 7973
rect 16669 8007 16727 8013
rect 16669 7973 16681 8007
rect 16715 8004 16727 8007
rect 16942 8004 16948 8016
rect 16715 7976 16948 8004
rect 16715 7973 16727 7976
rect 16669 7967 16727 7973
rect 16942 7964 16948 7976
rect 17000 8004 17006 8016
rect 17497 8007 17555 8013
rect 17000 7976 17448 8004
rect 17000 7964 17006 7976
rect 12066 7945 12072 7948
rect 12060 7936 12072 7945
rect 12027 7908 12072 7936
rect 12060 7899 12072 7908
rect 12066 7896 12072 7899
rect 12124 7896 12130 7948
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 13446 7936 13452 7948
rect 12492 7908 13452 7936
rect 12492 7896 12498 7908
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13716 7939 13774 7945
rect 13716 7905 13728 7939
rect 13762 7936 13774 7939
rect 17126 7936 17132 7948
rect 13762 7908 17132 7936
rect 13762 7905 13774 7908
rect 13716 7899 13774 7905
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7905 17279 7939
rect 17420 7936 17448 7976
rect 17497 7973 17509 8007
rect 17543 8004 17555 8007
rect 17678 8004 17684 8016
rect 17543 7976 17684 8004
rect 17543 7973 17555 7976
rect 17497 7967 17555 7973
rect 17678 7964 17684 7976
rect 17736 7964 17742 8016
rect 19153 8007 19211 8013
rect 19153 7973 19165 8007
rect 19199 8004 19211 8007
rect 20901 8007 20959 8013
rect 20901 8004 20913 8007
rect 19199 7976 20913 8004
rect 19199 7973 19211 7976
rect 19153 7967 19211 7973
rect 20901 7973 20913 7976
rect 20947 7973 20959 8007
rect 20901 7967 20959 7973
rect 17586 7936 17592 7948
rect 17420 7908 17592 7936
rect 17221 7899 17279 7905
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 4764 7704 11284 7732
rect 11808 7732 11836 7831
rect 16758 7828 16764 7880
rect 16816 7868 16822 7880
rect 16816 7840 16861 7868
rect 16816 7828 16822 7840
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 17236 7800 17264 7899
rect 17586 7896 17592 7908
rect 17644 7896 17650 7948
rect 19610 7896 19616 7948
rect 19668 7936 19674 7948
rect 19886 7936 19892 7948
rect 19668 7908 19892 7936
rect 19668 7896 19674 7908
rect 19886 7896 19892 7908
rect 19944 7936 19950 7948
rect 20165 7939 20223 7945
rect 20165 7936 20177 7939
rect 19944 7908 20177 7936
rect 19944 7896 19950 7908
rect 20165 7905 20177 7908
rect 20211 7905 20223 7939
rect 20165 7899 20223 7905
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 18932 7840 19349 7868
rect 18932 7828 18938 7840
rect 19337 7837 19349 7840
rect 19383 7837 19395 7871
rect 20254 7868 20260 7880
rect 20215 7840 20260 7868
rect 19337 7831 19395 7837
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 20438 7868 20444 7880
rect 20399 7840 20444 7868
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 15252 7772 17264 7800
rect 15252 7760 15258 7772
rect 12434 7732 12440 7744
rect 11808 7704 12440 7732
rect 4764 7692 4770 7704
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14516 7704 14841 7732
rect 14516 7692 14522 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 14829 7695 14887 7701
rect 18690 7692 18696 7744
rect 18748 7732 18754 7744
rect 18785 7735 18843 7741
rect 18785 7732 18797 7735
rect 18748 7704 18797 7732
rect 18748 7692 18754 7704
rect 18785 7701 18797 7704
rect 18831 7701 18843 7735
rect 18785 7695 18843 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11057 7531 11115 7537
rect 11057 7528 11069 7531
rect 10928 7500 11069 7528
rect 10928 7488 10934 7500
rect 11057 7497 11069 7500
rect 11103 7497 11115 7531
rect 11057 7491 11115 7497
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11698 7528 11704 7540
rect 11379 7500 11704 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 12802 7528 12808 7540
rect 12763 7500 12808 7528
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 16206 7528 16212 7540
rect 15304 7500 16212 7528
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 12768 7364 13369 7392
rect 12768 7352 12774 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13504 7364 13829 7392
rect 13504 7352 13510 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 11241 7327 11299 7333
rect 11241 7293 11253 7327
rect 11287 7324 11299 7327
rect 13906 7324 13912 7336
rect 11287 7296 13912 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 14084 7327 14142 7333
rect 14084 7293 14096 7327
rect 14130 7324 14142 7327
rect 15304 7324 15332 7500
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 19613 7463 19671 7469
rect 19613 7429 19625 7463
rect 19659 7460 19671 7463
rect 20714 7460 20720 7472
rect 19659 7432 20720 7460
rect 19659 7429 19671 7432
rect 19613 7423 19671 7429
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20346 7392 20352 7404
rect 20303 7364 20352 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 14130 7296 15332 7324
rect 15381 7327 15439 7333
rect 14130 7293 14142 7296
rect 14084 7287 14142 7293
rect 15381 7293 15393 7327
rect 15427 7324 15439 7327
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15427 7296 15485 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 15562 7284 15568 7336
rect 15620 7324 15626 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 15620 7296 17325 7324
rect 15620 7284 15626 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 12342 7256 12348 7268
rect 11747 7228 12348 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 13173 7259 13231 7265
rect 13173 7256 13185 7259
rect 12676 7228 13185 7256
rect 12676 7216 12682 7228
rect 13173 7225 13185 7228
rect 13219 7225 13231 7259
rect 15718 7259 15776 7265
rect 15718 7256 15730 7259
rect 13173 7219 13231 7225
rect 15212 7228 15730 7256
rect 11790 7188 11796 7200
rect 11751 7160 11796 7188
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 13262 7188 13268 7200
rect 13223 7160 13268 7188
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 15212 7197 15240 7228
rect 15718 7225 15730 7228
rect 15764 7256 15776 7259
rect 15838 7256 15844 7268
rect 15764 7228 15844 7256
rect 15764 7225 15776 7228
rect 15718 7219 15776 7225
rect 15838 7216 15844 7228
rect 15896 7216 15902 7268
rect 17586 7216 17592 7268
rect 17644 7256 17650 7268
rect 19981 7259 20039 7265
rect 19981 7256 19993 7259
rect 17644 7228 19993 7256
rect 17644 7216 17650 7228
rect 19981 7225 19993 7228
rect 20027 7225 20039 7259
rect 19981 7219 20039 7225
rect 15197 7191 15255 7197
rect 15197 7157 15209 7191
rect 15243 7157 15255 7191
rect 15197 7151 15255 7157
rect 15381 7191 15439 7197
rect 15381 7157 15393 7191
rect 15427 7188 15439 7191
rect 15930 7188 15936 7200
rect 15427 7160 15936 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16850 7188 16856 7200
rect 16811 7160 16856 7188
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 17129 7191 17187 7197
rect 17129 7157 17141 7191
rect 17175 7188 17187 7191
rect 17954 7188 17960 7200
rect 17175 7160 17960 7188
rect 17175 7157 17187 7160
rect 17129 7151 17187 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 20070 7148 20076 7200
rect 20128 7188 20134 7200
rect 20128 7160 20173 7188
rect 20128 7148 20134 7160
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 12066 6984 12072 6996
rect 12027 6956 12072 6984
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 12342 6984 12348 6996
rect 12303 6956 12348 6984
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 14553 6987 14611 6993
rect 14553 6953 14565 6987
rect 14599 6984 14611 6987
rect 15289 6987 15347 6993
rect 15289 6984 15301 6987
rect 14599 6956 15301 6984
rect 14599 6953 14611 6956
rect 14553 6947 14611 6953
rect 15289 6953 15301 6956
rect 15335 6953 15347 6987
rect 20070 6984 20076 6996
rect 15289 6947 15347 6953
rect 16776 6956 20076 6984
rect 1210 6876 1216 6928
rect 1268 6916 1274 6928
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 1268 6888 13185 6916
rect 1268 6876 1274 6888
rect 13173 6885 13185 6888
rect 13219 6885 13231 6919
rect 13173 6879 13231 6885
rect 13262 6876 13268 6928
rect 13320 6916 13326 6928
rect 16776 6916 16804 6956
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 20346 6916 20352 6928
rect 13320 6888 16804 6916
rect 19352 6888 20352 6916
rect 13320 6876 13326 6888
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10962 6857 10968 6860
rect 10376 6820 10732 6848
rect 10376 6808 10382 6820
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10704 6789 10732 6820
rect 10956 6811 10968 6857
rect 11020 6848 11026 6860
rect 11020 6820 11056 6848
rect 10962 6808 10968 6811
rect 11020 6808 11026 6820
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 15654 6848 15660 6860
rect 13136 6820 13400 6848
rect 15615 6820 15660 6848
rect 13136 6808 13142 6820
rect 13372 6789 13400 6820
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 16557 6851 16615 6857
rect 16557 6848 16569 6851
rect 15804 6820 15849 6848
rect 16040 6820 16569 6848
rect 15804 6808 15810 6820
rect 10689 6783 10747 6789
rect 10284 6752 10329 6780
rect 10284 6740 10290 6752
rect 10689 6749 10701 6783
rect 10735 6749 10747 6783
rect 10689 6743 10747 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 14642 6780 14648 6792
rect 14603 6752 14648 6780
rect 13357 6743 13415 6749
rect 9674 6712 9680 6724
rect 9635 6684 9680 6712
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 10704 6644 10732 6743
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6749 14887 6783
rect 15838 6780 15844 6792
rect 15799 6752 15844 6780
rect 14829 6743 14887 6749
rect 12805 6715 12863 6721
rect 12805 6681 12817 6715
rect 12851 6712 12863 6715
rect 13170 6712 13176 6724
rect 12851 6684 13176 6712
rect 12851 6681 12863 6684
rect 12805 6675 12863 6681
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 14844 6712 14872 6743
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 16040 6712 16068 6820
rect 16557 6817 16569 6820
rect 16603 6848 16615 6851
rect 16850 6848 16856 6860
rect 16603 6820 16856 6848
rect 16603 6817 16615 6820
rect 16557 6811 16615 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 18224 6851 18282 6857
rect 18224 6848 18236 6851
rect 17696 6820 18236 6848
rect 16301 6783 16359 6789
rect 16301 6749 16313 6783
rect 16347 6749 16359 6783
rect 16301 6743 16359 6749
rect 14844 6684 16068 6712
rect 11606 6644 11612 6656
rect 10704 6616 11612 6644
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 15194 6644 15200 6656
rect 14231 6616 15200 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16316 6644 16344 6743
rect 17696 6721 17724 6820
rect 18224 6817 18236 6820
rect 18270 6848 18282 6851
rect 19352 6848 19380 6888
rect 20346 6876 20352 6888
rect 20404 6876 20410 6928
rect 19978 6848 19984 6860
rect 18270 6820 19380 6848
rect 19939 6820 19984 6848
rect 18270 6817 18282 6820
rect 18224 6811 18282 6817
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 17954 6780 17960 6792
rect 17867 6752 17960 6780
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 20070 6780 20076 6792
rect 20031 6752 20076 6780
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 20220 6752 20265 6780
rect 20220 6740 20226 6752
rect 17681 6715 17739 6721
rect 17681 6681 17693 6715
rect 17727 6681 17739 6715
rect 17681 6675 17739 6681
rect 17034 6644 17040 6656
rect 15988 6616 17040 6644
rect 15988 6604 15994 6616
rect 17034 6604 17040 6616
rect 17092 6644 17098 6656
rect 17972 6644 18000 6740
rect 19613 6715 19671 6721
rect 19613 6681 19625 6715
rect 19659 6712 19671 6715
rect 19702 6712 19708 6724
rect 19659 6684 19708 6712
rect 19659 6681 19671 6684
rect 19613 6675 19671 6681
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 18874 6644 18880 6656
rect 17092 6616 18880 6644
rect 17092 6604 17098 6616
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 19337 6647 19395 6653
rect 19337 6613 19349 6647
rect 19383 6644 19395 6647
rect 20898 6644 20904 6656
rect 19383 6616 20904 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 10873 6443 10931 6449
rect 10873 6409 10885 6443
rect 10919 6440 10931 6443
rect 10962 6440 10968 6452
rect 10919 6412 10968 6440
rect 10919 6409 10931 6412
rect 10873 6403 10931 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11790 6440 11796 6452
rect 11195 6412 11796 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 14182 6440 14188 6452
rect 13495 6412 14188 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 15289 6443 15347 6449
rect 15289 6440 15301 6443
rect 14700 6412 15301 6440
rect 14700 6400 14706 6412
rect 15289 6409 15301 6412
rect 15335 6409 15347 6443
rect 18966 6440 18972 6452
rect 15289 6403 15347 6409
rect 16960 6412 18972 6440
rect 10980 6304 11008 6400
rect 16960 6372 16988 6412
rect 18966 6400 18972 6412
rect 19024 6400 19030 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 20128 6412 20361 6440
rect 20128 6400 20134 6412
rect 20349 6409 20361 6412
rect 20395 6409 20407 6443
rect 20349 6403 20407 6409
rect 16224 6344 16988 6372
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 10980 6276 11713 6304
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 14366 6304 14372 6316
rect 14139 6276 14372 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6304 14887 6307
rect 15654 6304 15660 6316
rect 14875 6276 15660 6304
rect 14875 6273 14887 6276
rect 14829 6267 14887 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 15838 6304 15844 6316
rect 15799 6276 15844 6304
rect 15838 6264 15844 6276
rect 15896 6264 15902 6316
rect 16224 6304 16252 6344
rect 15948 6276 16252 6304
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 7340 6208 7849 6236
rect 7340 6196 7346 6208
rect 7837 6205 7849 6208
rect 7883 6236 7895 6239
rect 9493 6239 9551 6245
rect 9493 6236 9505 6239
rect 7883 6208 9505 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 9493 6205 9505 6208
rect 9539 6236 9551 6239
rect 9582 6236 9588 6248
rect 9539 6208 9588 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9760 6239 9818 6245
rect 9760 6236 9772 6239
rect 9692 6208 9772 6236
rect 8104 6171 8162 6177
rect 8104 6137 8116 6171
rect 8150 6168 8162 6171
rect 8662 6168 8668 6180
rect 8150 6140 8668 6168
rect 8150 6137 8162 6140
rect 8104 6131 8162 6137
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 7377 6103 7435 6109
rect 7377 6100 7389 6103
rect 6696 6072 7389 6100
rect 6696 6060 6702 6072
rect 7377 6069 7389 6072
rect 7423 6069 7435 6103
rect 7377 6063 7435 6069
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 9692 6100 9720 6208
rect 9760 6205 9772 6208
rect 9806 6236 9818 6239
rect 10226 6236 10232 6248
rect 9806 6208 10232 6236
rect 9806 6205 9818 6208
rect 9760 6199 9818 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11112 6208 11621 6236
rect 11112 6196 11118 6208
rect 11609 6205 11621 6208
rect 11655 6236 11667 6239
rect 15948 6236 15976 6276
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16356 6276 16865 6304
rect 16356 6264 16362 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 11655 6208 15976 6236
rect 11655 6205 11667 6208
rect 11609 6199 11667 6205
rect 16022 6196 16028 6248
rect 16080 6236 16086 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16080 6208 16681 6236
rect 16080 6196 16086 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 16761 6239 16819 6245
rect 16761 6205 16773 6239
rect 16807 6236 16819 6239
rect 16960 6236 16988 6344
rect 20898 6304 20904 6316
rect 19720 6276 20904 6304
rect 16807 6208 16988 6236
rect 18693 6239 18751 6245
rect 16807 6205 16819 6208
rect 16761 6199 16819 6205
rect 18693 6205 18705 6239
rect 18739 6236 18751 6239
rect 18782 6236 18788 6248
rect 18739 6208 18788 6236
rect 18739 6205 18751 6208
rect 18693 6199 18751 6205
rect 15657 6171 15715 6177
rect 15657 6137 15669 6171
rect 15703 6168 15715 6171
rect 16684 6168 16712 6199
rect 18782 6196 18788 6208
rect 18840 6196 18846 6248
rect 18960 6239 19018 6245
rect 18960 6205 18972 6239
rect 19006 6236 19018 6239
rect 19518 6236 19524 6248
rect 19006 6208 19524 6236
rect 19006 6205 19018 6208
rect 18960 6199 19018 6205
rect 19518 6196 19524 6208
rect 19576 6236 19582 6248
rect 19720 6236 19748 6276
rect 20898 6264 20904 6276
rect 20956 6264 20962 6316
rect 20714 6236 20720 6248
rect 19576 6208 19748 6236
rect 20675 6208 20720 6236
rect 19576 6196 19582 6208
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 19058 6168 19064 6180
rect 15703 6140 16344 6168
rect 16684 6140 19064 6168
rect 15703 6137 15715 6140
rect 15657 6131 15715 6137
rect 9263 6072 9720 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11204 6072 11529 6100
rect 11204 6060 11210 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 11517 6063 11575 6069
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 15749 6103 15807 6109
rect 13964 6072 14009 6100
rect 13964 6060 13970 6072
rect 15749 6069 15761 6103
rect 15795 6100 15807 6103
rect 16114 6100 16120 6112
rect 15795 6072 16120 6100
rect 15795 6069 15807 6072
rect 15749 6063 15807 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 16316 6109 16344 6140
rect 19058 6128 19064 6140
rect 19116 6128 19122 6180
rect 16301 6103 16359 6109
rect 16301 6069 16313 6103
rect 16347 6069 16359 6103
rect 16301 6063 16359 6069
rect 18233 6103 18291 6109
rect 18233 6069 18245 6103
rect 18279 6100 18291 6103
rect 19242 6100 19248 6112
rect 18279 6072 19248 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 20070 6100 20076 6112
rect 20031 6072 20076 6100
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 20162 6060 20168 6112
rect 20220 6100 20226 6112
rect 20809 6103 20867 6109
rect 20809 6100 20821 6103
rect 20220 6072 20821 6100
rect 20220 6060 20226 6072
rect 20809 6069 20821 6072
rect 20855 6069 20867 6103
rect 20809 6063 20867 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 6638 5896 6644 5908
rect 6599 5868 6644 5896
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 10042 5896 10048 5908
rect 9723 5868 10048 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10410 5896 10416 5908
rect 10371 5868 10416 5896
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 14366 5896 14372 5908
rect 12360 5868 14372 5896
rect 6733 5831 6791 5837
rect 6733 5797 6745 5831
rect 6779 5828 6791 5831
rect 8110 5828 8116 5840
rect 6779 5800 8116 5828
rect 6779 5797 6791 5800
rect 6733 5791 6791 5797
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 10870 5828 10876 5840
rect 10336 5800 10876 5828
rect 7558 5769 7564 5772
rect 7552 5760 7564 5769
rect 6932 5732 7564 5760
rect 6932 5701 6960 5732
rect 7552 5723 7564 5732
rect 7558 5720 7564 5723
rect 7616 5720 7622 5772
rect 10336 5769 10364 5800
rect 10870 5788 10876 5800
rect 10928 5788 10934 5840
rect 11692 5831 11750 5837
rect 11164 5800 11652 5828
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11054 5760 11060 5772
rect 10827 5732 11060 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5661 6975 5695
rect 7282 5692 7288 5704
rect 7243 5664 7288 5692
rect 6917 5655 6975 5661
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 10870 5692 10876 5704
rect 10831 5664 10876 5692
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 10980 5624 11008 5655
rect 10836 5596 11008 5624
rect 10836 5584 10842 5596
rect 6273 5559 6331 5565
rect 6273 5525 6285 5559
rect 6319 5556 6331 5559
rect 7650 5556 7656 5568
rect 6319 5528 7656 5556
rect 6319 5525 6331 5528
rect 6273 5519 6331 5525
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8662 5556 8668 5568
rect 8575 5528 8668 5556
rect 8662 5516 8668 5528
rect 8720 5556 8726 5568
rect 9122 5556 9128 5568
rect 8720 5528 9128 5556
rect 8720 5516 8726 5528
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 10137 5559 10195 5565
rect 10137 5556 10149 5559
rect 9732 5528 10149 5556
rect 9732 5516 9738 5528
rect 10137 5525 10149 5528
rect 10183 5556 10195 5559
rect 10318 5556 10324 5568
rect 10183 5528 10324 5556
rect 10183 5525 10195 5528
rect 10137 5519 10195 5525
rect 10318 5516 10324 5528
rect 10376 5556 10382 5568
rect 11164 5556 11192 5800
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 11514 5760 11520 5772
rect 11471 5732 11520 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 11624 5760 11652 5800
rect 11692 5797 11704 5831
rect 11738 5828 11750 5831
rect 12360 5828 12388 5868
rect 14366 5856 14372 5868
rect 14424 5896 14430 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 14424 5868 14473 5896
rect 14424 5856 14430 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5896 15347 5899
rect 15746 5896 15752 5908
rect 15335 5868 15752 5896
rect 15335 5865 15347 5868
rect 15289 5859 15347 5865
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 16301 5899 16359 5905
rect 16301 5896 16313 5899
rect 16172 5868 16313 5896
rect 16172 5856 16178 5868
rect 16301 5865 16313 5868
rect 16347 5865 16359 5899
rect 16758 5896 16764 5908
rect 16671 5868 16764 5896
rect 16301 5859 16359 5865
rect 16758 5856 16764 5868
rect 16816 5896 16822 5908
rect 18598 5896 18604 5908
rect 16816 5868 18604 5896
rect 16816 5856 16822 5868
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 19242 5896 19248 5908
rect 19203 5868 19248 5896
rect 19242 5856 19248 5868
rect 19300 5856 19306 5908
rect 11738 5800 12388 5828
rect 11738 5797 11750 5800
rect 11692 5791 11750 5797
rect 15838 5788 15844 5840
rect 15896 5828 15902 5840
rect 19337 5831 19395 5837
rect 19337 5828 19349 5831
rect 15896 5800 19349 5828
rect 15896 5788 15902 5800
rect 19337 5797 19349 5800
rect 19383 5797 19395 5831
rect 19337 5791 19395 5797
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 11624 5732 13093 5760
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 13348 5763 13406 5769
rect 13348 5729 13360 5763
rect 13394 5760 13406 5763
rect 14458 5760 14464 5772
rect 13394 5732 14464 5760
rect 13394 5729 13406 5732
rect 13348 5723 13406 5729
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5760 16727 5763
rect 18782 5760 18788 5772
rect 16715 5732 18788 5760
rect 16715 5729 16727 5732
rect 16669 5723 16727 5729
rect 18782 5720 18788 5732
rect 18840 5720 18846 5772
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 20622 5720 20628 5772
rect 20680 5720 20686 5772
rect 14734 5692 14740 5704
rect 14695 5664 14740 5692
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 16298 5692 16304 5704
rect 15979 5664 16304 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 16298 5652 16304 5664
rect 16356 5692 16362 5704
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16356 5664 16865 5692
rect 16356 5652 16362 5664
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 19518 5692 19524 5704
rect 19479 5664 19524 5692
rect 16853 5655 16911 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 18877 5627 18935 5633
rect 18877 5593 18889 5627
rect 18923 5624 18935 5627
rect 19978 5624 19984 5636
rect 18923 5596 19984 5624
rect 18923 5593 18935 5596
rect 18877 5587 18935 5593
rect 19978 5584 19984 5596
rect 20036 5584 20042 5636
rect 20254 5584 20260 5636
rect 20312 5624 20318 5636
rect 20640 5624 20668 5720
rect 20312 5596 20668 5624
rect 20312 5584 20318 5596
rect 10376 5528 11192 5556
rect 10376 5516 10382 5528
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 11664 5528 12817 5556
rect 11664 5516 11670 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 12805 5519 12863 5525
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 20441 5559 20499 5565
rect 20441 5556 20453 5559
rect 19484 5528 20453 5556
rect 19484 5516 19490 5528
rect 20441 5525 20453 5528
rect 20487 5525 20499 5559
rect 20441 5519 20499 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 7616 5324 8217 5352
rect 7616 5312 7622 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 12989 5355 13047 5361
rect 12989 5321 13001 5355
rect 13035 5352 13047 5355
rect 13814 5352 13820 5364
rect 13035 5324 13820 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 13964 5324 14013 5352
rect 13964 5312 13970 5324
rect 14001 5321 14013 5324
rect 14047 5321 14059 5355
rect 14001 5315 14059 5321
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 17862 5352 17868 5364
rect 15804 5324 17868 5352
rect 15804 5312 15810 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 19150 5352 19156 5364
rect 18095 5324 19156 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 20162 5352 20168 5364
rect 19659 5324 20168 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 8110 5244 8116 5296
rect 8168 5284 8174 5296
rect 8481 5287 8539 5293
rect 8481 5284 8493 5287
rect 8168 5256 8493 5284
rect 8168 5244 8174 5256
rect 8481 5253 8493 5256
rect 8527 5253 8539 5287
rect 8481 5247 8539 5253
rect 15286 5244 15292 5296
rect 15344 5284 15350 5296
rect 19334 5284 19340 5296
rect 15344 5256 19340 5284
rect 15344 5244 15350 5256
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 9030 5216 9036 5228
rect 8991 5188 9036 5216
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14458 5216 14464 5228
rect 13679 5188 14464 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 14458 5176 14464 5188
rect 14516 5216 14522 5228
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 14516 5188 14565 5216
rect 14516 5176 14522 5188
rect 14553 5185 14565 5188
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 17828 5188 18613 5216
rect 17828 5176 17834 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 19886 5216 19892 5228
rect 18601 5179 18659 5185
rect 18708 5188 19892 5216
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7092 5151 7150 5157
rect 7092 5117 7104 5151
rect 7138 5148 7150 5151
rect 9048 5148 9076 5176
rect 7138 5120 9076 5148
rect 10229 5151 10287 5157
rect 7138 5117 7150 5120
rect 7092 5111 7150 5117
rect 10229 5117 10241 5151
rect 10275 5148 10287 5151
rect 10318 5148 10324 5160
rect 10275 5120 10324 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 6270 5040 6276 5092
rect 6328 5080 6334 5092
rect 6840 5080 6868 5111
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11885 5151 11943 5157
rect 11885 5148 11897 5151
rect 11112 5120 11897 5148
rect 11112 5108 11118 5120
rect 11885 5117 11897 5120
rect 11931 5117 11943 5151
rect 11885 5111 11943 5117
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 14734 5148 14740 5160
rect 13403 5120 14740 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 18708 5148 18736 5188
rect 19886 5176 19892 5188
rect 19944 5176 19950 5228
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5216 20315 5219
rect 20346 5216 20352 5228
rect 20303 5188 20352 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 20346 5176 20352 5188
rect 20404 5176 20410 5228
rect 19058 5148 19064 5160
rect 17276 5120 18736 5148
rect 19019 5120 19064 5148
rect 17276 5108 17282 5120
rect 19058 5108 19064 5120
rect 19116 5108 19122 5160
rect 19334 5108 19340 5160
rect 19392 5148 19398 5160
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19392 5120 20085 5148
rect 19392 5108 19398 5120
rect 20073 5117 20085 5120
rect 20119 5117 20131 5151
rect 20622 5148 20628 5160
rect 20583 5120 20628 5148
rect 20073 5111 20131 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 7282 5080 7288 5092
rect 6328 5052 7288 5080
rect 6328 5040 6334 5052
rect 7282 5040 7288 5052
rect 7340 5040 7346 5092
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 8941 5083 8999 5089
rect 8941 5080 8953 5083
rect 8812 5052 8953 5080
rect 8812 5040 8818 5052
rect 8941 5049 8953 5052
rect 8987 5049 8999 5083
rect 8941 5043 8999 5049
rect 10496 5083 10554 5089
rect 10496 5049 10508 5083
rect 10542 5080 10554 5083
rect 11514 5080 11520 5092
rect 10542 5052 11520 5080
rect 10542 5049 10554 5052
rect 10496 5043 10554 5049
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 14369 5083 14427 5089
rect 14369 5080 14381 5083
rect 14240 5052 14381 5080
rect 14240 5040 14246 5052
rect 14369 5049 14381 5052
rect 14415 5080 14427 5083
rect 15746 5080 15752 5092
rect 14415 5052 15752 5080
rect 14415 5049 14427 5052
rect 14369 5043 14427 5049
rect 15746 5040 15752 5052
rect 15804 5040 15810 5092
rect 16942 5040 16948 5092
rect 17000 5080 17006 5092
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 17000 5052 18429 5080
rect 17000 5040 17006 5052
rect 18417 5049 18429 5052
rect 18463 5049 18475 5083
rect 18417 5043 18475 5049
rect 18509 5083 18567 5089
rect 18509 5049 18521 5083
rect 18555 5080 18567 5083
rect 19702 5080 19708 5092
rect 18555 5052 19708 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 19702 5040 19708 5052
rect 19760 5040 19766 5092
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 5500 4984 8861 5012
rect 5500 4972 5506 4984
rect 8849 4981 8861 4984
rect 8895 4981 8907 5015
rect 8849 4975 8907 4981
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 10836 4984 11621 5012
rect 10836 4972 10842 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 13446 5012 13452 5024
rect 13407 4984 13452 5012
rect 11609 4975 11667 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 14332 4984 14473 5012
rect 14332 4972 14338 4984
rect 14461 4981 14473 4984
rect 14507 5012 14519 5015
rect 16758 5012 16764 5024
rect 14507 4984 16764 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 19245 5015 19303 5021
rect 19245 4981 19257 5015
rect 19291 5012 19303 5015
rect 19518 5012 19524 5024
rect 19291 4984 19524 5012
rect 19291 4981 19303 4984
rect 19245 4975 19303 4981
rect 19518 4972 19524 4984
rect 19576 4972 19582 5024
rect 19610 4972 19616 5024
rect 19668 5012 19674 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19668 4984 19993 5012
rect 19668 4972 19674 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 19981 4975 20039 4981
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 20809 5015 20867 5021
rect 20809 5012 20821 5015
rect 20772 4984 20821 5012
rect 20772 4972 20778 4984
rect 20809 4981 20821 4984
rect 20855 4981 20867 5015
rect 20809 4975 20867 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 9030 4808 9036 4820
rect 7699 4780 9036 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 10597 4811 10655 4817
rect 10597 4777 10609 4811
rect 10643 4808 10655 4811
rect 10870 4808 10876 4820
rect 10643 4780 10876 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 14182 4808 14188 4820
rect 14143 4780 14188 4808
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 14274 4768 14280 4820
rect 14332 4808 14338 4820
rect 14332 4780 14377 4808
rect 14332 4768 14338 4780
rect 18598 4768 18604 4820
rect 18656 4808 18662 4820
rect 20346 4808 20352 4820
rect 18656 4780 20352 4808
rect 18656 4768 18662 4780
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 6540 4743 6598 4749
rect 6540 4709 6552 4743
rect 6586 4740 6598 4743
rect 10778 4740 10784 4752
rect 6586 4712 10784 4740
rect 6586 4709 6598 4712
rect 6540 4703 6598 4709
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 17954 4740 17960 4752
rect 17052 4712 17960 4740
rect 17052 4684 17080 4712
rect 17954 4700 17960 4712
rect 18012 4740 18018 4752
rect 19420 4743 19478 4749
rect 18012 4712 19196 4740
rect 18012 4700 18018 4712
rect 6270 4672 6276 4684
rect 6231 4644 6276 4672
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 8938 4672 8944 4684
rect 8899 4644 8944 4672
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9033 4675 9091 4681
rect 9033 4641 9045 4675
rect 9079 4672 9091 4675
rect 9950 4672 9956 4684
rect 9079 4644 9956 4672
rect 9079 4641 9091 4644
rect 9033 4635 9091 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10244 4644 10977 4672
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9180 4576 9225 4604
rect 9180 4564 9186 4576
rect 8573 4539 8631 4545
rect 8573 4505 8585 4539
rect 8619 4536 8631 4539
rect 10134 4536 10140 4548
rect 8619 4508 10140 4536
rect 8619 4505 8631 4508
rect 8573 4499 8631 4505
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 10244 4468 10272 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 17034 4672 17040 4684
rect 15252 4644 17040 4672
rect 15252 4632 15258 4644
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 17310 4681 17316 4684
rect 17304 4635 17316 4681
rect 17368 4672 17374 4684
rect 19168 4681 19196 4712
rect 19420 4709 19432 4743
rect 19466 4740 19478 4743
rect 20070 4740 20076 4752
rect 19466 4712 20076 4740
rect 19466 4709 19478 4712
rect 19420 4703 19478 4709
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 19153 4675 19211 4681
rect 17368 4644 17404 4672
rect 17310 4632 17316 4635
rect 17368 4632 17374 4644
rect 19153 4641 19165 4675
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 10594 4564 10600 4616
rect 10652 4604 10658 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10652 4576 11069 4604
rect 10652 4564 10658 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4604 11299 4607
rect 11606 4604 11612 4616
rect 11287 4576 11612 4604
rect 11287 4573 11299 4576
rect 11241 4567 11299 4573
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 13814 4468 13820 4480
rect 4212 4440 10272 4468
rect 13775 4440 13820 4468
rect 4212 4428 4218 4440
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 17828 4440 18429 4468
rect 17828 4428 17834 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 20530 4468 20536 4480
rect 20491 4440 20536 4468
rect 18417 4431 18475 4437
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 13446 4264 13452 4276
rect 9824 4236 13452 4264
rect 9824 4224 9830 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 16942 4264 16948 4276
rect 16903 4236 16948 4264
rect 16942 4224 16948 4236
rect 17000 4224 17006 4276
rect 19429 4267 19487 4273
rect 19429 4264 19441 4267
rect 17512 4236 19441 4264
rect 9232 4196 9260 4224
rect 13906 4196 13912 4208
rect 9232 4168 9987 4196
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7340 4100 7849 4128
rect 7340 4088 7346 4100
rect 7837 4097 7849 4100
rect 7883 4097 7895 4131
rect 9766 4128 9772 4140
rect 7837 4091 7895 4097
rect 8864 4100 9772 4128
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 8864 4060 8892 4100
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9959 4128 9987 4168
rect 12360 4168 13912 4196
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9959 4100 10057 4128
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10744 4100 11069 4128
rect 10744 4088 10750 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 9950 4060 9956 4072
rect 4028 4032 8892 4060
rect 9863 4032 9956 4060
rect 4028 4020 4034 4032
rect 9950 4020 9956 4032
rect 10008 4060 10014 4072
rect 12360 4060 12388 4168
rect 13906 4156 13912 4168
rect 13964 4156 13970 4208
rect 17310 4156 17316 4208
rect 17368 4196 17374 4208
rect 17512 4196 17540 4236
rect 19429 4233 19441 4236
rect 19475 4233 19487 4267
rect 19702 4264 19708 4276
rect 19663 4236 19708 4264
rect 19429 4227 19487 4233
rect 17368 4168 17540 4196
rect 17368 4156 17374 4168
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13170 4088 13176 4140
rect 13228 4128 13234 4140
rect 13228 4100 13952 4128
rect 13228 4088 13234 4100
rect 10008 4032 12388 4060
rect 12989 4063 13047 4069
rect 10008 4020 10014 4032
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13814 4060 13820 4072
rect 13035 4032 13820 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 13924 4060 13952 4100
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14332 4100 14657 4128
rect 14332 4088 14338 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 15194 4128 15200 4140
rect 15155 4100 15200 4128
rect 14645 4091 14703 4097
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 17512 4137 17540 4168
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4097 17555 4131
rect 18046 4128 18052 4140
rect 18007 4100 18052 4128
rect 17497 4091 17555 4097
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 19444 4128 19472 4227
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 19444 4100 20269 4128
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 22462 4128 22468 4140
rect 20864 4100 22468 4128
rect 20864 4088 20870 4100
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 15286 4060 15292 4072
rect 13924 4032 15292 4060
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 15464 4063 15522 4069
rect 15464 4029 15476 4063
rect 15510 4060 15522 4063
rect 17770 4060 17776 4072
rect 15510 4032 17776 4060
rect 15510 4029 15522 4032
rect 15464 4023 15522 4029
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 19426 4060 19432 4072
rect 18656 4032 19432 4060
rect 18656 4020 18662 4032
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 20680 4032 20729 4060
rect 20680 4020 20686 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 8104 3995 8162 4001
rect 8104 3961 8116 3995
rect 8150 3992 8162 3995
rect 8478 3992 8484 4004
rect 8150 3964 8484 3992
rect 8150 3961 8162 3964
rect 8104 3955 8162 3961
rect 8478 3952 8484 3964
rect 8536 3952 8542 4004
rect 9861 3995 9919 4001
rect 9861 3992 9873 3995
rect 8588 3964 9873 3992
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 5442 3924 5448 3936
rect 2924 3896 5448 3924
rect 2924 3884 2930 3896
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 8588 3924 8616 3964
rect 9861 3961 9873 3964
rect 9907 3961 9919 3995
rect 17862 3992 17868 4004
rect 9861 3955 9919 3961
rect 10336 3964 17868 3992
rect 9490 3924 9496 3936
rect 6696 3896 8616 3924
rect 9451 3896 9496 3924
rect 6696 3884 6702 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 10336 3924 10364 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 18322 4001 18328 4004
rect 18316 3992 18328 4001
rect 18283 3964 18328 3992
rect 18316 3955 18328 3964
rect 18322 3952 18328 3955
rect 18380 3952 18386 4004
rect 18414 3952 18420 4004
rect 18472 3992 18478 4004
rect 18472 3964 20944 3992
rect 18472 3952 18478 3964
rect 10502 3924 10508 3936
rect 9640 3896 10364 3924
rect 10463 3896 10508 3924
rect 9640 3884 9646 3896
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10870 3924 10876 3936
rect 10831 3896 10876 3924
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11020 3896 11065 3924
rect 11020 3884 11026 3896
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11756 3896 11805 3924
rect 11756 3884 11762 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 12526 3924 12532 3936
rect 12487 3896 12532 3924
rect 11793 3887 11851 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14458 3924 14464 3936
rect 14419 3896 14464 3924
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14553 3927 14611 3933
rect 14553 3893 14565 3927
rect 14599 3924 14611 3927
rect 15102 3924 15108 3936
rect 14599 3896 15108 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 16482 3884 16488 3936
rect 16540 3924 16546 3936
rect 16577 3927 16635 3933
rect 16577 3924 16589 3927
rect 16540 3896 16589 3924
rect 16540 3884 16546 3896
rect 16577 3893 16589 3896
rect 16623 3893 16635 3927
rect 16577 3887 16635 3893
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 17092 3896 17325 3924
rect 17092 3884 17098 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 17313 3887 17371 3893
rect 17405 3927 17463 3933
rect 17405 3893 17417 3927
rect 17451 3924 17463 3927
rect 17494 3924 17500 3936
rect 17451 3896 17500 3924
rect 17451 3893 17463 3896
rect 17405 3887 17463 3893
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 18966 3884 18972 3936
rect 19024 3924 19030 3936
rect 19702 3924 19708 3936
rect 19024 3896 19708 3924
rect 19024 3884 19030 3896
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20916 3933 20944 3964
rect 20901 3927 20959 3933
rect 20220 3896 20265 3924
rect 20220 3884 20226 3896
rect 20901 3893 20913 3927
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 4154 3720 4160 3732
rect 3476 3692 4160 3720
rect 3476 3680 3482 3692
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 6086 3680 6092 3732
rect 6144 3720 6150 3732
rect 8294 3720 8300 3732
rect 6144 3692 8300 3720
rect 6144 3680 6150 3692
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 8478 3680 8484 3692
rect 8536 3720 8542 3732
rect 9030 3720 9036 3732
rect 8536 3692 9036 3720
rect 8536 3680 8542 3692
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9125 3723 9183 3729
rect 9125 3689 9137 3723
rect 9171 3720 9183 3723
rect 10870 3720 10876 3732
rect 9171 3692 10876 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 12713 3723 12771 3729
rect 12713 3720 12725 3723
rect 11164 3692 12725 3720
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 9944 3655 10002 3661
rect 6788 3624 8340 3652
rect 6788 3612 6794 3624
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6880 3556 7113 3584
rect 6880 3544 6886 3556
rect 7101 3553 7113 3556
rect 7147 3584 7159 3587
rect 7190 3584 7196 3596
rect 7147 3556 7196 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7368 3587 7426 3593
rect 7368 3553 7380 3587
rect 7414 3584 7426 3587
rect 8202 3584 8208 3596
rect 7414 3556 8208 3584
rect 7414 3553 7426 3556
rect 7368 3547 7426 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8312 3584 8340 3624
rect 9944 3621 9956 3655
rect 9990 3652 10002 3655
rect 11164 3652 11192 3692
rect 12713 3689 12725 3692
rect 12759 3720 12771 3723
rect 13078 3720 13084 3732
rect 12759 3692 13084 3720
rect 12759 3689 12771 3692
rect 12713 3683 12771 3689
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 14366 3720 14372 3732
rect 13464 3692 14372 3720
rect 9990 3624 11192 3652
rect 9990 3621 10002 3624
rect 9944 3615 10002 3621
rect 11146 3584 11152 3596
rect 8312 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11600 3587 11658 3593
rect 11600 3553 11612 3587
rect 11646 3584 11658 3587
rect 11974 3584 11980 3596
rect 11646 3556 11980 3584
rect 11646 3553 11658 3556
rect 11600 3547 11658 3553
rect 11974 3544 11980 3556
rect 12032 3584 12038 3596
rect 13464 3584 13492 3692
rect 14366 3680 14372 3692
rect 14424 3720 14430 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14424 3692 14657 3720
rect 14424 3680 14430 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 15105 3723 15163 3729
rect 15105 3689 15117 3723
rect 15151 3720 15163 3723
rect 16574 3720 16580 3732
rect 15151 3692 16580 3720
rect 15151 3689 15163 3692
rect 15105 3683 15163 3689
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 17034 3720 17040 3732
rect 16995 3692 17040 3720
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 17494 3720 17500 3732
rect 17455 3692 17500 3720
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 17862 3720 17868 3732
rect 17823 3692 17868 3720
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 17957 3723 18015 3729
rect 17957 3689 17969 3723
rect 18003 3720 18015 3723
rect 18046 3720 18052 3732
rect 18003 3692 18052 3720
rect 18003 3689 18015 3692
rect 17957 3683 18015 3689
rect 18046 3680 18052 3692
rect 18104 3720 18110 3732
rect 18966 3720 18972 3732
rect 18104 3692 18972 3720
rect 18104 3680 18110 3692
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 19076 3692 19257 3720
rect 14182 3612 14188 3664
rect 14240 3652 14246 3664
rect 18414 3652 18420 3664
rect 14240 3624 18420 3652
rect 14240 3612 14246 3624
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 19076 3652 19104 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 19429 3723 19487 3729
rect 19429 3689 19441 3723
rect 19475 3720 19487 3723
rect 20070 3720 20076 3732
rect 19475 3692 20076 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 20622 3720 20628 3732
rect 20404 3692 20628 3720
rect 20404 3680 20410 3692
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 18524 3624 19104 3652
rect 12032 3556 13492 3584
rect 13532 3587 13590 3593
rect 12032 3544 12038 3556
rect 13532 3553 13544 3587
rect 13578 3584 13590 3587
rect 14274 3584 14280 3596
rect 13578 3556 14280 3584
rect 13578 3553 13590 3556
rect 13532 3547 13590 3553
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15252 3556 15301 3584
rect 15252 3544 15258 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15556 3587 15614 3593
rect 15556 3553 15568 3587
rect 15602 3584 15614 3587
rect 16482 3584 16488 3596
rect 15602 3556 16488 3584
rect 15602 3553 15614 3556
rect 15556 3547 15614 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 9692 3392 9720 3479
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 10928 3488 11345 3516
rect 10928 3476 10934 3488
rect 11333 3485 11345 3488
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13044 3488 13277 3516
rect 13044 3476 13050 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 18322 3516 18328 3528
rect 18187 3488 18328 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 18322 3476 18328 3488
rect 18380 3516 18386 3528
rect 18524 3516 18552 3624
rect 19150 3612 19156 3664
rect 19208 3652 19214 3664
rect 20714 3652 20720 3664
rect 19208 3624 20720 3652
rect 19208 3612 19214 3624
rect 20714 3612 20720 3624
rect 20772 3612 20778 3664
rect 18874 3584 18880 3596
rect 18835 3556 18880 3584
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 19797 3587 19855 3593
rect 19797 3584 19809 3587
rect 19300 3556 19809 3584
rect 19300 3544 19306 3556
rect 19797 3553 19809 3556
rect 19843 3553 19855 3587
rect 19797 3547 19855 3553
rect 19904 3556 20668 3584
rect 18380 3488 18552 3516
rect 18380 3476 18386 3488
rect 19702 3476 19708 3528
rect 19760 3516 19766 3528
rect 19904 3525 19932 3556
rect 19889 3519 19947 3525
rect 19889 3516 19901 3519
rect 19760 3488 19901 3516
rect 19760 3476 19766 3488
rect 19889 3485 19901 3488
rect 19935 3485 19947 3519
rect 19889 3479 19947 3485
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20530 3516 20536 3528
rect 20119 3488 20536 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 10888 3448 10916 3476
rect 10612 3420 10916 3448
rect 19245 3451 19303 3457
rect 2314 3340 2320 3392
rect 2372 3380 2378 3392
rect 8938 3380 8944 3392
rect 2372 3352 8944 3380
rect 2372 3340 2378 3352
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9674 3380 9680 3392
rect 9587 3352 9680 3380
rect 9674 3340 9680 3352
rect 9732 3380 9738 3392
rect 10318 3380 10324 3392
rect 9732 3352 10324 3380
rect 9732 3340 9738 3352
rect 10318 3340 10324 3352
rect 10376 3380 10382 3392
rect 10612 3380 10640 3420
rect 19245 3417 19257 3451
rect 19291 3448 19303 3451
rect 19794 3448 19800 3460
rect 19291 3420 19800 3448
rect 19291 3417 19303 3420
rect 19245 3411 19303 3417
rect 19794 3408 19800 3420
rect 19852 3448 19858 3460
rect 20088 3448 20116 3479
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20640 3516 20668 3556
rect 20714 3516 20720 3528
rect 20640 3488 20720 3516
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 19852 3420 20116 3448
rect 19852 3408 19858 3420
rect 10376 3352 10640 3380
rect 10376 3340 10382 3352
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10836 3352 11069 3380
rect 10836 3340 10842 3352
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 11057 3343 11115 3349
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 15105 3383 15163 3389
rect 15105 3380 15117 3383
rect 11204 3352 15117 3380
rect 11204 3340 11210 3352
rect 15105 3349 15117 3352
rect 15151 3349 15163 3383
rect 15105 3343 15163 3349
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 15988 3352 16681 3380
rect 15988 3340 15994 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 16669 3343 16727 3349
rect 19061 3383 19119 3389
rect 19061 3349 19073 3383
rect 19107 3380 19119 3383
rect 20070 3380 20076 3392
rect 19107 3352 20076 3380
rect 19107 3349 19119 3352
rect 19061 3343 19119 3349
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 8202 3176 8208 3188
rect 8163 3148 8208 3176
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 8444 3148 8493 3176
rect 8444 3136 8450 3148
rect 8481 3145 8493 3148
rect 8527 3145 8539 3179
rect 10686 3176 10692 3188
rect 8481 3139 8539 3145
rect 8772 3148 10692 3176
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 8772 3040 8800 3148
rect 10686 3136 10692 3148
rect 10744 3176 10750 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10744 3148 10977 3176
rect 10744 3136 10750 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 12894 3176 12900 3188
rect 11379 3148 12900 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 14274 3176 14280 3188
rect 14235 3148 14280 3176
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14369 3179 14427 3185
rect 14369 3145 14381 3179
rect 14415 3176 14427 3179
rect 14737 3179 14795 3185
rect 14737 3176 14749 3179
rect 14415 3148 14749 3176
rect 14415 3145 14427 3148
rect 14369 3139 14427 3145
rect 14737 3145 14749 3148
rect 14783 3145 14795 3179
rect 15102 3176 15108 3188
rect 15063 3148 15108 3176
rect 14737 3139 14795 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 16025 3179 16083 3185
rect 16025 3145 16037 3179
rect 16071 3176 16083 3179
rect 16574 3176 16580 3188
rect 16071 3148 16580 3176
rect 16071 3145 16083 3148
rect 16025 3139 16083 3145
rect 16574 3136 16580 3148
rect 16632 3176 16638 3188
rect 19334 3176 19340 3188
rect 16632 3148 19340 3176
rect 16632 3136 16638 3148
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19429 3179 19487 3185
rect 19429 3145 19441 3179
rect 19475 3176 19487 3179
rect 20162 3176 20168 3188
rect 19475 3148 20168 3176
rect 19475 3145 19487 3148
rect 19429 3139 19487 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 8846 3068 8852 3120
rect 8904 3068 8910 3120
rect 10870 3068 10876 3120
rect 10928 3108 10934 3120
rect 10928 3080 12940 3108
rect 10928 3068 10934 3080
rect 8312 3012 8800 3040
rect 1762 2932 1768 2984
rect 1820 2972 1826 2984
rect 6730 2972 6736 2984
rect 1820 2944 6736 2972
rect 1820 2932 1826 2944
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 7092 2975 7150 2981
rect 7092 2941 7104 2975
rect 7138 2972 7150 2975
rect 8312 2972 8340 3012
rect 8864 2981 8892 3068
rect 9030 3040 9036 3052
rect 8991 3012 9036 3040
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 11974 3040 11980 3052
rect 10652 3012 11836 3040
rect 11935 3012 11980 3040
rect 10652 3000 10658 3012
rect 7138 2944 8340 2972
rect 8849 2975 8907 2981
rect 7138 2941 7150 2944
rect 7092 2935 7150 2941
rect 8849 2941 8861 2975
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 9585 2975 9643 2981
rect 9585 2941 9597 2975
rect 9631 2972 9643 2975
rect 9674 2972 9680 2984
rect 9631 2944 9680 2972
rect 9631 2941 9643 2944
rect 9585 2935 9643 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9852 2975 9910 2981
rect 9852 2941 9864 2975
rect 9898 2972 9910 2975
rect 10778 2972 10784 2984
rect 9898 2944 10784 2972
rect 9898 2941 9910 2944
rect 9852 2935 9910 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11698 2972 11704 2984
rect 11659 2944 11704 2972
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 11808 2972 11836 3012
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12912 2981 12940 3080
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 13964 3080 16151 3108
rect 13964 3068 13970 3080
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 13924 3012 15761 3040
rect 12897 2975 12955 2981
rect 11808 2944 12848 2972
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8941 2907 8999 2913
rect 8941 2904 8953 2907
rect 8352 2876 8953 2904
rect 8352 2864 8358 2876
rect 8941 2873 8953 2876
rect 8987 2873 8999 2907
rect 11790 2904 11796 2916
rect 11751 2876 11796 2904
rect 8941 2867 8999 2873
rect 11790 2864 11796 2876
rect 11848 2864 11854 2916
rect 12618 2904 12624 2916
rect 11900 2876 12624 2904
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 11900 2836 11928 2876
rect 12618 2864 12624 2876
rect 12676 2864 12682 2916
rect 5684 2808 11928 2836
rect 5684 2796 5690 2808
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12820 2836 12848 2944
rect 12897 2941 12909 2975
rect 12943 2972 12955 2975
rect 12986 2972 12992 2984
rect 12943 2944 12992 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 12986 2932 12992 2944
rect 13044 2932 13050 2984
rect 13164 2975 13222 2981
rect 13164 2941 13176 2975
rect 13210 2972 13222 2975
rect 13630 2972 13636 2984
rect 13210 2944 13636 2972
rect 13210 2941 13222 2944
rect 13164 2935 13222 2941
rect 13630 2932 13636 2944
rect 13688 2972 13694 2984
rect 13924 2972 13952 3012
rect 15749 3009 15761 3012
rect 15795 3040 15807 3043
rect 15930 3040 15936 3052
rect 15795 3012 15936 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 14550 2972 14556 2984
rect 13688 2944 13952 2972
rect 14511 2944 14556 2972
rect 13688 2932 13694 2944
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15304 2944 16037 2972
rect 13722 2864 13728 2916
rect 13780 2904 13786 2916
rect 14369 2907 14427 2913
rect 14369 2904 14381 2907
rect 13780 2876 14381 2904
rect 13780 2864 13786 2876
rect 14369 2873 14381 2876
rect 14415 2873 14427 2907
rect 14369 2867 14427 2873
rect 15304 2836 15332 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16123 2972 16151 3080
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 18233 3111 18291 3117
rect 18233 3108 18245 3111
rect 17092 3080 18245 3108
rect 17092 3068 17098 3080
rect 18233 3077 18245 3080
rect 18279 3077 18291 3111
rect 18233 3071 18291 3077
rect 18874 3068 18880 3120
rect 18932 3108 18938 3120
rect 20717 3111 20775 3117
rect 20717 3108 20729 3111
rect 18932 3080 20729 3108
rect 18932 3068 18938 3080
rect 20717 3077 20729 3080
rect 20763 3077 20775 3111
rect 20717 3071 20775 3077
rect 16206 3000 16212 3052
rect 16264 3040 16270 3052
rect 16482 3040 16488 3052
rect 16264 3012 16488 3040
rect 16264 3000 16270 3012
rect 16482 3000 16488 3012
rect 16540 3040 16546 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16540 3012 16681 3040
rect 16540 3000 16546 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 16776 3012 18828 3040
rect 16776 2972 16804 3012
rect 16123 2944 16804 2972
rect 17405 2975 17463 2981
rect 16025 2935 16083 2941
rect 15470 2836 15476 2848
rect 12492 2808 12537 2836
rect 12820 2808 15332 2836
rect 15431 2808 15476 2836
rect 12492 2796 12498 2808
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 16500 2845 16528 2944
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 17678 2972 17684 2984
rect 17451 2944 17684 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 17678 2932 17684 2944
rect 17736 2932 17742 2984
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2972 18107 2975
rect 18506 2972 18512 2984
rect 18095 2944 18512 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18506 2932 18512 2944
rect 18564 2932 18570 2984
rect 18690 2972 18696 2984
rect 18651 2944 18696 2972
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 18800 2972 18828 3012
rect 18966 3000 18972 3052
rect 19024 3040 19030 3052
rect 19242 3040 19248 3052
rect 19024 3012 19248 3040
rect 19024 3000 19030 3012
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 19794 3000 19800 3052
rect 19852 3040 19858 3052
rect 19981 3043 20039 3049
rect 19981 3040 19993 3043
rect 19852 3012 19993 3040
rect 19852 3000 19858 3012
rect 19981 3009 19993 3012
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 20438 3000 20444 3052
rect 20496 3000 20502 3052
rect 19426 2972 19432 2984
rect 18800 2944 19432 2972
rect 19426 2932 19432 2944
rect 19484 2972 19490 2984
rect 19610 2972 19616 2984
rect 19484 2944 19616 2972
rect 19484 2932 19490 2944
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 20456 2972 20484 3000
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 20456 2944 20545 2972
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 18874 2864 18880 2916
rect 18932 2904 18938 2916
rect 18969 2907 19027 2913
rect 18969 2904 18981 2907
rect 18932 2876 18981 2904
rect 18932 2864 18938 2876
rect 18969 2873 18981 2876
rect 19015 2873 19027 2907
rect 18969 2867 19027 2873
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 21358 2904 21364 2916
rect 19300 2876 21364 2904
rect 19300 2864 19306 2876
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 15565 2839 15623 2845
rect 15565 2805 15577 2839
rect 15611 2836 15623 2839
rect 16117 2839 16175 2845
rect 16117 2836 16129 2839
rect 15611 2808 16129 2836
rect 15611 2805 15623 2808
rect 15565 2799 15623 2805
rect 16117 2805 16129 2808
rect 16163 2805 16175 2839
rect 16117 2799 16175 2805
rect 16485 2839 16543 2845
rect 16485 2805 16497 2839
rect 16531 2805 16543 2839
rect 16485 2799 16543 2805
rect 16574 2796 16580 2848
rect 16632 2836 16638 2848
rect 16632 2808 16677 2836
rect 16632 2796 16638 2808
rect 17494 2796 17500 2848
rect 17552 2836 17558 2848
rect 17589 2839 17647 2845
rect 17589 2836 17601 2839
rect 17552 2808 17601 2836
rect 17552 2796 17558 2808
rect 17589 2805 17601 2808
rect 17635 2805 17647 2839
rect 19794 2836 19800 2848
rect 19755 2808 19800 2836
rect 17589 2799 17647 2805
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 19889 2839 19947 2845
rect 19889 2805 19901 2839
rect 19935 2836 19947 2839
rect 20622 2836 20628 2848
rect 19935 2808 20628 2836
rect 19935 2805 19947 2808
rect 19889 2799 19947 2805
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 8294 2632 8300 2644
rect 7423 2604 8300 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 8846 2632 8852 2644
rect 8435 2604 8852 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10962 2632 10968 2644
rect 10183 2604 10968 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 12492 2604 13369 2632
rect 12492 2592 12498 2604
rect 13357 2601 13369 2604
rect 13403 2601 13415 2635
rect 13357 2595 13415 2601
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 15841 2635 15899 2641
rect 15841 2632 15853 2635
rect 15528 2604 15853 2632
rect 15528 2592 15534 2604
rect 15841 2601 15853 2604
rect 15887 2601 15899 2635
rect 15841 2595 15899 2601
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 17586 2632 17592 2644
rect 16255 2604 17592 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 17865 2635 17923 2641
rect 17865 2601 17877 2635
rect 17911 2632 17923 2635
rect 19242 2632 19248 2644
rect 17911 2604 19248 2632
rect 17911 2601 17923 2604
rect 17865 2595 17923 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 20717 2635 20775 2641
rect 20717 2601 20729 2635
rect 20763 2601 20775 2635
rect 20717 2595 20775 2601
rect 7834 2524 7840 2576
rect 7892 2564 7898 2576
rect 10505 2567 10563 2573
rect 10505 2564 10517 2567
rect 7892 2536 10517 2564
rect 7892 2524 7898 2536
rect 10505 2533 10517 2536
rect 10551 2533 10563 2567
rect 10505 2527 10563 2533
rect 10594 2524 10600 2576
rect 10652 2564 10658 2576
rect 10652 2536 10697 2564
rect 10652 2524 10658 2536
rect 15378 2524 15384 2576
rect 15436 2564 15442 2576
rect 20732 2564 20760 2595
rect 15436 2536 20760 2564
rect 15436 2524 15442 2536
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 7248 2468 7757 2496
rect 7248 2456 7254 2468
rect 7745 2465 7757 2468
rect 7791 2465 7803 2499
rect 7745 2459 7803 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11882 2496 11888 2508
rect 11471 2468 11888 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 13998 2496 14004 2508
rect 12023 2468 14004 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 13998 2456 14004 2468
rect 14056 2456 14062 2508
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2496 16359 2499
rect 16945 2499 17003 2505
rect 16347 2468 16896 2496
rect 16347 2465 16359 2468
rect 16301 2459 16359 2465
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8202 2428 8208 2440
rect 8067 2400 8208 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 7852 2360 7880 2391
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 10778 2428 10784 2440
rect 10739 2400 10784 2428
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 10888 2400 13461 2428
rect 8294 2360 8300 2372
rect 7852 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 8846 2320 8852 2372
rect 8904 2360 8910 2372
rect 10888 2360 10916 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13630 2428 13636 2440
rect 13591 2400 13636 2428
rect 13449 2391 13507 2397
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 16393 2431 16451 2437
rect 16393 2428 16405 2431
rect 16264 2400 16405 2428
rect 16264 2388 16270 2400
rect 16393 2397 16405 2400
rect 16439 2397 16451 2431
rect 16868 2428 16896 2468
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17402 2496 17408 2508
rect 16991 2468 17408 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17402 2456 17408 2468
rect 17460 2456 17466 2508
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2496 17739 2499
rect 17954 2496 17960 2508
rect 17727 2468 17960 2496
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 18417 2499 18475 2505
rect 18417 2465 18429 2499
rect 18463 2496 18475 2499
rect 18874 2496 18880 2508
rect 18463 2468 18880 2496
rect 18463 2465 18475 2468
rect 18417 2459 18475 2465
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19116 2468 19441 2496
rect 19116 2456 19122 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 19886 2456 19892 2508
rect 19944 2496 19950 2508
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19944 2468 19993 2496
rect 19944 2456 19950 2468
rect 19981 2465 19993 2468
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 20438 2456 20444 2508
rect 20496 2496 20502 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20496 2468 20545 2496
rect 20496 2456 20502 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 17126 2428 17132 2440
rect 16868 2400 17132 2428
rect 16393 2391 16451 2397
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 8904 2332 10916 2360
rect 12989 2363 13047 2369
rect 8904 2320 8910 2332
rect 12989 2329 13001 2363
rect 13035 2360 13047 2363
rect 14458 2360 14464 2372
rect 13035 2332 14464 2360
rect 13035 2329 13047 2332
rect 12989 2323 13047 2329
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 14826 2320 14832 2372
rect 14884 2360 14890 2372
rect 19613 2363 19671 2369
rect 14884 2332 18736 2360
rect 14884 2320 14890 2332
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 12161 2295 12219 2301
rect 12161 2261 12173 2295
rect 12207 2292 12219 2295
rect 12618 2292 12624 2304
rect 12207 2264 12624 2292
rect 12207 2261 12219 2264
rect 12161 2255 12219 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 16482 2252 16488 2304
rect 16540 2292 16546 2304
rect 17129 2295 17187 2301
rect 17129 2292 17141 2295
rect 16540 2264 17141 2292
rect 16540 2252 16546 2264
rect 17129 2261 17141 2264
rect 17175 2261 17187 2295
rect 17129 2255 17187 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 18601 2295 18659 2301
rect 18601 2292 18613 2295
rect 18012 2264 18613 2292
rect 18012 2252 18018 2264
rect 18601 2261 18613 2264
rect 18647 2261 18659 2295
rect 18708 2292 18736 2332
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 20806 2360 20812 2372
rect 19659 2332 20812 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 20806 2320 20812 2332
rect 20864 2320 20870 2372
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 18708 2264 20177 2292
rect 18601 2255 18659 2261
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 8294 2048 8300 2100
rect 8352 2088 8358 2100
rect 8754 2088 8760 2100
rect 8352 2060 8760 2088
rect 8352 2048 8358 2060
rect 8754 2048 8760 2060
rect 8812 2088 8818 2100
rect 18782 2088 18788 2100
rect 8812 2060 18788 2088
rect 8812 2048 8818 2060
rect 18782 2048 18788 2060
rect 18840 2088 18846 2100
rect 19794 2088 19800 2100
rect 18840 2060 19800 2088
rect 18840 2048 18846 2060
rect 19794 2048 19800 2060
rect 19852 2048 19858 2100
rect 9950 1164 9956 1216
rect 10008 1204 10014 1216
rect 15838 1204 15844 1216
rect 10008 1176 15844 1204
rect 10008 1164 10014 1176
rect 15838 1164 15844 1176
rect 15896 1164 15902 1216
rect 10502 824 10508 876
rect 10560 864 10566 876
rect 15654 864 15660 876
rect 10560 836 15660 864
rect 10560 824 10566 836
rect 15654 824 15660 836
rect 15712 824 15718 876
rect 8294 620 8300 672
rect 8352 660 8358 672
rect 11790 660 11796 672
rect 8352 632 11796 660
rect 8352 620 8358 632
rect 11790 620 11796 632
rect 11848 620 11854 672
rect 12066 552 12072 604
rect 12124 592 12130 604
rect 15010 592 15016 604
rect 12124 564 15016 592
rect 12124 552 12130 564
rect 15010 552 15016 564
rect 15068 552 15074 604
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 20628 20000 20680 20052
rect 19892 19864 19944 19916
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 15936 19252 15988 19304
rect 17868 19252 17920 19304
rect 18880 19252 18932 19304
rect 19064 19252 19116 19304
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 5724 19184 5776 19236
rect 17776 19116 17828 19168
rect 18512 19159 18564 19168
rect 18512 19125 18521 19159
rect 18521 19125 18555 19159
rect 18555 19125 18564 19159
rect 18512 19116 18564 19125
rect 20812 19116 20864 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 15752 18844 15804 18896
rect 15936 18887 15988 18896
rect 15936 18853 15945 18887
rect 15945 18853 15979 18887
rect 15979 18853 15988 18887
rect 15936 18844 15988 18853
rect 17868 18887 17920 18896
rect 17868 18853 17877 18887
rect 17877 18853 17911 18887
rect 17911 18853 17920 18887
rect 17868 18844 17920 18853
rect 19892 18887 19944 18896
rect 19892 18853 19901 18887
rect 19901 18853 19935 18887
rect 19935 18853 19944 18887
rect 19892 18844 19944 18853
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 11704 18776 11756 18828
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 19616 18819 19668 18828
rect 19616 18785 19625 18819
rect 19625 18785 19659 18819
rect 19659 18785 19668 18819
rect 19616 18776 19668 18785
rect 19984 18640 20036 18692
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 20168 18411 20220 18420
rect 20168 18377 20177 18411
rect 20177 18377 20211 18411
rect 20211 18377 20220 18411
rect 20168 18368 20220 18377
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 15752 18232 15804 18284
rect 7656 18164 7708 18216
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 17868 17824 17920 17876
rect 20444 17867 20496 17876
rect 20444 17833 20453 17867
rect 20453 17833 20487 17867
rect 20487 17833 20496 17867
rect 20444 17824 20496 17833
rect 11888 17688 11940 17740
rect 14464 17688 14516 17740
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 14464 17187 14516 17196
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 14188 17119 14240 17128
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 19892 17076 19944 17128
rect 17316 17008 17368 17060
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 17316 16711 17368 16720
rect 17316 16677 17325 16711
rect 17325 16677 17359 16711
rect 17359 16677 17368 16711
rect 17316 16668 17368 16677
rect 19892 16711 19944 16720
rect 19892 16677 19901 16711
rect 19901 16677 19935 16711
rect 19935 16677 19944 16711
rect 19892 16668 19944 16677
rect 16396 16600 16448 16652
rect 19524 16600 19576 16652
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 20536 16031 20588 16040
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 20536 15580 20588 15632
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 13912 15555 13964 15564
rect 13912 15521 13921 15555
rect 13921 15521 13955 15555
rect 13955 15521 13964 15555
rect 13912 15512 13964 15521
rect 20260 15555 20312 15564
rect 20260 15521 20269 15555
rect 20269 15521 20303 15555
rect 20303 15521 20312 15555
rect 20260 15512 20312 15521
rect 19984 15376 20036 15428
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 9588 14943 9640 14952
rect 9588 14909 9597 14943
rect 9597 14909 9631 14943
rect 9631 14909 9640 14943
rect 9588 14900 9640 14909
rect 16488 14900 16540 14952
rect 20260 14832 20312 14884
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 19892 14603 19944 14612
rect 19892 14569 19901 14603
rect 19901 14569 19935 14603
rect 19935 14569 19944 14603
rect 19892 14560 19944 14569
rect 20444 14603 20496 14612
rect 20444 14569 20453 14603
rect 20453 14569 20487 14603
rect 20487 14569 20496 14603
rect 20444 14560 20496 14569
rect 8392 14467 8444 14476
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 16488 14356 16540 14408
rect 11060 14288 11112 14340
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 16304 14016 16356 14068
rect 19248 14016 19300 14068
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 19892 13880 19944 13932
rect 10508 13812 10560 13864
rect 16120 13855 16172 13864
rect 16120 13821 16129 13855
rect 16129 13821 16163 13855
rect 16163 13821 16172 13855
rect 16120 13812 16172 13821
rect 17132 13812 17184 13864
rect 19432 13812 19484 13864
rect 20076 13812 20128 13864
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 19248 13515 19300 13524
rect 19248 13481 19257 13515
rect 19257 13481 19291 13515
rect 19291 13481 19300 13515
rect 19248 13472 19300 13481
rect 19708 13404 19760 13456
rect 19340 13336 19392 13388
rect 12532 13268 12584 13320
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 15660 12928 15712 12980
rect 17592 12928 17644 12980
rect 19248 12971 19300 12980
rect 19248 12937 19257 12971
rect 19257 12937 19291 12971
rect 19291 12937 19300 12971
rect 19248 12928 19300 12937
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 17592 12835 17644 12844
rect 17592 12801 17601 12835
rect 17601 12801 17635 12835
rect 17635 12801 17644 12835
rect 17592 12792 17644 12801
rect 19432 12792 19484 12844
rect 14096 12724 14148 12776
rect 16488 12656 16540 12708
rect 17684 12724 17736 12776
rect 19800 12724 19852 12776
rect 19432 12656 19484 12708
rect 19892 12656 19944 12708
rect 20260 12656 20312 12708
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 17316 12631 17368 12640
rect 15568 12588 15620 12597
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 15476 12384 15528 12436
rect 20444 12427 20496 12436
rect 13452 12316 13504 12368
rect 15384 12248 15436 12300
rect 16120 12316 16172 12368
rect 20444 12393 20453 12427
rect 20453 12393 20487 12427
rect 20487 12393 20496 12427
rect 20444 12384 20496 12393
rect 16764 12248 16816 12300
rect 17592 12316 17644 12368
rect 19340 12316 19392 12368
rect 19156 12248 19208 12300
rect 20260 12291 20312 12300
rect 20260 12257 20269 12291
rect 20269 12257 20303 12291
rect 20303 12257 20312 12291
rect 20260 12248 20312 12257
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 15844 12044 15896 12096
rect 18880 12044 18932 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 15660 11840 15712 11892
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 13452 11704 13504 11756
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 17316 11704 17368 11756
rect 13636 11636 13688 11688
rect 15660 11679 15712 11688
rect 15660 11645 15694 11679
rect 15694 11645 15712 11679
rect 15660 11636 15712 11645
rect 18512 11704 18564 11756
rect 20628 11704 20680 11756
rect 18420 11636 18472 11688
rect 18880 11679 18932 11688
rect 18880 11645 18914 11679
rect 18914 11645 18932 11679
rect 18880 11636 18932 11645
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 15844 11568 15896 11620
rect 19616 11568 19668 11620
rect 13176 11500 13228 11509
rect 21916 11568 21968 11620
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 20260 11543 20312 11552
rect 20260 11509 20269 11543
rect 20269 11509 20303 11543
rect 20303 11509 20312 11543
rect 20260 11500 20312 11509
rect 20444 11500 20496 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 664 11296 716 11348
rect 4068 11228 4120 11280
rect 13636 11296 13688 11348
rect 15568 11296 15620 11348
rect 15936 11296 15988 11348
rect 19340 11296 19392 11348
rect 13084 11160 13136 11212
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 15568 11160 15620 11212
rect 15844 11135 15896 11144
rect 12440 11092 12492 11101
rect 13452 11024 13504 11076
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 18880 11228 18932 11280
rect 19984 11228 20036 11280
rect 20628 11160 20680 11212
rect 17592 10956 17644 11008
rect 18420 11092 18472 11144
rect 17960 10956 18012 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 19524 10752 19576 10804
rect 16488 10616 16540 10668
rect 16764 10616 16816 10668
rect 17960 10616 18012 10668
rect 19984 10616 20036 10668
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 20628 10659 20680 10668
rect 20628 10625 20637 10659
rect 20637 10625 20671 10659
rect 20671 10625 20680 10659
rect 20628 10616 20680 10625
rect 11980 10480 12032 10532
rect 15292 10480 15344 10532
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 16580 10548 16632 10600
rect 18052 10548 18104 10600
rect 19340 10548 19392 10600
rect 20260 10548 20312 10600
rect 16580 10412 16632 10464
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 18604 10412 18656 10464
rect 20444 10455 20496 10464
rect 20444 10421 20453 10455
rect 20453 10421 20487 10455
rect 20487 10421 20496 10455
rect 20444 10412 20496 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 13912 10208 13964 10260
rect 15752 10208 15804 10260
rect 17960 10140 18012 10192
rect 20444 10140 20496 10192
rect 12992 10072 13044 10124
rect 15384 10072 15436 10124
rect 15844 10072 15896 10124
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 19708 10115 19760 10124
rect 19708 10081 19717 10115
rect 19717 10081 19751 10115
rect 19751 10081 19760 10115
rect 19708 10072 19760 10081
rect 20352 10072 20404 10124
rect 12808 10004 12860 10056
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 18972 9979 19024 9988
rect 18972 9945 18981 9979
rect 18981 9945 19015 9979
rect 19015 9945 19024 9979
rect 18972 9936 19024 9945
rect 13728 9868 13780 9920
rect 16488 9868 16540 9920
rect 19064 9868 19116 9920
rect 19340 9868 19392 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 11888 9664 11940 9716
rect 11796 9596 11848 9648
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 10876 9460 10928 9512
rect 15384 9664 15436 9716
rect 17592 9664 17644 9716
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 10416 9392 10468 9444
rect 13728 9503 13780 9512
rect 13728 9469 13762 9503
rect 13762 9469 13780 9503
rect 11888 9392 11940 9444
rect 13728 9460 13780 9469
rect 17960 9528 18012 9580
rect 16488 9460 16540 9512
rect 17592 9460 17644 9512
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 18972 9460 19024 9512
rect 19248 9460 19300 9512
rect 15016 9392 15068 9444
rect 10324 9324 10376 9376
rect 11060 9324 11112 9376
rect 15844 9324 15896 9376
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 19800 9367 19852 9376
rect 19800 9333 19809 9367
rect 19809 9333 19843 9367
rect 19843 9333 19852 9367
rect 19800 9324 19852 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 9588 9120 9640 9172
rect 5080 9052 5132 9104
rect 13728 9120 13780 9172
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 15936 9120 15988 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 9496 8916 9548 8968
rect 9312 8848 9364 8900
rect 10324 8916 10376 8968
rect 11612 8984 11664 9036
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12716 9027 12768 9036
rect 12440 8984 12492 8993
rect 12716 8993 12750 9027
rect 12750 8993 12768 9027
rect 12716 8984 12768 8993
rect 18604 9052 18656 9104
rect 19248 9052 19300 9104
rect 19800 9052 19852 9104
rect 17500 8984 17552 9036
rect 18420 8984 18472 9036
rect 14004 8916 14056 8968
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 17132 8916 17184 8968
rect 18972 8916 19024 8968
rect 12716 8780 12768 8832
rect 13360 8780 13412 8832
rect 19432 8780 19484 8832
rect 20444 8823 20496 8832
rect 20444 8789 20453 8823
rect 20453 8789 20487 8823
rect 20487 8789 20496 8823
rect 20444 8780 20496 8789
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 10324 8372 10376 8424
rect 13360 8372 13412 8424
rect 18880 8576 18932 8628
rect 15568 8551 15620 8560
rect 15568 8517 15577 8551
rect 15577 8517 15611 8551
rect 15611 8517 15620 8551
rect 15568 8508 15620 8517
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 9312 8304 9364 8356
rect 10968 8304 11020 8356
rect 14556 8304 14608 8356
rect 13912 8236 13964 8288
rect 15936 8372 15988 8424
rect 18972 8415 19024 8424
rect 18972 8381 18981 8415
rect 18981 8381 19015 8415
rect 19015 8381 19024 8415
rect 18972 8372 19024 8381
rect 16764 8304 16816 8356
rect 18788 8304 18840 8356
rect 20444 8372 20496 8424
rect 17132 8236 17184 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 8300 8032 8352 8084
rect 9312 8075 9364 8084
rect 8576 7964 8628 8016
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 11060 8032 11112 8084
rect 13084 8032 13136 8084
rect 16856 8032 16908 8084
rect 9220 7896 9272 7948
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 10968 7760 11020 7812
rect 4712 7692 4764 7744
rect 16948 7964 17000 8016
rect 12072 7939 12124 7948
rect 12072 7905 12106 7939
rect 12106 7905 12124 7939
rect 12072 7896 12124 7905
rect 12440 7896 12492 7948
rect 13452 7939 13504 7948
rect 13452 7905 13461 7939
rect 13461 7905 13495 7939
rect 13495 7905 13504 7939
rect 13452 7896 13504 7905
rect 17132 7896 17184 7948
rect 17684 7964 17736 8016
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 15200 7760 15252 7812
rect 17592 7896 17644 7948
rect 19616 7896 19668 7948
rect 19892 7896 19944 7948
rect 18880 7828 18932 7880
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 12440 7692 12492 7744
rect 14464 7692 14516 7744
rect 18696 7692 18748 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 10876 7488 10928 7540
rect 11704 7488 11756 7540
rect 12808 7531 12860 7540
rect 12808 7497 12817 7531
rect 12817 7497 12851 7531
rect 12851 7497 12860 7531
rect 12808 7488 12860 7497
rect 12072 7352 12124 7404
rect 12716 7352 12768 7404
rect 13452 7352 13504 7404
rect 13912 7284 13964 7336
rect 16212 7488 16264 7540
rect 20720 7420 20772 7472
rect 20352 7352 20404 7404
rect 15568 7284 15620 7336
rect 12348 7216 12400 7268
rect 12624 7216 12676 7268
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 15844 7216 15896 7268
rect 17592 7216 17644 7268
rect 15936 7148 15988 7200
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 17960 7148 18012 7200
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 12072 6987 12124 6996
rect 12072 6953 12081 6987
rect 12081 6953 12115 6987
rect 12115 6953 12124 6987
rect 12072 6944 12124 6953
rect 12348 6987 12400 6996
rect 12348 6953 12357 6987
rect 12357 6953 12391 6987
rect 12391 6953 12400 6987
rect 12348 6944 12400 6953
rect 1216 6876 1268 6928
rect 13268 6919 13320 6928
rect 13268 6885 13277 6919
rect 13277 6885 13311 6919
rect 13311 6885 13320 6919
rect 20076 6944 20128 6996
rect 13268 6876 13320 6885
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10324 6808 10376 6860
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10968 6851 11020 6860
rect 10968 6817 11002 6851
rect 11002 6817 11020 6851
rect 10968 6808 11020 6817
rect 13084 6808 13136 6860
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 10232 6740 10284 6749
rect 14648 6783 14700 6792
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 14648 6749 14657 6783
rect 14657 6749 14691 6783
rect 14691 6749 14700 6783
rect 14648 6740 14700 6749
rect 15844 6783 15896 6792
rect 13176 6672 13228 6724
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 16856 6808 16908 6860
rect 11612 6604 11664 6656
rect 15200 6604 15252 6656
rect 15936 6604 15988 6656
rect 20352 6876 20404 6928
rect 19984 6851 20036 6860
rect 19984 6817 19993 6851
rect 19993 6817 20027 6851
rect 20027 6817 20036 6851
rect 19984 6808 20036 6817
rect 17960 6783 18012 6792
rect 17960 6749 17969 6783
rect 17969 6749 18003 6783
rect 18003 6749 18012 6783
rect 17960 6740 18012 6749
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 17040 6604 17092 6656
rect 19708 6672 19760 6724
rect 18880 6604 18932 6656
rect 20904 6604 20956 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 10968 6400 11020 6452
rect 11796 6400 11848 6452
rect 14188 6400 14240 6452
rect 14648 6400 14700 6452
rect 18972 6400 19024 6452
rect 20076 6400 20128 6452
rect 14372 6264 14424 6316
rect 15660 6264 15712 6316
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 7288 6196 7340 6248
rect 9588 6196 9640 6248
rect 8668 6128 8720 6180
rect 6644 6060 6696 6112
rect 10232 6196 10284 6248
rect 11060 6196 11112 6248
rect 16304 6264 16356 6316
rect 16028 6196 16080 6248
rect 20904 6307 20956 6316
rect 18788 6196 18840 6248
rect 19524 6196 19576 6248
rect 20904 6273 20913 6307
rect 20913 6273 20947 6307
rect 20947 6273 20956 6307
rect 20904 6264 20956 6273
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 11152 6060 11204 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 16120 6060 16172 6112
rect 19064 6128 19116 6180
rect 19248 6060 19300 6112
rect 20076 6103 20128 6112
rect 20076 6069 20085 6103
rect 20085 6069 20119 6103
rect 20119 6069 20128 6103
rect 20076 6060 20128 6069
rect 20168 6060 20220 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 6644 5899 6696 5908
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 10048 5856 10100 5908
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 8116 5788 8168 5840
rect 7564 5763 7616 5772
rect 7564 5729 7598 5763
rect 7598 5729 7616 5763
rect 7564 5720 7616 5729
rect 10876 5788 10928 5840
rect 11060 5720 11112 5772
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 10784 5584 10836 5636
rect 7656 5516 7708 5568
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 9128 5516 9180 5568
rect 9680 5516 9732 5568
rect 10324 5516 10376 5568
rect 11520 5720 11572 5772
rect 14372 5856 14424 5908
rect 15752 5856 15804 5908
rect 16120 5856 16172 5908
rect 16764 5899 16816 5908
rect 16764 5865 16773 5899
rect 16773 5865 16807 5899
rect 16807 5865 16816 5899
rect 16764 5856 16816 5865
rect 18604 5856 18656 5908
rect 19248 5899 19300 5908
rect 19248 5865 19257 5899
rect 19257 5865 19291 5899
rect 19291 5865 19300 5899
rect 19248 5856 19300 5865
rect 15844 5788 15896 5840
rect 14464 5720 14516 5772
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 18788 5720 18840 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 20628 5720 20680 5772
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 16304 5652 16356 5704
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 19984 5584 20036 5636
rect 20260 5584 20312 5636
rect 11612 5516 11664 5568
rect 19432 5516 19484 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 7564 5312 7616 5364
rect 13820 5312 13872 5364
rect 13912 5312 13964 5364
rect 15752 5312 15804 5364
rect 17868 5312 17920 5364
rect 19156 5312 19208 5364
rect 20168 5312 20220 5364
rect 8116 5244 8168 5296
rect 15292 5244 15344 5296
rect 19340 5244 19392 5296
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 14464 5176 14516 5228
rect 17776 5176 17828 5228
rect 6276 5040 6328 5092
rect 10324 5108 10376 5160
rect 11060 5108 11112 5160
rect 14740 5108 14792 5160
rect 17224 5108 17276 5160
rect 19892 5176 19944 5228
rect 20352 5176 20404 5228
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 19340 5108 19392 5160
rect 20628 5151 20680 5160
rect 20628 5117 20637 5151
rect 20637 5117 20671 5151
rect 20671 5117 20680 5151
rect 20628 5108 20680 5117
rect 7288 5040 7340 5092
rect 8760 5040 8812 5092
rect 11520 5040 11572 5092
rect 14188 5040 14240 5092
rect 15752 5040 15804 5092
rect 16948 5040 17000 5092
rect 19708 5040 19760 5092
rect 5448 4972 5500 5024
rect 10784 4972 10836 5024
rect 13452 5015 13504 5024
rect 13452 4981 13461 5015
rect 13461 4981 13495 5015
rect 13495 4981 13504 5015
rect 13452 4972 13504 4981
rect 14280 4972 14332 5024
rect 16764 4972 16816 5024
rect 19524 4972 19576 5024
rect 19616 4972 19668 5024
rect 20720 4972 20772 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 9036 4768 9088 4820
rect 10876 4768 10928 4820
rect 14188 4811 14240 4820
rect 14188 4777 14197 4811
rect 14197 4777 14231 4811
rect 14231 4777 14240 4811
rect 14188 4768 14240 4777
rect 14280 4811 14332 4820
rect 14280 4777 14289 4811
rect 14289 4777 14323 4811
rect 14323 4777 14332 4811
rect 14280 4768 14332 4777
rect 18604 4768 18656 4820
rect 20352 4768 20404 4820
rect 10784 4700 10836 4752
rect 17960 4700 18012 4752
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 9956 4632 10008 4684
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 10140 4496 10192 4548
rect 4160 4428 4212 4480
rect 15200 4632 15252 4684
rect 17040 4675 17092 4684
rect 17040 4641 17049 4675
rect 17049 4641 17083 4675
rect 17083 4641 17092 4675
rect 17040 4632 17092 4641
rect 17316 4675 17368 4684
rect 17316 4641 17350 4675
rect 17350 4641 17368 4675
rect 20076 4700 20128 4752
rect 17316 4632 17368 4641
rect 10600 4564 10652 4616
rect 11612 4564 11664 4616
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 13820 4471 13872 4480
rect 13820 4437 13829 4471
rect 13829 4437 13863 4471
rect 13863 4437 13872 4471
rect 13820 4428 13872 4437
rect 17776 4428 17828 4480
rect 20536 4471 20588 4480
rect 20536 4437 20545 4471
rect 20545 4437 20579 4471
rect 20579 4437 20588 4471
rect 20536 4428 20588 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 9772 4224 9824 4276
rect 13452 4224 13504 4276
rect 16948 4267 17000 4276
rect 16948 4233 16957 4267
rect 16957 4233 16991 4267
rect 16991 4233 17000 4267
rect 16948 4224 17000 4233
rect 7288 4088 7340 4140
rect 3976 4020 4028 4072
rect 9772 4088 9824 4140
rect 10692 4088 10744 4140
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 13912 4156 13964 4208
rect 17316 4156 17368 4208
rect 19708 4267 19760 4276
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13176 4088 13228 4140
rect 9956 4020 10008 4029
rect 13820 4020 13872 4072
rect 14280 4088 14332 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 20812 4088 20864 4140
rect 22468 4088 22520 4140
rect 15292 4020 15344 4072
rect 17776 4020 17828 4072
rect 18604 4020 18656 4072
rect 19432 4020 19484 4072
rect 20628 4020 20680 4072
rect 8484 3952 8536 4004
rect 2872 3884 2924 3936
rect 5448 3884 5500 3936
rect 6644 3884 6696 3936
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 9588 3884 9640 3936
rect 17868 3952 17920 4004
rect 18328 3995 18380 4004
rect 18328 3961 18362 3995
rect 18362 3961 18380 3995
rect 18328 3952 18380 3961
rect 18420 3952 18472 4004
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 10876 3927 10928 3936
rect 10876 3893 10885 3927
rect 10885 3893 10919 3927
rect 10919 3893 10928 3927
rect 10876 3884 10928 3893
rect 10968 3927 11020 3936
rect 10968 3893 10977 3927
rect 10977 3893 11011 3927
rect 11011 3893 11020 3927
rect 10968 3884 11020 3893
rect 11704 3884 11756 3936
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 14464 3927 14516 3936
rect 14464 3893 14473 3927
rect 14473 3893 14507 3927
rect 14507 3893 14516 3927
rect 14464 3884 14516 3893
rect 15108 3884 15160 3936
rect 16488 3884 16540 3936
rect 17040 3884 17092 3936
rect 17500 3884 17552 3936
rect 18972 3884 19024 3936
rect 19708 3884 19760 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3424 3680 3476 3732
rect 4160 3680 4212 3732
rect 6092 3680 6144 3732
rect 8300 3680 8352 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 9036 3680 9088 3732
rect 10876 3680 10928 3732
rect 6736 3612 6788 3664
rect 6828 3544 6880 3596
rect 7196 3544 7248 3596
rect 8208 3544 8260 3596
rect 13084 3680 13136 3732
rect 11152 3544 11204 3596
rect 11980 3544 12032 3596
rect 14372 3680 14424 3732
rect 16580 3680 16632 3732
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 17500 3723 17552 3732
rect 17500 3689 17509 3723
rect 17509 3689 17543 3723
rect 17543 3689 17552 3723
rect 17500 3680 17552 3689
rect 17868 3723 17920 3732
rect 17868 3689 17877 3723
rect 17877 3689 17911 3723
rect 17911 3689 17920 3723
rect 17868 3680 17920 3689
rect 18052 3680 18104 3732
rect 18972 3680 19024 3732
rect 14188 3612 14240 3664
rect 18420 3612 18472 3664
rect 20076 3680 20128 3732
rect 20352 3680 20404 3732
rect 20628 3680 20680 3732
rect 14280 3544 14332 3596
rect 15200 3544 15252 3596
rect 16488 3544 16540 3596
rect 10876 3476 10928 3528
rect 12992 3476 13044 3528
rect 18328 3476 18380 3528
rect 19156 3612 19208 3664
rect 20720 3612 20772 3664
rect 18880 3587 18932 3596
rect 18880 3553 18889 3587
rect 18889 3553 18923 3587
rect 18923 3553 18932 3587
rect 18880 3544 18932 3553
rect 19248 3544 19300 3596
rect 19708 3476 19760 3528
rect 2320 3340 2372 3392
rect 8944 3340 8996 3392
rect 9680 3340 9732 3392
rect 10324 3340 10376 3392
rect 19800 3408 19852 3460
rect 20536 3476 20588 3528
rect 20720 3476 20772 3528
rect 10784 3340 10836 3392
rect 11152 3340 11204 3392
rect 15936 3340 15988 3392
rect 20076 3340 20128 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 8392 3136 8444 3188
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 10692 3136 10744 3188
rect 12900 3136 12952 3188
rect 14280 3179 14332 3188
rect 14280 3145 14289 3179
rect 14289 3145 14323 3179
rect 14323 3145 14332 3179
rect 14280 3136 14332 3145
rect 15108 3179 15160 3188
rect 15108 3145 15117 3179
rect 15117 3145 15151 3179
rect 15151 3145 15160 3179
rect 15108 3136 15160 3145
rect 16580 3136 16632 3188
rect 19340 3136 19392 3188
rect 20168 3136 20220 3188
rect 8852 3068 8904 3120
rect 10876 3068 10928 3120
rect 1768 2932 1820 2984
rect 6736 2932 6788 2984
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 10600 3000 10652 3052
rect 11980 3043 12032 3052
rect 9680 2932 9732 2984
rect 10784 2932 10836 2984
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 13912 3068 13964 3120
rect 8300 2864 8352 2916
rect 11796 2907 11848 2916
rect 11796 2873 11805 2907
rect 11805 2873 11839 2907
rect 11839 2873 11848 2907
rect 11796 2864 11848 2873
rect 5632 2796 5684 2848
rect 12624 2864 12676 2916
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12992 2932 13044 2984
rect 13636 2932 13688 2984
rect 15936 3000 15988 3052
rect 14556 2975 14608 2984
rect 14556 2941 14565 2975
rect 14565 2941 14599 2975
rect 14599 2941 14608 2975
rect 14556 2932 14608 2941
rect 13728 2864 13780 2916
rect 17040 3068 17092 3120
rect 18880 3068 18932 3120
rect 16212 3000 16264 3052
rect 16488 3000 16540 3052
rect 15476 2839 15528 2848
rect 12440 2796 12492 2805
rect 15476 2805 15485 2839
rect 15485 2805 15519 2839
rect 15519 2805 15528 2839
rect 15476 2796 15528 2805
rect 17684 2932 17736 2984
rect 18512 2932 18564 2984
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 18972 3000 19024 3052
rect 19248 3000 19300 3052
rect 19800 3000 19852 3052
rect 20444 3000 20496 3052
rect 19432 2932 19484 2984
rect 19616 2932 19668 2984
rect 18880 2864 18932 2916
rect 19248 2864 19300 2916
rect 21364 2864 21416 2916
rect 16580 2839 16632 2848
rect 16580 2805 16589 2839
rect 16589 2805 16623 2839
rect 16623 2805 16632 2839
rect 16580 2796 16632 2805
rect 17500 2796 17552 2848
rect 19800 2839 19852 2848
rect 19800 2805 19809 2839
rect 19809 2805 19843 2839
rect 19843 2805 19852 2839
rect 19800 2796 19852 2805
rect 20628 2796 20680 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 8300 2592 8352 2644
rect 8852 2592 8904 2644
rect 10968 2592 11020 2644
rect 12440 2592 12492 2644
rect 15476 2592 15528 2644
rect 17592 2592 17644 2644
rect 19248 2592 19300 2644
rect 7840 2524 7892 2576
rect 10600 2567 10652 2576
rect 10600 2533 10609 2567
rect 10609 2533 10643 2567
rect 10643 2533 10652 2567
rect 10600 2524 10652 2533
rect 15384 2524 15436 2576
rect 7196 2456 7248 2508
rect 11888 2456 11940 2508
rect 14004 2456 14056 2508
rect 8208 2388 8260 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 8300 2320 8352 2372
rect 8852 2320 8904 2372
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 16212 2388 16264 2440
rect 17408 2456 17460 2508
rect 17960 2456 18012 2508
rect 18880 2456 18932 2508
rect 19064 2456 19116 2508
rect 19892 2456 19944 2508
rect 20444 2456 20496 2508
rect 17132 2388 17184 2440
rect 14464 2320 14516 2372
rect 14832 2320 14884 2372
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 12624 2252 12676 2304
rect 16488 2252 16540 2304
rect 17960 2252 18012 2304
rect 20812 2320 20864 2372
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 8300 2048 8352 2100
rect 8760 2048 8812 2100
rect 18788 2048 18840 2100
rect 19800 2048 19852 2100
rect 9956 1164 10008 1216
rect 15844 1164 15896 1216
rect 10508 824 10560 876
rect 15660 824 15712 876
rect 8300 620 8352 672
rect 11796 620 11848 672
rect 12072 552 12124 604
rect 15016 552 15068 604
<< metal2 >>
rect 5722 22320 5778 22800
rect 17130 22320 17186 22800
rect 18878 22536 18934 22545
rect 18878 22471 18934 22480
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 5736 19242 5764 22320
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 15948 18902 15976 19246
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4066 11520 4122 11529
rect 4066 11455 4122 11464
rect 664 11348 716 11354
rect 664 11290 716 11296
rect 202 3632 258 3641
rect 202 3567 258 3576
rect 216 480 244 3567
rect 676 480 704 11290
rect 4080 11286 4108 11455
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 1216 6928 1268 6934
rect 1216 6870 1268 6876
rect 1228 480 1256 6870
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 480 1808 2926
rect 2332 480 2360 3334
rect 2884 480 2912 3878
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3436 480 3464 3674
rect 3988 480 4016 4014
rect 4172 3738 4200 4422
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 1986 4752 7686
rect 4540 1958 4752 1986
rect 4540 480 4568 1958
rect 5092 480 5120 9046
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5914 6684 6054
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 7300 5710 7328 6190
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7300 5098 7328 5646
rect 7576 5370 7604 5714
rect 7668 5574 7696 18158
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 8128 5302 8156 5782
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 3942 5488 4966
rect 6288 4690 6316 5034
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 7300 4146 7328 5034
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 480 5672 2790
rect 6104 480 6132 3674
rect 6656 480 6684 3878
rect 6736 3664 6788 3670
rect 7300 3618 7328 4082
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8312 3738 8340 8026
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 6736 3606 6788 3612
rect 6748 2990 6776 3606
rect 7208 3602 7328 3618
rect 8298 3632 8354 3641
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 7196 3596 7328 3602
rect 7248 3590 7328 3596
rect 8208 3596 8260 3602
rect 7196 3538 7248 3544
rect 8298 3567 8354 3576
rect 8208 3538 8260 3544
rect 6840 3058 6868 3538
rect 8220 3194 8248 3538
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7208 480 7236 2450
rect 7852 1306 7880 2518
rect 8220 2446 8248 3130
rect 8312 3097 8340 3567
rect 8404 3194 8432 14418
rect 9600 9178 9628 14894
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 8022 8616 8366
rect 9324 8362 9352 8842
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 8090 9352 8298
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8680 5574 8708 6122
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8496 3738 8524 3946
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8298 3088 8354 3097
rect 8298 3023 8354 3032
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8312 2650 8340 2858
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8312 2106 8340 2314
rect 8772 2106 8800 5034
rect 9048 4826 9076 5170
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8956 3398 8984 4626
rect 9140 4622 9168 5510
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9232 4282 9260 7890
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9508 3942 9536 8910
rect 9692 6730 9720 18770
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 11072 13938 11100 14282
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 8974 10364 9318
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8430 10364 8910
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10336 6866 10364 8366
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9588 6248 9640 6254
rect 9640 6196 9720 6202
rect 9588 6190 9720 6196
rect 9600 6174 9720 6190
rect 9692 5574 9720 6174
rect 10060 5914 10088 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9784 4146 9812 4218
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9968 4078 9996 4626
rect 10152 4554 10180 6734
rect 10244 6254 10272 6734
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10428 5914 10456 9386
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10336 5166 10364 5510
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8864 2650 8892 3062
rect 9048 3058 9076 3674
rect 9600 3482 9628 3878
rect 9416 3454 9628 3482
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 8760 2100 8812 2106
rect 8760 2042 8812 2048
rect 7760 1278 7880 1306
rect 7760 480 7788 1278
rect 8300 672 8352 678
rect 8300 614 8352 620
rect 8312 480 8340 614
rect 8864 480 8892 2314
rect 9416 480 9444 3454
rect 10336 3398 10364 5102
rect 10520 3942 10548 13806
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10888 7546 10916 9454
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 7818 11008 8298
rect 11072 8090 11100 9318
rect 11624 9042 11652 9522
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8634 11652 8978
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10888 5846 10916 7482
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6458 11008 6802
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11072 6254 11100 7822
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11716 7546 11744 18770
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 9654 11836 15506
rect 11900 9722 11928 17682
rect 14476 17202 14504 17682
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11900 8498 11928 9386
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11060 6248 11112 6254
rect 11624 6202 11652 6598
rect 11808 6458 11836 7142
rect 11992 6610 12020 10474
rect 12452 9042 12480 11086
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12452 7954 12480 8978
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12084 7410 12112 7890
rect 12452 7750 12480 7890
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 7002 12112 7346
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12360 7002 12388 7210
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 11900 6582 12020 6610
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11060 6190 11112 6196
rect 11532 6174 11652 6202
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 5030 10824 5578
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4758 10824 4966
rect 10888 4826 10916 5646
rect 11072 5166 11100 5714
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 9692 2990 9720 3334
rect 10612 3058 10640 4558
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 3194 10732 4082
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10888 3738 10916 3878
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 10612 2582 10640 2994
rect 10796 2990 10824 3334
rect 10888 3126 10916 3470
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10796 2446 10824 2926
rect 10980 2650 11008 3878
rect 11164 3602 11192 6054
rect 11532 5778 11560 6174
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11624 5114 11652 5510
rect 11532 5098 11652 5114
rect 11520 5092 11652 5098
rect 11572 5086 11652 5092
rect 11520 5034 11572 5040
rect 11624 4622 11652 5086
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11152 3392 11204 3398
rect 11072 3352 11152 3380
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 9956 1216 10008 1222
rect 9956 1158 10008 1164
rect 9968 480 9996 1158
rect 10508 876 10560 882
rect 10508 818 10560 824
rect 10520 480 10548 818
rect 11072 480 11100 3352
rect 11152 3334 11204 3340
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11716 2990 11744 3878
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11624 480 11652 2246
rect 11808 678 11836 2858
rect 11900 2514 11928 6582
rect 12544 3942 12572 13262
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13464 11762 13492 12310
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 8838 12756 8978
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 7410 12756 8774
rect 12820 7546 12848 9998
rect 13004 9586 13032 10066
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13096 8090 13124 11154
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11992 3058 12020 3538
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12636 2922 12664 7210
rect 13096 6866 13124 8026
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13188 6730 13216 11494
rect 13464 11082 13492 11698
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13648 11354 13676 11630
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13924 10266 13952 15506
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9518 13768 9862
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 9178 13768 9454
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8430 13400 8774
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7410 13492 7890
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13924 7342 13952 8230
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13280 6934 13308 7142
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13832 5370 13860 6054
rect 13924 5370 13952 6054
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13464 4282 13492 4966
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3194 12940 3878
rect 13096 3738 13124 4082
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13004 2990 13032 3470
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2650 12480 2790
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 11796 672 11848 678
rect 11796 614 11848 620
rect 12072 604 12124 610
rect 12072 546 12124 552
rect 12084 480 12112 546
rect 12636 480 12664 2246
rect 13188 480 13216 4082
rect 13832 4078 13860 4422
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13924 3126 13952 4150
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13648 2446 13676 2926
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13740 480 13768 2858
rect 14016 2514 14044 8910
rect 14108 3942 14136 12718
rect 14200 6458 14228 17070
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15672 12986 15700 18770
rect 15764 18290 15792 18838
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15488 12442 15516 12582
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15396 11762 15424 12242
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15580 11354 15608 12582
rect 15672 11898 15700 12786
rect 16132 12374 16160 13806
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15672 11694 15700 11834
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15856 11626 15884 12038
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14384 5914 14412 6258
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14476 5778 14504 7686
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14476 5234 14504 5714
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14200 4826 14228 5034
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14292 4826 14320 4966
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14200 1986 14228 3606
rect 14292 3602 14320 4082
rect 14384 3738 14412 4558
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14292 3194 14320 3538
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14476 2378 14504 3878
rect 14568 2990 14596 8298
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14660 6458 14688 6734
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14752 5166 14780 5646
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 14200 1958 14320 1986
rect 14292 480 14320 1958
rect 14844 480 14872 2314
rect 15028 610 15056 9386
rect 15304 9178 15332 10474
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15396 9722 15424 10066
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15580 8566 15608 11154
rect 15856 11150 15884 11562
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10266 15792 10406
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 9382 15884 10066
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 8974 15884 9318
rect 15948 9178 15976 11290
rect 15936 9172 15988 9178
rect 15988 9132 16068 9160
rect 15936 9114 15988 9120
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15212 6662 15240 7754
rect 15580 7342 15608 8502
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15672 6322 15700 6802
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15764 5914 15792 6802
rect 15856 6798 15884 7210
rect 15948 7206 15976 8366
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 6322 15884 6734
rect 15948 6662 15976 7142
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 16040 6254 16068 9132
rect 16316 7562 16344 14010
rect 16408 9178 16436 16594
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16500 14414 16528 14894
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 17144 13870 17172 22320
rect 18510 21584 18566 21593
rect 18510 21519 18566 21528
rect 17774 21176 17830 21185
rect 17774 21111 17830 21120
rect 17788 19174 17816 21111
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17880 18902 17908 19246
rect 18524 19174 18552 21519
rect 18892 19310 18920 22471
rect 20074 22128 20130 22137
rect 20074 22063 20130 22072
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17328 16726 17356 17002
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17604 12986 17632 18770
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17866 18320 17922 18329
rect 17866 18255 17922 18264
rect 17880 17882 17908 18255
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16500 10826 16528 12650
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11898 16804 12242
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16500 10798 16620 10826
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16500 9926 16528 10610
rect 16592 10606 16620 10798
rect 16776 10674 16804 11834
rect 17328 11762 17356 12582
rect 17604 12374 17632 12786
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17604 11014 17632 12174
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9518 16528 9862
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16224 7546 16344 7562
rect 16212 7540 16344 7546
rect 16264 7534 16344 7540
rect 16212 7482 16264 7488
rect 16316 6322 16344 7534
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5914 16160 6054
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15212 4146 15240 4626
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15120 3194 15148 3878
rect 15212 3602 15240 4082
rect 15304 4078 15332 5238
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15488 2650 15516 2790
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 15016 604 15068 610
rect 15016 546 15068 552
rect 15396 480 15424 2518
rect 15672 882 15700 5714
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15764 5370 15792 5646
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15764 5098 15792 5306
rect 15752 5092 15804 5098
rect 15752 5034 15804 5040
rect 15856 1222 15884 5782
rect 16316 5710 16344 6258
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16500 3602 16528 3878
rect 16592 3738 16620 10406
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 8362 16804 9318
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16776 7886 16804 8298
rect 16868 8090 16896 8910
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16960 8022 16988 10406
rect 17604 10062 17632 10950
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9722 17632 9998
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17604 9518 17632 9658
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8294 17172 8910
rect 17512 8498 17540 8978
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 17144 7954 17172 8230
rect 17696 8022 17724 12718
rect 18510 12472 18566 12481
rect 18510 12407 18566 12416
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18524 11762 18552 12407
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18892 11694 18920 12038
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18432 11150 18460 11630
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10674 18000 10950
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17972 10198 18000 10610
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 18064 10010 18092 10542
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 17972 9982 18092 10010
rect 17972 9586 18000 9982
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18432 9042 18460 9454
rect 18616 9110 18644 10406
rect 18786 9752 18842 9761
rect 18786 9687 18842 9696
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18800 8480 18828 9687
rect 18892 8634 18920 11222
rect 19076 10033 19104 19246
rect 19904 18902 19932 19858
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19246 14376 19302 14385
rect 19246 14311 19302 14320
rect 19260 14074 19288 14311
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19432 13864 19484 13870
rect 19246 13832 19302 13841
rect 19432 13806 19484 13812
rect 19246 13767 19302 13776
rect 19260 13530 19288 13767
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19246 13016 19302 13025
rect 19246 12951 19248 12960
rect 19300 12951 19302 12960
rect 19248 12922 19300 12928
rect 19352 12374 19380 13330
rect 19444 12850 19472 13806
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19062 10024 19118 10033
rect 18972 9988 19024 9994
rect 19062 9959 19118 9968
rect 18972 9930 19024 9936
rect 18984 9518 19012 9930
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18616 8452 18828 8480
rect 17684 8016 17736 8022
rect 17406 7984 17462 7993
rect 17132 7948 17184 7954
rect 17684 7958 17736 7964
rect 17406 7919 17462 7928
rect 17592 7948 17644 7954
rect 17132 7890 17184 7896
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6866 16896 7142
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16776 5030 16804 5850
rect 16948 5092 17000 5098
rect 16948 5034 17000 5040
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16960 4282 16988 5034
rect 17052 4690 17080 6598
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17052 3738 17080 3878
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 3058 15976 3334
rect 16026 3088 16082 3097
rect 15936 3052 15988 3058
rect 16500 3058 16528 3538
rect 17236 3233 17264 5102
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17328 4214 17356 4626
rect 17316 4208 17368 4214
rect 17316 4150 17368 4156
rect 17222 3224 17278 3233
rect 16580 3188 16632 3194
rect 17222 3159 17278 3168
rect 16580 3130 16632 3136
rect 16026 3023 16082 3032
rect 16212 3052 16264 3058
rect 15936 2994 15988 3000
rect 16040 1578 16068 3023
rect 16212 2994 16264 3000
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16224 2446 16252 2994
rect 16592 2854 16620 3130
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 15948 1550 16068 1578
rect 15844 1216 15896 1222
rect 15844 1158 15896 1164
rect 15660 876 15712 882
rect 15660 818 15712 824
rect 15948 480 15976 1550
rect 16500 480 16528 2246
rect 17052 480 17080 3062
rect 17130 2816 17186 2825
rect 17130 2751 17186 2760
rect 17144 2446 17172 2751
rect 17420 2514 17448 7919
rect 17592 7890 17644 7896
rect 17604 7274 17632 7890
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18510 7440 18566 7449
rect 18510 7375 18566 7384
rect 17592 7268 17644 7274
rect 17592 7210 17644 7216
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17512 3738 17540 3878
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17604 2961 17632 7210
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17682 7032 17738 7041
rect 17682 6967 17738 6976
rect 17696 2990 17724 6967
rect 17972 6798 18000 7142
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17788 4486 17816 5170
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4078 17816 4422
rect 17880 4162 17908 5306
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 17972 4264 18000 4694
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17972 4236 18092 4264
rect 17880 4134 18000 4162
rect 18064 4146 18092 4236
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17972 4026 18000 4134
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17868 4004 17920 4010
rect 17972 3998 18092 4026
rect 17868 3946 17920 3952
rect 17880 3738 17908 3946
rect 17958 3768 18014 3777
rect 17868 3732 17920 3738
rect 18064 3738 18092 3998
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 17958 3703 18014 3712
rect 18052 3732 18104 3738
rect 17868 3674 17920 3680
rect 17684 2984 17736 2990
rect 17590 2952 17646 2961
rect 17684 2926 17736 2932
rect 17590 2887 17646 2896
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17512 480 17540 2790
rect 17604 2650 17632 2887
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17972 2514 18000 3703
rect 18052 3674 18104 3680
rect 18340 3534 18368 3946
rect 18432 3670 18460 3946
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18524 2990 18552 7375
rect 18616 5914 18644 8452
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18616 4826 18644 5850
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 1170 18000 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18092 1170
rect 18064 480 18092 1142
rect 18616 480 18644 4014
rect 18708 2990 18736 7686
rect 18800 6644 18828 8298
rect 18892 7886 18920 8570
rect 18984 8430 19012 8910
rect 19076 8498 19104 9862
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18880 6656 18932 6662
rect 18800 6616 18880 6644
rect 18800 6254 18828 6616
rect 18880 6598 18932 6604
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18788 5772 18840 5778
rect 18788 5714 18840 5720
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18800 2106 18828 5714
rect 18878 4720 18934 4729
rect 18878 4655 18934 4664
rect 18892 3602 18920 4655
rect 18984 3942 19012 6394
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19076 5250 19104 6122
rect 19168 5370 19196 12242
rect 19246 11656 19302 11665
rect 19246 11591 19302 11600
rect 19260 9518 19288 11591
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19352 10606 19380 11290
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 19260 8498 19288 9046
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5914 19288 6054
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19352 5302 19380 9862
rect 19444 8838 19472 12650
rect 19536 10810 19564 16594
rect 19628 11626 19656 18770
rect 19996 18698 20024 19246
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19904 16726 19932 17070
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19996 15434 20024 15982
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19890 14784 19946 14793
rect 19890 14719 19946 14728
rect 19904 14618 19932 14719
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19720 13462 19748 14418
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19708 13456 19760 13462
rect 19708 13398 19760 13404
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19706 10160 19762 10169
rect 19616 10124 19668 10130
rect 19706 10095 19708 10104
rect 19616 10066 19668 10072
rect 19760 10095 19762 10104
rect 19708 10066 19760 10072
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19628 7954 19656 10066
rect 19812 9466 19840 12718
rect 19904 12714 19932 13874
rect 20088 13870 20116 22063
rect 20626 20768 20682 20777
rect 20626 20703 20682 20712
rect 20166 20224 20222 20233
rect 20166 20159 20222 20168
rect 20180 19514 20208 20159
rect 20640 20058 20668 20703
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20166 19408 20222 19417
rect 20166 19343 20222 19352
rect 20180 18426 20208 19343
rect 20442 18864 20498 18873
rect 20442 18799 20498 18808
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20456 17882 20484 18799
rect 20732 18426 20760 19751
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20718 18048 20774 18057
rect 20718 17983 20774 17992
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20166 17504 20222 17513
rect 20166 17439 20222 17448
rect 20180 17338 20208 17439
rect 20732 17338 20760 17983
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20718 17096 20774 17105
rect 20718 17031 20774 17040
rect 20166 16552 20222 16561
rect 20166 16487 20222 16496
rect 20180 16250 20208 16487
rect 20732 16250 20760 17031
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20442 16144 20498 16153
rect 20442 16079 20498 16088
rect 20456 15706 20484 16079
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20548 15638 20576 15982
rect 20718 15736 20774 15745
rect 20718 15671 20774 15680
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20272 14890 20300 15506
rect 20442 15192 20498 15201
rect 20732 15162 20760 15671
rect 20442 15127 20498 15136
rect 20720 15156 20772 15162
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20456 14618 20484 15127
rect 20720 15098 20772 15104
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 20442 13424 20498 13433
rect 20442 13359 20498 13368
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 20272 12306 20300 12650
rect 20456 12442 20484 13359
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20626 12064 20682 12073
rect 20626 11999 20682 12008
rect 20640 11762 20668 11999
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 19996 11286 20024 11494
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19996 10674 20024 11222
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 20272 10606 20300 11494
rect 20350 10704 20406 10713
rect 20350 10639 20406 10648
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20364 10130 20392 10639
rect 20456 10470 20484 11494
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20534 11112 20590 11121
rect 20534 11047 20590 11056
rect 20548 10674 20576 11047
rect 20640 10674 20668 11154
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 10198 20484 10406
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20534 9752 20590 9761
rect 20534 9687 20590 9696
rect 19720 9438 19840 9466
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19720 6730 19748 9438
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19890 9344 19946 9353
rect 19812 9110 19840 9318
rect 19890 9279 19946 9288
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19904 8922 19932 9279
rect 19812 8894 19932 8922
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19536 5710 19564 6190
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19340 5296 19392 5302
rect 19076 5222 19288 5250
rect 19340 5238 19392 5244
rect 19064 5160 19116 5166
rect 19062 5128 19064 5137
rect 19116 5128 19118 5137
rect 19062 5063 19118 5072
rect 19062 4312 19118 4321
rect 19062 4247 19118 4256
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18984 3369 19012 3674
rect 18970 3360 19026 3369
rect 18970 3295 19026 3304
rect 18880 3120 18932 3126
rect 18878 3088 18880 3097
rect 18932 3088 18934 3097
rect 18878 3023 18934 3032
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18892 2514 18920 2858
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18984 2417 19012 2994
rect 19076 2514 19104 4247
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 18970 2408 19026 2417
rect 18970 2343 19026 2352
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 19168 480 19196 3606
rect 19260 3602 19288 5222
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 3058 19288 3538
rect 19352 3194 19380 5102
rect 19444 4078 19472 5510
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19260 2650 19288 2858
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3974 0 4030 480
rect 4526 0 4582 480
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6090 0 6146 480
rect 6642 0 6698 480
rect 7194 0 7250 480
rect 7746 0 7802 480
rect 8298 0 8354 480
rect 8850 0 8906 480
rect 9402 0 9458 480
rect 9954 0 10010 480
rect 10506 0 10562 480
rect 11058 0 11114 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12622 0 12678 480
rect 13174 0 13230 480
rect 13726 0 13782 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 17038 0 17094 480
rect 17498 0 17554 480
rect 18050 0 18106 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19352 241 19380 3130
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 1057 19472 2926
rect 19536 2530 19564 4966
rect 19628 2990 19656 4966
rect 19720 4282 19748 5034
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19812 3890 19840 8894
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20456 8430 20484 8774
rect 20444 8424 20496 8430
rect 20350 8392 20406 8401
rect 20444 8366 20496 8372
rect 20350 8327 20406 8336
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19904 5234 19932 7890
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20088 7002 20116 7142
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 20088 6905 20116 6938
rect 20074 6896 20130 6905
rect 19984 6860 20036 6866
rect 20074 6831 20130 6840
rect 19984 6802 20036 6808
rect 19996 5642 20024 6802
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20088 6458 20116 6734
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20180 6202 20208 6734
rect 20272 6633 20300 7822
rect 20364 7562 20392 8327
rect 20456 7886 20484 8366
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20364 7534 20484 7562
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20364 6934 20392 7346
rect 20352 6928 20404 6934
rect 20352 6870 20404 6876
rect 20258 6624 20314 6633
rect 20258 6559 20314 6568
rect 20088 6174 20208 6202
rect 20088 6118 20116 6174
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20258 6080 20314 6089
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 20088 4758 20116 6054
rect 20180 5370 20208 6054
rect 20258 6015 20314 6024
rect 20272 5778 20300 6015
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20076 3936 20128 3942
rect 19720 3534 19748 3878
rect 19812 3862 19932 3890
rect 20076 3878 20128 3884
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19812 3058 19840 3402
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19536 2502 19748 2530
rect 19430 1048 19486 1057
rect 19430 983 19486 992
rect 19720 480 19748 2502
rect 19812 2106 19840 2790
rect 19904 2514 19932 3862
rect 20088 3738 20116 3878
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 20088 2666 20116 3334
rect 20180 3194 20208 3878
rect 20272 3482 20300 5578
rect 20364 5234 20392 6870
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20364 3738 20392 4762
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20272 3454 20392 3482
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20364 2904 20392 3454
rect 20456 3058 20484 7534
rect 20548 4570 20576 9687
rect 20626 8800 20682 8809
rect 20626 8735 20682 8744
rect 20640 5778 20668 8735
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20732 6254 20760 7414
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20626 5672 20682 5681
rect 20626 5607 20682 5616
rect 20640 5166 20668 5607
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20548 4542 20668 4570
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 3534 20576 4422
rect 20640 4078 20668 4542
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20364 2876 20484 2904
rect 20088 2638 20300 2666
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 19812 649 19840 2042
rect 19798 640 19854 649
rect 19798 575 19854 584
rect 20272 480 20300 2638
rect 20456 2514 20484 2876
rect 20640 2854 20668 3674
rect 20732 3670 20760 4966
rect 20824 4146 20852 19110
rect 21916 11620 21968 11626
rect 21916 11562 21968 11568
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20916 6322 20944 6598
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 20732 1601 20760 3470
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20812 2372 20864 2378
rect 20812 2314 20864 2320
rect 20718 1592 20774 1601
rect 20718 1527 20774 1536
rect 20824 480 20852 2314
rect 21376 480 21404 2858
rect 21928 480 21956 11562
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22480 480 22508 4082
rect 19338 232 19394 241
rect 19338 167 19394 176
rect 19706 0 19762 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
<< via2 >>
rect 18878 22480 18934 22536
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 11464 4122 11520
rect 202 3576 258 3632
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 8298 3576 8354 3632
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8298 3032 8354 3088
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 18510 21528 18566 21584
rect 17774 21120 17830 21176
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 20074 22072 20130 22128
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 17866 18264 17922 18320
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18510 12416 18566 12472
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18786 9696 18842 9752
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 19246 14320 19302 14376
rect 19246 13776 19302 13832
rect 19246 12980 19302 13016
rect 19246 12960 19248 12980
rect 19248 12960 19300 12980
rect 19300 12960 19302 12980
rect 19062 9968 19118 10024
rect 17406 7928 17462 7984
rect 16026 3032 16082 3088
rect 17222 3168 17278 3224
rect 17130 2760 17186 2816
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18510 7384 18566 7440
rect 17682 6976 17738 7032
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17958 3712 18014 3768
rect 17590 2896 17646 2952
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18878 4664 18934 4720
rect 19246 11600 19302 11656
rect 19890 14728 19946 14784
rect 19706 10124 19762 10160
rect 19706 10104 19708 10124
rect 19708 10104 19760 10124
rect 19760 10104 19762 10124
rect 20626 20712 20682 20768
rect 20166 20168 20222 20224
rect 20718 19760 20774 19816
rect 20166 19352 20222 19408
rect 20442 18808 20498 18864
rect 20718 17992 20774 18048
rect 20166 17448 20222 17504
rect 20718 17040 20774 17096
rect 20166 16496 20222 16552
rect 20442 16088 20498 16144
rect 20718 15680 20774 15736
rect 20442 15136 20498 15192
rect 20442 13368 20498 13424
rect 20626 12008 20682 12064
rect 20350 10648 20406 10704
rect 20534 11056 20590 11112
rect 20534 9696 20590 9752
rect 19890 9288 19946 9344
rect 19062 5108 19064 5128
rect 19064 5108 19116 5128
rect 19116 5108 19118 5128
rect 19062 5072 19118 5108
rect 19062 4256 19118 4312
rect 18970 3304 19026 3360
rect 18878 3068 18880 3088
rect 18880 3068 18932 3088
rect 18932 3068 18934 3088
rect 18878 3032 18934 3068
rect 18970 2352 19026 2408
rect 20350 8336 20406 8392
rect 20074 6840 20130 6896
rect 20258 6568 20314 6624
rect 20258 6024 20314 6080
rect 19430 992 19486 1048
rect 20626 8744 20682 8800
rect 20626 5616 20682 5672
rect 19798 584 19854 640
rect 20718 1536 20774 1592
rect 19338 176 19394 232
<< metal3 >>
rect 18873 22538 18939 22541
rect 22320 22538 22800 22568
rect 18873 22536 22800 22538
rect 18873 22480 18878 22536
rect 18934 22480 22800 22536
rect 18873 22478 22800 22480
rect 18873 22475 18939 22478
rect 22320 22448 22800 22478
rect 20069 22130 20135 22133
rect 22320 22130 22800 22160
rect 20069 22128 22800 22130
rect 20069 22072 20074 22128
rect 20130 22072 22800 22128
rect 20069 22070 22800 22072
rect 20069 22067 20135 22070
rect 22320 22040 22800 22070
rect 18505 21586 18571 21589
rect 22320 21586 22800 21616
rect 18505 21584 22800 21586
rect 18505 21528 18510 21584
rect 18566 21528 22800 21584
rect 18505 21526 22800 21528
rect 18505 21523 18571 21526
rect 22320 21496 22800 21526
rect 17769 21178 17835 21181
rect 22320 21178 22800 21208
rect 17769 21176 22800 21178
rect 17769 21120 17774 21176
rect 17830 21120 22800 21176
rect 17769 21118 22800 21120
rect 17769 21115 17835 21118
rect 22320 21088 22800 21118
rect 20621 20770 20687 20773
rect 22320 20770 22800 20800
rect 20621 20768 22800 20770
rect 20621 20712 20626 20768
rect 20682 20712 22800 20768
rect 20621 20710 22800 20712
rect 20621 20707 20687 20710
rect 22320 20680 22800 20710
rect 20161 20226 20227 20229
rect 22320 20226 22800 20256
rect 20161 20224 22800 20226
rect 20161 20168 20166 20224
rect 20222 20168 22800 20224
rect 20161 20166 22800 20168
rect 20161 20163 20227 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 20713 19818 20779 19821
rect 22320 19818 22800 19848
rect 20713 19816 22800 19818
rect 20713 19760 20718 19816
rect 20774 19760 22800 19816
rect 20713 19758 22800 19760
rect 20713 19755 20779 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 20161 19410 20227 19413
rect 22320 19410 22800 19440
rect 20161 19408 22800 19410
rect 20161 19352 20166 19408
rect 20222 19352 22800 19408
rect 20161 19350 22800 19352
rect 20161 19347 20227 19350
rect 22320 19320 22800 19350
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 20437 18866 20503 18869
rect 22320 18866 22800 18896
rect 20437 18864 22800 18866
rect 20437 18808 20442 18864
rect 20498 18808 22800 18864
rect 20437 18806 22800 18808
rect 20437 18803 20503 18806
rect 22320 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 22320 18458 22800 18488
rect 18646 18398 22800 18458
rect 17861 18322 17927 18325
rect 18646 18322 18706 18398
rect 22320 18368 22800 18398
rect 17861 18320 18706 18322
rect 17861 18264 17866 18320
rect 17922 18264 18706 18320
rect 17861 18262 18706 18264
rect 17861 18259 17927 18262
rect 20713 18050 20779 18053
rect 22320 18050 22800 18080
rect 20713 18048 22800 18050
rect 20713 17992 20718 18048
rect 20774 17992 22800 18048
rect 20713 17990 22800 17992
rect 20713 17987 20779 17990
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 22320 17960 22800 17990
rect 14672 17919 14992 17920
rect 20161 17506 20227 17509
rect 22320 17506 22800 17536
rect 20161 17504 22800 17506
rect 20161 17448 20166 17504
rect 20222 17448 22800 17504
rect 20161 17446 22800 17448
rect 20161 17443 20227 17446
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 22320 17416 22800 17446
rect 18104 17375 18424 17376
rect 20713 17098 20779 17101
rect 22320 17098 22800 17128
rect 20713 17096 22800 17098
rect 20713 17040 20718 17096
rect 20774 17040 22800 17096
rect 20713 17038 22800 17040
rect 20713 17035 20779 17038
rect 22320 17008 22800 17038
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 20161 16554 20227 16557
rect 22320 16554 22800 16584
rect 20161 16552 22800 16554
rect 20161 16496 20166 16552
rect 20222 16496 22800 16552
rect 20161 16494 22800 16496
rect 20161 16491 20227 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 20437 16146 20503 16149
rect 22320 16146 22800 16176
rect 20437 16144 22800 16146
rect 20437 16088 20442 16144
rect 20498 16088 22800 16144
rect 20437 16086 22800 16088
rect 20437 16083 20503 16086
rect 22320 16056 22800 16086
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 20713 15738 20779 15741
rect 22320 15738 22800 15768
rect 20713 15736 22800 15738
rect 20713 15680 20718 15736
rect 20774 15680 22800 15736
rect 20713 15678 22800 15680
rect 20713 15675 20779 15678
rect 22320 15648 22800 15678
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 20437 15194 20503 15197
rect 22320 15194 22800 15224
rect 20437 15192 22800 15194
rect 20437 15136 20442 15192
rect 20498 15136 22800 15192
rect 20437 15134 22800 15136
rect 20437 15131 20503 15134
rect 22320 15104 22800 15134
rect 19885 14786 19951 14789
rect 22320 14786 22800 14816
rect 19885 14784 22800 14786
rect 19885 14728 19890 14784
rect 19946 14728 22800 14784
rect 19885 14726 22800 14728
rect 19885 14723 19951 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 22320 14696 22800 14726
rect 14672 14655 14992 14656
rect 19241 14378 19307 14381
rect 22320 14378 22800 14408
rect 19241 14376 22800 14378
rect 19241 14320 19246 14376
rect 19302 14320 22800 14376
rect 19241 14318 22800 14320
rect 19241 14315 19307 14318
rect 22320 14288 22800 14318
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 19241 13834 19307 13837
rect 22320 13834 22800 13864
rect 19241 13832 22800 13834
rect 19241 13776 19246 13832
rect 19302 13776 22800 13832
rect 19241 13774 22800 13776
rect 19241 13771 19307 13774
rect 22320 13744 22800 13774
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 20437 13426 20503 13429
rect 22320 13426 22800 13456
rect 20437 13424 22800 13426
rect 20437 13368 20442 13424
rect 20498 13368 22800 13424
rect 20437 13366 22800 13368
rect 20437 13363 20503 13366
rect 22320 13336 22800 13366
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 19241 13018 19307 13021
rect 22320 13018 22800 13048
rect 19241 13016 22800 13018
rect 19241 12960 19246 13016
rect 19302 12960 22800 13016
rect 19241 12958 22800 12960
rect 19241 12955 19307 12958
rect 22320 12928 22800 12958
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 18505 12474 18571 12477
rect 22320 12474 22800 12504
rect 18505 12472 22800 12474
rect 18505 12416 18510 12472
rect 18566 12416 22800 12472
rect 18505 12414 22800 12416
rect 18505 12411 18571 12414
rect 22320 12384 22800 12414
rect 20621 12066 20687 12069
rect 22320 12066 22800 12096
rect 20621 12064 22800 12066
rect 20621 12008 20626 12064
rect 20682 12008 22800 12064
rect 20621 12006 22800 12008
rect 20621 12003 20687 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 22320 11976 22800 12006
rect 18104 11935 18424 11936
rect 19241 11658 19307 11661
rect 22320 11658 22800 11688
rect 19241 11656 22800 11658
rect 19241 11600 19246 11656
rect 19302 11600 22800 11656
rect 19241 11598 22800 11600
rect 19241 11595 19307 11598
rect 22320 11568 22800 11598
rect 0 11522 480 11552
rect 4061 11522 4127 11525
rect 0 11520 4127 11522
rect 0 11464 4066 11520
rect 4122 11464 4127 11520
rect 0 11462 4127 11464
rect 0 11432 480 11462
rect 4061 11459 4127 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 20529 11114 20595 11117
rect 22320 11114 22800 11144
rect 20529 11112 22800 11114
rect 20529 11056 20534 11112
rect 20590 11056 22800 11112
rect 20529 11054 22800 11056
rect 20529 11051 20595 11054
rect 22320 11024 22800 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 20345 10706 20411 10709
rect 22320 10706 22800 10736
rect 20345 10704 22800 10706
rect 20345 10648 20350 10704
rect 20406 10648 22800 10704
rect 20345 10646 22800 10648
rect 20345 10643 20411 10646
rect 22320 10616 22800 10646
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 19701 10162 19767 10165
rect 22320 10162 22800 10192
rect 19701 10160 22800 10162
rect 19701 10104 19706 10160
rect 19762 10104 22800 10160
rect 19701 10102 22800 10104
rect 19701 10099 19767 10102
rect 22320 10072 22800 10102
rect 19057 10026 19123 10029
rect 18646 10024 19123 10026
rect 18646 9968 19062 10024
rect 19118 9968 19123 10024
rect 18646 9966 19123 9968
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 18646 9754 18706 9966
rect 19057 9963 19123 9966
rect 18781 9754 18847 9757
rect 18646 9752 18847 9754
rect 18646 9696 18786 9752
rect 18842 9696 18847 9752
rect 18646 9694 18847 9696
rect 18781 9691 18847 9694
rect 20529 9754 20595 9757
rect 22320 9754 22800 9784
rect 20529 9752 22800 9754
rect 20529 9696 20534 9752
rect 20590 9696 22800 9752
rect 20529 9694 22800 9696
rect 20529 9691 20595 9694
rect 22320 9664 22800 9694
rect 19885 9346 19951 9349
rect 22320 9346 22800 9376
rect 19885 9344 22800 9346
rect 19885 9288 19890 9344
rect 19946 9288 22800 9344
rect 19885 9286 22800 9288
rect 19885 9283 19951 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 22320 9256 22800 9286
rect 14672 9215 14992 9216
rect 20621 8802 20687 8805
rect 22320 8802 22800 8832
rect 20621 8800 22800 8802
rect 20621 8744 20626 8800
rect 20682 8744 22800 8800
rect 20621 8742 22800 8744
rect 20621 8739 20687 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 22320 8712 22800 8742
rect 18104 8671 18424 8672
rect 20345 8394 20411 8397
rect 22320 8394 22800 8424
rect 20345 8392 22800 8394
rect 20345 8336 20350 8392
rect 20406 8336 22800 8392
rect 20345 8334 22800 8336
rect 20345 8331 20411 8334
rect 22320 8304 22800 8334
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 17401 7986 17467 7989
rect 22320 7986 22800 8016
rect 17401 7984 22800 7986
rect 17401 7928 17406 7984
rect 17462 7928 22800 7984
rect 17401 7926 22800 7928
rect 17401 7923 17467 7926
rect 22320 7896 22800 7926
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 18505 7442 18571 7445
rect 22320 7442 22800 7472
rect 18505 7440 22800 7442
rect 18505 7384 18510 7440
rect 18566 7384 22800 7440
rect 18505 7382 22800 7384
rect 18505 7379 18571 7382
rect 22320 7352 22800 7382
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 17677 7034 17743 7037
rect 22320 7034 22800 7064
rect 17677 7032 22800 7034
rect 17677 6976 17682 7032
rect 17738 6976 22800 7032
rect 17677 6974 22800 6976
rect 17677 6971 17743 6974
rect 22320 6944 22800 6974
rect 20069 6900 20135 6901
rect 20069 6898 20116 6900
rect 20024 6896 20116 6898
rect 20024 6840 20074 6896
rect 20024 6838 20116 6840
rect 20069 6836 20116 6838
rect 20180 6836 20186 6900
rect 20069 6835 20135 6836
rect 20253 6626 20319 6629
rect 22320 6626 22800 6656
rect 20253 6624 22800 6626
rect 20253 6568 20258 6624
rect 20314 6568 22800 6624
rect 20253 6566 22800 6568
rect 20253 6563 20319 6566
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 22320 6536 22800 6566
rect 18104 6495 18424 6496
rect 20253 6082 20319 6085
rect 22320 6082 22800 6112
rect 20253 6080 22800 6082
rect 20253 6024 20258 6080
rect 20314 6024 22800 6080
rect 20253 6022 22800 6024
rect 20253 6019 20319 6022
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 22320 5992 22800 6022
rect 14672 5951 14992 5952
rect 20621 5674 20687 5677
rect 22320 5674 22800 5704
rect 20621 5672 22800 5674
rect 20621 5616 20626 5672
rect 20682 5616 22800 5672
rect 20621 5614 22800 5616
rect 20621 5611 20687 5614
rect 22320 5584 22800 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 19057 5130 19123 5133
rect 22320 5130 22800 5160
rect 19057 5128 22800 5130
rect 19057 5072 19062 5128
rect 19118 5072 22800 5128
rect 19057 5070 22800 5072
rect 19057 5067 19123 5070
rect 22320 5040 22800 5070
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 18873 4722 18939 4725
rect 22320 4722 22800 4752
rect 18873 4720 22800 4722
rect 18873 4664 18878 4720
rect 18934 4664 22800 4720
rect 18873 4662 22800 4664
rect 18873 4659 18939 4662
rect 22320 4632 22800 4662
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 19057 4314 19123 4317
rect 22320 4314 22800 4344
rect 19057 4312 22800 4314
rect 19057 4256 19062 4312
rect 19118 4256 22800 4312
rect 19057 4254 22800 4256
rect 19057 4251 19123 4254
rect 22320 4224 22800 4254
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 17953 3770 18019 3773
rect 22320 3770 22800 3800
rect 17953 3768 22800 3770
rect 17953 3712 17958 3768
rect 18014 3712 22800 3768
rect 17953 3710 22800 3712
rect 17953 3707 18019 3710
rect 22320 3680 22800 3710
rect 197 3634 263 3637
rect 8293 3634 8359 3637
rect 197 3632 2698 3634
rect 197 3576 202 3632
rect 258 3600 2698 3632
rect 2822 3632 8359 3634
rect 2822 3600 8298 3632
rect 258 3576 8298 3600
rect 8354 3576 8359 3632
rect 197 3574 8359 3576
rect 197 3571 263 3574
rect 2638 3540 2882 3574
rect 8293 3571 8359 3574
rect 18965 3362 19031 3365
rect 22320 3362 22800 3392
rect 18965 3360 19442 3362
rect 18965 3304 18970 3360
rect 19026 3304 19442 3360
rect 18965 3302 19442 3304
rect 18965 3299 19031 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 17217 3226 17283 3229
rect 11654 3224 17283 3226
rect 11654 3168 17222 3224
rect 17278 3168 17283 3224
rect 11654 3166 17283 3168
rect 19382 3226 19442 3302
rect 19566 3302 22800 3362
rect 19566 3226 19626 3302
rect 22320 3272 22800 3302
rect 19382 3166 19626 3226
rect 8293 3090 8359 3093
rect 11654 3090 11714 3166
rect 17217 3163 17283 3166
rect 8293 3088 11714 3090
rect 8293 3032 8298 3088
rect 8354 3032 11714 3088
rect 8293 3030 11714 3032
rect 16021 3090 16087 3093
rect 18873 3090 18939 3093
rect 16021 3088 18939 3090
rect 16021 3032 16026 3088
rect 16082 3032 18878 3088
rect 18934 3032 18939 3088
rect 16021 3030 18939 3032
rect 8293 3027 8359 3030
rect 16021 3027 16087 3030
rect 18873 3027 18939 3030
rect 17585 2954 17651 2957
rect 22320 2954 22800 2984
rect 17585 2952 22800 2954
rect 17585 2896 17590 2952
rect 17646 2896 22800 2952
rect 17585 2894 22800 2896
rect 17585 2891 17651 2894
rect 22320 2864 22800 2894
rect 17125 2818 17191 2821
rect 20110 2818 20116 2820
rect 17125 2816 20116 2818
rect 17125 2760 17130 2816
rect 17186 2760 20116 2816
rect 17125 2758 20116 2760
rect 17125 2755 17191 2758
rect 20110 2756 20116 2758
rect 20180 2756 20186 2820
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 18965 2410 19031 2413
rect 22320 2410 22800 2440
rect 18965 2408 22800 2410
rect 18965 2352 18970 2408
rect 19026 2352 22800 2408
rect 18965 2350 22800 2352
rect 18965 2347 19031 2350
rect 22320 2320 22800 2350
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 20110 1940 20116 2004
rect 20180 2002 20186 2004
rect 22320 2002 22800 2032
rect 20180 1942 22800 2002
rect 20180 1940 20186 1942
rect 22320 1912 22800 1942
rect 20713 1594 20779 1597
rect 22320 1594 22800 1624
rect 20713 1592 22800 1594
rect 20713 1536 20718 1592
rect 20774 1536 22800 1592
rect 20713 1534 22800 1536
rect 20713 1531 20779 1534
rect 22320 1504 22800 1534
rect 19425 1050 19491 1053
rect 22320 1050 22800 1080
rect 19425 1048 22800 1050
rect 19425 992 19430 1048
rect 19486 992 22800 1048
rect 19425 990 22800 992
rect 19425 987 19491 990
rect 22320 960 22800 990
rect 19793 642 19859 645
rect 22320 642 22800 672
rect 19793 640 22800 642
rect 19793 584 19798 640
rect 19854 584 22800 640
rect 19793 582 22800 584
rect 19793 579 19859 582
rect 22320 552 22800 582
rect 19333 234 19399 237
rect 22320 234 22800 264
rect 19333 232 22800 234
rect 19333 176 19338 232
rect 19394 176 22800 232
rect 19333 174 22800 176
rect 19333 171 19399 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 20116 6896 20180 6900
rect 20116 6840 20130 6896
rect 20130 6840 20180 6896
rect 20116 6836 20180 6840
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 20116 2756 20180 2820
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 20116 1940 20180 2004
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 20115 6900 20181 6901
rect 20115 6836 20116 6900
rect 20180 6836 20181 6900
rect 20115 6835 20181 6836
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 20118 2821 20178 6835
rect 20115 2820 20181 2821
rect 20115 2756 20116 2820
rect 20180 2756 20181 2820
rect 20115 2755 20181 2756
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 20118 2005 20178 2755
rect 20115 2004 20181 2005
rect 20115 1940 20116 2004
rect 20180 1940 20181 2004
rect 20115 1939 20181 1940
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606821651
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606821651
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7360 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1606821651
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82
timestamp 1606821651
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1606821651
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9568 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10120 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1606821651
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_89
timestamp 1606821651
transform 1 0 9292 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp 1606821651
transform 1 0 11040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1606821651
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1606821651
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11316 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _88_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606821651
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1606821651
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606821651
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12880 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12972 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_0_138
timestamp 1606821651
transform 1 0 13800 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 1606821651
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1606821651
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1606821651
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1606821651
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1606821651
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15088 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606821651
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1606821651
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15824 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16100 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1606821651
transform 1 0 16652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_176
timestamp 1606821651
transform 1 0 17296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1606821651
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1606821651
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606821651
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606821651
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606821651
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606821651
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1606821651
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_188
timestamp 1606821651
transform 1 0 18400 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_192
timestamp 1606821651
transform 1 0 18768 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 18676 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606821651
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1606821651
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_198
timestamp 1606821651
transform 1 0 19320 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19412 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606821651
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp 1606821651
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1606821651
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606821651
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606821651
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606821651
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606821651
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1606821651
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606821651
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_56
timestamp 1606821651
transform 1 0 6256 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7084 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1606821651
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_81
timestamp 1606821651
transform 1 0 8556 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1606821651
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1606821651
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11316 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_109
timestamp 1606821651
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13248 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_127
timestamp 1606821651
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_131
timestamp 1606821651
transform 1 0 13156 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1606821651
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1606821651
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606821651
transform 1 0 17020 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 17480 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_170
timestamp 1606821651
transform 1 0 16744 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1606821651
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_187
timestamp 1606821651
transform 1 0 18308 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 18860 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19412 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1606821651
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_208
timestamp 1606821651
transform 1 0 20240 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606821651
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606821651
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606821651
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606821651
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_70
timestamp 1606821651
transform 1 0 7544 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9476 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1606821651
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1606821651
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1606821651
transform 1 0 11776 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_111
timestamp 1606821651
transform 1 0 11316 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_115
timestamp 1606821651
transform 1 0 11684 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606821651
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14076 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_133
timestamp 1606821651
transform 1 0 13340 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15180 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_150
timestamp 1606821651
transform 1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16928 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1606821651
transform 1 0 16652 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606821651
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1606821651
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606821651
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1606821651
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1606821651
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606821651
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6256 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606821651
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_72
timestamp 1606821651
transform 1 0 7728 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_80
timestamp 1606821651
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1606821651
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1606821651
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_112
timestamp 1606821651
transform 1 0 11408 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_124
timestamp 1606821651
transform 1 0 12512 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13800 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_136
timestamp 1606821651
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_147
timestamp 1606821651
transform 1 0 14628 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_166
timestamp 1606821651
transform 1 0 16376 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 17020 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_172
timestamp 1606821651
transform 1 0 16928 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1606821651
transform 1 0 18492 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1606821651
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606821651
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606821651
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606821651
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1606821651
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10212 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_89
timestamp 1606821651
transform 1 0 9292 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1606821651
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606821651
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1606821651
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606821651
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_123
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12972 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1606821651
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1606821651
transform 1 0 14812 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_161
timestamp 1606821651
transform 1 0 15916 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_173
timestamp 1606821651
transform 1 0 17020 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606821651
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 19044 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1606821651
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1606821651
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 20608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1606821651
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1606821651
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606821651
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606821651
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606821651
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606821651
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6256 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606821651
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606821651
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606821651
transform 1 0 7360 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7268 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7820 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1606821651
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_83
timestamp 1606821651
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1606821651
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9476 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10396 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10120 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1606821651
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_96
timestamp 1606821651
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_89
timestamp 1606821651
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11408 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1606821651
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1606821651
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606821651
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13064 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13432 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1606821651
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_131
timestamp 1606821651
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_143
timestamp 1606821651
transform 1 0 14260 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_152
timestamp 1606821651
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606821651
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1606821651
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15272 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1606821651
transform 1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606821651
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_163
timestamp 1606821651
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1606821651
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16284 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16284 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1606821651
transform 1 0 18216 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_174
timestamp 1606821651
transform 1 0 17112 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_186
timestamp 1606821651
transform 1 0 18216 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_174
timestamp 1606821651
transform 1 0 17112 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1606821651
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606821651
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 18676 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18860 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_192
timestamp 1606821651
transform 1 0 18768 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_202
timestamp 1606821651
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_189
timestamp 1606821651
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_207
timestamp 1606821651
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 20332 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606821651
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_218
timestamp 1606821651
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606821651
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606821651
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606821651
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606821651
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1606821651
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10672 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1606821651
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606821651
transform 1 0 12328 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1606821651
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1606821651
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_136
timestamp 1606821651
transform 1 0 13616 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16284 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606821651
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606821651
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17940 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1606821651
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 19596 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1606821651
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1606821651
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606821651
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606821651
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1606821651
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1606821651
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1606821651
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606821651
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1606821651
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1606821651
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_98
timestamp 1606821651
transform 1 0 10120 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1606821651
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606821651
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13800 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12788 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1606821651
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15456 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1606821651
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 17112 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1606821651
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1606821651
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_196
timestamp 1606821651
transform 1 0 19136 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_200
timestamp 1606821651
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_210
timestamp 1606821651
transform 1 0 20424 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_218
timestamp 1606821651
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606821651
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606821651
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606821651
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606821651
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_68
timestamp 1606821651
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10580 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606821651
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1606821651
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11776 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1606821651
transform 1 0 11408 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13432 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1606821651
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16192 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1606821651
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_162
timestamp 1606821651
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17204 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1606821651
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_181
timestamp 1606821651
transform 1 0 17756 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19780 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18768 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp 1606821651
transform 1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_201
timestamp 1606821651
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1606821651
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1606821651
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606821651
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606821651
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606821651
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1606821651
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8556 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_74
timestamp 1606821651
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_80
timestamp 1606821651
transform 1 0 8464 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10212 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1606821651
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1606821651
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1606821651
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_123
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12972 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15824 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14812 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1606821651
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606821651
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1606821651
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1606821651
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 19688 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18584 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_199
timestamp 1606821651
transform 1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_218
timestamp 1606821651
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606821651
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606821651
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606821651
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606821651
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606821651
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_80
timestamp 1606821651
transform 1 0 8464 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1606821651
transform 1 0 9108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_86
timestamp 1606821651
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10764 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1606821651
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13892 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1606821651
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16376 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_163
timestamp 1606821651
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_175
timestamp 1606821651
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_187
timestamp 1606821651
transform 1 0 18308 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1606821651
transform 1 0 18584 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19044 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1606821651
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1606821651
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606821651
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606821651
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606821651
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1606821651
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1606821651
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606821651
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606821651
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1606821651
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1606821651
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1606821651
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1606821651
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1606821651
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1606821651
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_98
timestamp 1606821651
transform 1 0 10120 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_104
timestamp 1606821651
transform 1 0 10672 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11040 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 10764 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1606821651
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1606821651
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1606821651
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1606821651
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1606821651
transform 1 0 12972 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13432 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1606821651
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_129
timestamp 1606821651
transform 1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1606821651
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15364 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1606821651
transform 1 0 14904 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_154
timestamp 1606821651
transform 1 0 15272 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_175
timestamp 1606821651
transform 1 0 17204 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1606821651
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_177
timestamp 1606821651
transform 1 0 17388 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_171
timestamp 1606821651
transform 1 0 16836 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1606821651
transform 1 0 16928 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606821651
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1606821651
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17572 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606821651
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18400 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_204
timestamp 1606821651
transform 1 0 19872 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_195
timestamp 1606821651
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1606821651
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1606821651
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_210
timestamp 1606821651
transform 1 0 20424 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1606821651
transform 1 0 20516 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606821651
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606821651
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606821651
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606821651
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1606821651
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1606821651
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1606821651
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606821651
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1606821651
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1606821651
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1606821651
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1606821651
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1606821651
transform 1 0 12972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_141
timestamp 1606821651
transform 1 0 14076 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1606821651
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_164
timestamp 1606821651
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16468 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_176
timestamp 1606821651
transform 1 0 17296 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1606821651
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19044 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 20056 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1606821651
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_204
timestamp 1606821651
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1606821651
transform 1 0 20884 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1606821651
transform 1 0 21252 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606821651
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1606821651
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1606821651
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1606821651
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1606821651
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1606821651
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_117
timestamp 1606821651
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606821651
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_139
timestamp 1606821651
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1606821651
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606821651
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16836 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1606821651
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1606821651
transform 1 0 18308 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1606821651
transform 1 0 18676 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19136 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1606821651
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1606821651
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606821651
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606821651
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606821651
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606821651
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606821651
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1606821651
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1606821651
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1606821651
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1606821651
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13708 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12696 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1606821651
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15364 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_153
timestamp 1606821651
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606821651
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_171
timestamp 1606821651
transform 1 0 16836 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_177
timestamp 1606821651
transform 1 0 17388 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606821651
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18584 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 20240 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1606821651
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1606821651
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1606821651
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606821651
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1606821651
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1606821651
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1606821651
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1606821651
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1606821651
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1606821651
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_129
timestamp 1606821651
transform 1 0 12972 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606821651
transform 1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15916 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1606821651
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1606821651
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_158
timestamp 1606821651
transform 1 0 15640 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17572 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1606821651
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19412 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_195
timestamp 1606821651
transform 1 0 19044 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_205
timestamp 1606821651
transform 1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606821651
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606821651
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606821651
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606821651
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606821651
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606821651
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606821651
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606821651
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606821651
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1606821651
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1606821651
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1606821651
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1606821651
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1606821651
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1606821651
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1606821651
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1606821651
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1606821651
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1606821651
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1606821651
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1606821651
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1606821651
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15088 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1606821651
transform 1 0 14628 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_151
timestamp 1606821651
transform 1 0 14996 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_161
timestamp 1606821651
transform 1 0 15916 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1606821651
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1606821651
transform 1 0 16652 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606821651
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606821651
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_194
timestamp 1606821651
transform 1 0 18952 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_190
timestamp 1606821651
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_192
timestamp 1606821651
transform 1 0 18768 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1606821651
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1606821651
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19596 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19596 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606821651
transform 1 0 19044 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 19044 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1606821651
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1606821651
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20332 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1606821651
transform 1 0 20884 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1606821651
transform 1 0 21252 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1606821651
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606821651
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1606821651
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1606821651
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606821651
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606821651
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1606821651
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1606821651
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_98
timestamp 1606821651
transform 1 0 10120 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_104
timestamp 1606821651
transform 1 0 10672 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10764 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_111
timestamp 1606821651
transform 1 0 11316 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1606821651
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1606821651
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16100 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1606821651
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1606821651
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1606821651
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 19228 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_196
timestamp 1606821651
transform 1 0 19136 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_201
timestamp 1606821651
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1606821651
transform 1 0 20884 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_219
timestamp 1606821651
transform 1 0 21252 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606821651
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606821651
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1606821651
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_68
timestamp 1606821651
transform 1 0 7360 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_76
timestamp 1606821651
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1606821651
transform 1 0 8924 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1606821651
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1606821651
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1606821651
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1606821651
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1606821651
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1606821651
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1606821651
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606821651
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606821651
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1606821651
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1606821651
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1606821651
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606821651
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606821651
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1606821651
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1606821651
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1606821651
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606821651
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1606821651
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9568 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_86
timestamp 1606821651
transform 1 0 9016 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1606821651
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1606821651
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1606821651
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1606821651
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1606821651
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1606821651
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1606821651
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_208
timestamp 1606821651
transform 1 0 20240 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606821651
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606821651
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606821651
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1606821651
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606821651
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1606821651
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1606821651
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1606821651
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1606821651
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11776 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_105
timestamp 1606821651
transform 1 0 10764 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_113
timestamp 1606821651
transform 1 0 11500 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_122
timestamp 1606821651
transform 1 0 12328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13892 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_134
timestamp 1606821651
transform 1 0 13432 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_138
timestamp 1606821651
transform 1 0 13800 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1606821651
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606821651
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606821651
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606821651
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606821651
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_202
timestamp 1606821651
transform 1 0 19688 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606821651
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1606821651
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1606821651
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1606821651
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1606821651
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1606821651
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1606821651
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1606821651
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1606821651
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606821651
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1606821651
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1606821651
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1606821651
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606821651
transform 1 0 19964 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1606821651
transform 1 0 19136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1606821651
transform 1 0 19872 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606821651
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1606821651
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606821651
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606821651
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606821651
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1606821651
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1606821651
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1606821651
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1606821651
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606821651
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1606821651
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1606821651
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606821651
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1606821651
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1606821651
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1606821651
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1606821651
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1606821651
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1606821651
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1606821651
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1606821651
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14168 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1606821651
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1606821651
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_135
timestamp 1606821651
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1606821651
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_166
timestamp 1606821651
transform 1 0 16376 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_148
timestamp 1606821651
transform 1 0 14720 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_160
timestamp 1606821651
transform 1 0 15824 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17020 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_172
timestamp 1606821651
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_179
timestamp 1606821651
transform 1 0 17572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_172
timestamp 1606821651
transform 1 0 16928 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1606821651
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606821651
transform 1 0 19964 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19596 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_191
timestamp 1606821651
transform 1 0 18676 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1606821651
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_207
timestamp 1606821651
transform 1 0 20148 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1606821651
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1606821651
transform 1 0 19872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1606821651
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1606821651
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606821651
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606821651
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606821651
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1606821651
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1606821651
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606821651
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606821651
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1606821651
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1606821651
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11408 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_105
timestamp 1606821651
transform 1 0 10764 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_111
timestamp 1606821651
transform 1 0 11316 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_118
timestamp 1606821651
transform 1 0 11960 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_130
timestamp 1606821651
transform 1 0 13064 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_142
timestamp 1606821651
transform 1 0 14168 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1606821651
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_158
timestamp 1606821651
transform 1 0 15640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_170
timestamp 1606821651
transform 1 0 16744 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_182
timestamp 1606821651
transform 1 0 17848 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606821651
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_194
timestamp 1606821651
transform 1 0 18952 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1606821651
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606821651
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606821651
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1606821651
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1606821651
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1606821651
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1606821651
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606821651
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_62
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 7728 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_70
timestamp 1606821651
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_78
timestamp 1606821651
transform 1 0 8280 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_90
timestamp 1606821651
transform 1 0 9384 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_102
timestamp 1606821651
transform 1 0 10488 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1606821651
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1606821651
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1606821651
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1606821651
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606821651
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606821651
transform 1 0 19964 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_196
timestamp 1606821651
transform 1 0 19136 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1606821651
transform 1 0 19872 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606821651
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1606821651
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606821651
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606821651
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1606821651
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1606821651
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606821651
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1606821651
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1606821651
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1606821651
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1606821651
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12052 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_111
timestamp 1606821651
transform 1 0 11316 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_125
timestamp 1606821651
transform 1 0 12604 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_137
timestamp 1606821651
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15640 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1606821651
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_164
timestamp 1606821651
transform 1 0 16192 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17572 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_176
timestamp 1606821651
transform 1 0 17296 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_185
timestamp 1606821651
transform 1 0 18124 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19596 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1606821651
transform 1 0 19228 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_207
timestamp 1606821651
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1606821651
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606821651
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1606821651
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1606821651
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1606821651
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606821651
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1606821651
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1606821651
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1606821651
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1606821651
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1606821651
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1606821651
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1606821651
transform 1 0 15732 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606821651
transform 1 0 18308 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606821651
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1606821651
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_184
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606821651
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_191
timestamp 1606821651
transform 1 0 18676 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1606821651
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606821651
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1606821651
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606821651
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606821651
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606821651
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606821651
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606821651
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606821651
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606821651
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606821651
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606821651
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606821651
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606821651
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606821651
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606821651
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1606821651
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606821651
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606821651
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 5722 22320 5778 22800 6 SC_IN_TOP
port 0 nsew default input
rlabel metal2 s 22466 0 22522 480 6 SC_OUT_BOT
port 1 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_1_
port 2 nsew default input
rlabel metal2 s 17130 22320 17186 22800 6 ccff_head
port 3 nsew default input
rlabel metal3 s 0 11432 480 11552 6 ccff_tail
port 4 nsew default tristate
rlabel metal3 s 22320 3680 22800 3800 6 chanx_right_in[0]
port 5 nsew default input
rlabel metal3 s 22320 8304 22800 8424 6 chanx_right_in[10]
port 6 nsew default input
rlabel metal3 s 22320 8712 22800 8832 6 chanx_right_in[11]
port 7 nsew default input
rlabel metal3 s 22320 9256 22800 9376 6 chanx_right_in[12]
port 8 nsew default input
rlabel metal3 s 22320 9664 22800 9784 6 chanx_right_in[13]
port 9 nsew default input
rlabel metal3 s 22320 10072 22800 10192 6 chanx_right_in[14]
port 10 nsew default input
rlabel metal3 s 22320 10616 22800 10736 6 chanx_right_in[15]
port 11 nsew default input
rlabel metal3 s 22320 11024 22800 11144 6 chanx_right_in[16]
port 12 nsew default input
rlabel metal3 s 22320 11568 22800 11688 6 chanx_right_in[17]
port 13 nsew default input
rlabel metal3 s 22320 11976 22800 12096 6 chanx_right_in[18]
port 14 nsew default input
rlabel metal3 s 22320 12384 22800 12504 6 chanx_right_in[19]
port 15 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 16 nsew default input
rlabel metal3 s 22320 4632 22800 4752 6 chanx_right_in[2]
port 17 nsew default input
rlabel metal3 s 22320 5040 22800 5160 6 chanx_right_in[3]
port 18 nsew default input
rlabel metal3 s 22320 5584 22800 5704 6 chanx_right_in[4]
port 19 nsew default input
rlabel metal3 s 22320 5992 22800 6112 6 chanx_right_in[5]
port 20 nsew default input
rlabel metal3 s 22320 6536 22800 6656 6 chanx_right_in[6]
port 21 nsew default input
rlabel metal3 s 22320 6944 22800 7064 6 chanx_right_in[7]
port 22 nsew default input
rlabel metal3 s 22320 7352 22800 7472 6 chanx_right_in[8]
port 23 nsew default input
rlabel metal3 s 22320 7896 22800 8016 6 chanx_right_in[9]
port 24 nsew default input
rlabel metal3 s 22320 12928 22800 13048 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal3 s 22320 17416 22800 17536 6 chanx_right_out[10]
port 26 nsew default tristate
rlabel metal3 s 22320 17960 22800 18080 6 chanx_right_out[11]
port 27 nsew default tristate
rlabel metal3 s 22320 18368 22800 18488 6 chanx_right_out[12]
port 28 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[13]
port 29 nsew default tristate
rlabel metal3 s 22320 19320 22800 19440 6 chanx_right_out[14]
port 30 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[15]
port 31 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[16]
port 32 nsew default tristate
rlabel metal3 s 22320 20680 22800 20800 6 chanx_right_out[17]
port 33 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[18]
port 34 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[19]
port 35 nsew default tristate
rlabel metal3 s 22320 13336 22800 13456 6 chanx_right_out[1]
port 36 nsew default tristate
rlabel metal3 s 22320 13744 22800 13864 6 chanx_right_out[2]
port 37 nsew default tristate
rlabel metal3 s 22320 14288 22800 14408 6 chanx_right_out[3]
port 38 nsew default tristate
rlabel metal3 s 22320 14696 22800 14816 6 chanx_right_out[4]
port 39 nsew default tristate
rlabel metal3 s 22320 15104 22800 15224 6 chanx_right_out[5]
port 40 nsew default tristate
rlabel metal3 s 22320 15648 22800 15768 6 chanx_right_out[6]
port 41 nsew default tristate
rlabel metal3 s 22320 16056 22800 16176 6 chanx_right_out[7]
port 42 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[8]
port 43 nsew default tristate
rlabel metal3 s 22320 17008 22800 17128 6 chanx_right_out[9]
port 44 nsew default tristate
rlabel metal2 s 662 0 718 480 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[10]
port 46 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[11]
port 47 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[12]
port 48 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[13]
port 49 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chany_bottom_in[14]
port 50 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[15]
port 51 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[16]
port 52 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[17]
port 53 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[18]
port 54 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[19]
port 55 nsew default input
rlabel metal2 s 1214 0 1270 480 6 chany_bottom_in[1]
port 56 nsew default input
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_in[2]
port 57 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[3]
port 58 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[4]
port 59 nsew default input
rlabel metal2 s 3422 0 3478 480 6 chany_bottom_in[5]
port 60 nsew default input
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_in[6]
port 61 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[7]
port 62 nsew default input
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[8]
port 63 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chany_bottom_in[9]
port 64 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_out[0]
port 65 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[10]
port 66 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chany_bottom_out[11]
port 67 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[12]
port 68 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[13]
port 69 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[14]
port 70 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[15]
port 71 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[16]
port 72 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[17]
port 73 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[18]
port 74 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[19]
port 75 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_out[1]
port 76 nsew default tristate
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_out[2]
port 77 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[3]
port 78 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[4]
port 79 nsew default tristate
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_out[5]
port 80 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_out[6]
port 81 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[7]
port 82 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[8]
port 83 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[9]
port 84 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 prog_clk_0_E_in
port 85 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 86 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 87 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 88 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 89 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 90 nsew default input
rlabel metal3 s 22320 2320 22800 2440 6 right_bottom_grid_pin_39_
port 91 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 92 nsew default input
rlabel metal3 s 22320 3272 22800 3392 6 right_bottom_grid_pin_41_
port 93 nsew default input
rlabel metal3 s 22320 22448 22800 22568 6 right_top_grid_pin_1_
port 94 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 95 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 96 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
